##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Mon May 30 03:23:00 2022
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO azadi_soc_top_caravel
  CLASS BLOCK ;
  SIZE 2399.820000 BY 2500.020000 ;
  FOREIGN azadi_soc_top_caravel 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 4.680000 0.000000 4.980000 0.800000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2496.850000 0.800000 2497.150000 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 505.620000 0.000000 505.920000 0.800000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 169.820000 0.000000 170.120000 0.800000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 510.680000 0.000000 510.980000 0.800000 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 501.020000 0.000000 501.320000 0.800000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 495.960000 0.000000 496.260000 0.800000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 491.360000 0.000000 491.660000 0.800000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 486.300000 0.000000 486.600000 0.800000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 325.760000 0.000000 326.060000 0.800000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 320.700000 0.000000 321.000000 0.800000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 316.100000 0.000000 316.400000 0.800000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 311.040000 0.000000 311.340000 0.800000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 306.440000 0.000000 306.740000 0.800000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 301.380000 0.000000 301.680000 0.800000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.320000 0.000000 296.620000 0.800000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 291.720000 0.000000 292.020000 0.800000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 286.660000 0.000000 286.960000 0.800000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 282.060000 0.000000 282.360000 0.800000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 277.000000 0.000000 277.300000 0.800000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 272.400000 0.000000 272.700000 0.800000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 267.340000 0.000000 267.640000 0.800000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.280000 0.000000 262.580000 0.800000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 257.680000 0.000000 257.980000 0.800000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 252.620000 0.000000 252.920000 0.800000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 248.020000 0.000000 248.320000 0.800000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 242.960000 0.000000 243.260000 0.800000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 237.900000 0.000000 238.200000 0.800000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 233.300000 0.000000 233.600000 0.800000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 228.240000 0.000000 228.540000 0.800000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 223.640000 0.000000 223.940000 0.800000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.580000 0.000000 218.880000 0.800000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.980000 0.000000 214.280000 0.800000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 208.920000 0.000000 209.220000 0.800000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 203.860000 0.000000 204.160000 0.800000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 199.260000 0.000000 199.560000 0.800000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 194.200000 0.000000 194.500000 0.800000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 189.600000 0.000000 189.900000 0.800000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 184.540000 0.000000 184.840000 0.800000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 179.480000 0.000000 179.780000 0.800000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 174.880000 0.000000 175.180000 0.800000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 165.220000 0.000000 165.520000 0.800000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 160.160000 0.000000 160.460000 0.800000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 155.560000 0.000000 155.860000 0.800000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 150.500000 0.000000 150.800000 0.800000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 145.440000 0.000000 145.740000 0.800000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.840000 0.000000 141.140000 0.800000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 135.780000 0.000000 136.080000 0.800000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.180000 0.000000 131.480000 0.800000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.120000 0.000000 126.420000 0.800000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.520000 0.000000 121.820000 0.800000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.460000 0.000000 116.760000 0.800000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.400000 0.000000 111.700000 0.800000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.800000 0.000000 107.100000 0.800000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.740000 0.000000 102.040000 0.800000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 97.140000 0.000000 97.440000 0.800000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 92.080000 0.000000 92.380000 0.800000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 87.020000 0.000000 87.320000 0.800000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 82.420000 0.000000 82.720000 0.800000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 77.360000 0.000000 77.660000 0.800000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 72.760000 0.000000 73.060000 0.800000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 67.700000 0.000000 68.000000 0.800000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 63.100000 0.000000 63.400000 0.800000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 58.040000 0.000000 58.340000 0.800000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 52.980000 0.000000 53.280000 0.800000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 48.380000 0.000000 48.680000 0.800000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 43.320000 0.000000 43.620000 0.800000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 38.720000 0.000000 39.020000 0.800000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 33.660000 0.000000 33.960000 0.800000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.600000 0.000000 28.900000 0.800000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 24.000000 0.000000 24.300000 0.800000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 18.940000 0.000000 19.240000 0.800000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 14.340000 0.000000 14.640000 0.800000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 9.280000 0.000000 9.580000 0.800000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 481.240000 0.000000 481.540000 0.800000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.640000 0.000000 476.940000 0.800000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 471.580000 0.000000 471.880000 0.800000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 466.980000 0.000000 467.280000 0.800000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.920000 0.000000 462.220000 0.800000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 457.320000 0.000000 457.620000 0.800000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 452.260000 0.000000 452.560000 0.800000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 447.200000 0.000000 447.500000 0.800000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 442.600000 0.000000 442.900000 0.800000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 437.540000 0.000000 437.840000 0.800000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 432.940000 0.000000 433.240000 0.800000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.880000 0.000000 428.180000 0.800000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 423.280000 0.000000 423.580000 0.800000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 418.220000 0.000000 418.520000 0.800000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 413.160000 0.000000 413.460000 0.800000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 408.560000 0.000000 408.860000 0.800000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 403.500000 0.000000 403.800000 0.800000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 398.900000 0.000000 399.200000 0.800000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.840000 0.000000 394.140000 0.800000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 388.780000 0.000000 389.080000 0.800000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 384.180000 0.000000 384.480000 0.800000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 379.120000 0.000000 379.420000 0.800000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 374.520000 0.000000 374.820000 0.800000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 369.460000 0.000000 369.760000 0.800000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 364.860000 0.000000 365.160000 0.800000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 359.800000 0.000000 360.100000 0.800000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 354.740000 0.000000 355.040000 0.800000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 350.140000 0.000000 350.440000 0.800000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 345.080000 0.000000 345.380000 0.800000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 340.480000 0.000000 340.780000 0.800000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 335.420000 0.000000 335.720000 0.800000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 330.360000 0.000000 330.660000 0.800000 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1133.520000 0.000000 1133.820000 0.800000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1128.920000 0.000000 1129.220000 0.800000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1123.860000 0.000000 1124.160000 0.800000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1119.260000 0.000000 1119.560000 0.800000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1114.200000 0.000000 1114.500000 0.800000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1109.140000 0.000000 1109.440000 0.800000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1104.540000 0.000000 1104.840000 0.800000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1099.480000 0.000000 1099.780000 0.800000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1094.880000 0.000000 1095.180000 0.800000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1089.820000 0.000000 1090.120000 0.800000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1084.760000 0.000000 1085.060000 0.800000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1080.160000 0.000000 1080.460000 0.800000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1075.100000 0.000000 1075.400000 0.800000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1070.500000 0.000000 1070.800000 0.800000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1065.440000 0.000000 1065.740000 0.800000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1060.840000 0.000000 1061.140000 0.800000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1055.780000 0.000000 1056.080000 0.800000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1050.720000 0.000000 1051.020000 0.800000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1046.120000 0.000000 1046.420000 0.800000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1041.060000 0.000000 1041.360000 0.800000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1036.460000 0.000000 1036.760000 0.800000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1031.400000 0.000000 1031.700000 0.800000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1026.340000 0.000000 1026.640000 0.800000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1021.740000 0.000000 1022.040000 0.800000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1016.680000 0.000000 1016.980000 0.800000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1012.080000 0.000000 1012.380000 0.800000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1007.020000 0.000000 1007.320000 0.800000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1002.420000 0.000000 1002.720000 0.800000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 997.360000 0.000000 997.660000 0.800000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 992.300000 0.000000 992.600000 0.800000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 987.700000 0.000000 988.000000 0.800000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 982.640000 0.000000 982.940000 0.800000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 978.040000 0.000000 978.340000 0.800000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 972.980000 0.000000 973.280000 0.800000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 968.380000 0.000000 968.680000 0.800000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 963.320000 0.000000 963.620000 0.800000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 958.260000 0.000000 958.560000 0.800000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 953.660000 0.000000 953.960000 0.800000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 948.600000 0.000000 948.900000 0.800000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 944.000000 0.000000 944.300000 0.800000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 938.940000 0.000000 939.240000 0.800000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 933.880000 0.000000 934.180000 0.800000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 929.280000 0.000000 929.580000 0.800000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 924.220000 0.000000 924.520000 0.800000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 919.620000 0.000000 919.920000 0.800000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 914.560000 0.000000 914.860000 0.800000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 909.960000 0.000000 910.260000 0.800000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 904.900000 0.000000 905.200000 0.800000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 899.840000 0.000000 900.140000 0.800000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 895.240000 0.000000 895.540000 0.800000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.180000 0.000000 890.480000 0.800000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 885.580000 0.000000 885.880000 0.800000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 880.520000 0.000000 880.820000 0.800000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 875.460000 0.000000 875.760000 0.800000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 870.860000 0.000000 871.160000 0.800000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 865.800000 0.000000 866.100000 0.800000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 861.200000 0.000000 861.500000 0.800000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 856.140000 0.000000 856.440000 0.800000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 851.540000 0.000000 851.840000 0.800000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.480000 0.000000 846.780000 0.800000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 841.420000 0.000000 841.720000 0.800000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.820000 0.000000 837.120000 0.800000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 831.760000 0.000000 832.060000 0.800000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 827.160000 0.000000 827.460000 0.800000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 822.100000 0.000000 822.400000 0.800000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.500000 0.000000 817.800000 0.800000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 812.440000 0.000000 812.740000 0.800000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 807.380000 0.000000 807.680000 0.800000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 802.780000 0.000000 803.080000 0.800000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 797.720000 0.000000 798.020000 0.800000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 793.120000 0.000000 793.420000 0.800000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 788.060000 0.000000 788.360000 0.800000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 783.000000 0.000000 783.300000 0.800000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 778.400000 0.000000 778.700000 0.800000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 773.340000 0.000000 773.640000 0.800000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 768.740000 0.000000 769.040000 0.800000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 763.680000 0.000000 763.980000 0.800000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 759.080000 0.000000 759.380000 0.800000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 754.020000 0.000000 754.320000 0.800000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 748.960000 0.000000 749.260000 0.800000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 744.360000 0.000000 744.660000 0.800000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 739.300000 0.000000 739.600000 0.800000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 734.700000 0.000000 735.000000 0.800000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 729.640000 0.000000 729.940000 0.800000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 724.580000 0.000000 724.880000 0.800000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 719.980000 0.000000 720.280000 0.800000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 714.920000 0.000000 715.220000 0.800000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 710.320000 0.000000 710.620000 0.800000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 705.260000 0.000000 705.560000 0.800000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 700.660000 0.000000 700.960000 0.800000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 695.600000 0.000000 695.900000 0.800000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 690.540000 0.000000 690.840000 0.800000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 685.940000 0.000000 686.240000 0.800000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 680.880000 0.000000 681.180000 0.800000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.280000 0.000000 676.580000 0.800000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 671.220000 0.000000 671.520000 0.800000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 666.620000 0.000000 666.920000 0.800000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 661.560000 0.000000 661.860000 0.800000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 656.500000 0.000000 656.800000 0.800000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 651.900000 0.000000 652.200000 0.800000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.840000 0.000000 647.140000 0.800000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 642.240000 0.000000 642.540000 0.800000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 637.180000 0.000000 637.480000 0.800000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 632.120000 0.000000 632.420000 0.800000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 627.520000 0.000000 627.820000 0.800000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 622.460000 0.000000 622.760000 0.800000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 617.860000 0.000000 618.160000 0.800000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 612.800000 0.000000 613.100000 0.800000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 608.200000 0.000000 608.500000 0.800000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 603.140000 0.000000 603.440000 0.800000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 598.080000 0.000000 598.380000 0.800000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 593.480000 0.000000 593.780000 0.800000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 588.420000 0.000000 588.720000 0.800000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.820000 0.000000 584.120000 0.800000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 578.760000 0.000000 579.060000 0.800000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 573.700000 0.000000 574.000000 0.800000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 569.100000 0.000000 569.400000 0.800000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 564.040000 0.000000 564.340000 0.800000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 559.440000 0.000000 559.740000 0.800000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 554.380000 0.000000 554.680000 0.800000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 549.780000 0.000000 550.080000 0.800000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 544.720000 0.000000 545.020000 0.800000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 539.660000 0.000000 539.960000 0.800000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 535.060000 0.000000 535.360000 0.800000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 530.000000 0.000000 530.300000 0.800000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 525.400000 0.000000 525.700000 0.800000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 520.340000 0.000000 520.640000 0.800000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 515.740000 0.000000 516.040000 0.800000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1756.820000 0.000000 1757.120000 0.800000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1751.760000 0.000000 1752.060000 0.800000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1746.700000 0.000000 1747.000000 0.800000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1742.100000 0.000000 1742.400000 0.800000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1737.040000 0.000000 1737.340000 0.800000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1732.440000 0.000000 1732.740000 0.800000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1727.380000 0.000000 1727.680000 0.800000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1722.320000 0.000000 1722.620000 0.800000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1717.720000 0.000000 1718.020000 0.800000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1712.660000 0.000000 1712.960000 0.800000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1708.060000 0.000000 1708.360000 0.800000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1703.000000 0.000000 1703.300000 0.800000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1698.400000 0.000000 1698.700000 0.800000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1693.340000 0.000000 1693.640000 0.800000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1688.280000 0.000000 1688.580000 0.800000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1683.680000 0.000000 1683.980000 0.800000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1678.620000 0.000000 1678.920000 0.800000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1674.020000 0.000000 1674.320000 0.800000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1668.960000 0.000000 1669.260000 0.800000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1664.360000 0.000000 1664.660000 0.800000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1659.300000 0.000000 1659.600000 0.800000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1654.240000 0.000000 1654.540000 0.800000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1649.640000 0.000000 1649.940000 0.800000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1644.580000 0.000000 1644.880000 0.800000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1639.980000 0.000000 1640.280000 0.800000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1634.920000 0.000000 1635.220000 0.800000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1629.860000 0.000000 1630.160000 0.800000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1625.260000 0.000000 1625.560000 0.800000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1620.200000 0.000000 1620.500000 0.800000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1615.600000 0.000000 1615.900000 0.800000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1610.540000 0.000000 1610.840000 0.800000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1605.940000 0.000000 1606.240000 0.800000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1600.880000 0.000000 1601.180000 0.800000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1595.820000 0.000000 1596.120000 0.800000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1591.220000 0.000000 1591.520000 0.800000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1586.160000 0.000000 1586.460000 0.800000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.560000 0.000000 1581.860000 0.800000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1576.500000 0.000000 1576.800000 0.800000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1571.440000 0.000000 1571.740000 0.800000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1566.840000 0.000000 1567.140000 0.800000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1561.780000 0.000000 1562.080000 0.800000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1557.180000 0.000000 1557.480000 0.800000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1552.120000 0.000000 1552.420000 0.800000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1547.520000 0.000000 1547.820000 0.800000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1542.460000 0.000000 1542.760000 0.800000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1537.400000 0.000000 1537.700000 0.800000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1532.800000 0.000000 1533.100000 0.800000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1527.740000 0.000000 1528.040000 0.800000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1523.140000 0.000000 1523.440000 0.800000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1518.080000 0.000000 1518.380000 0.800000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1513.480000 0.000000 1513.780000 0.800000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1508.420000 0.000000 1508.720000 0.800000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1503.360000 0.000000 1503.660000 0.800000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1498.760000 0.000000 1499.060000 0.800000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1493.700000 0.000000 1494.000000 0.800000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1489.100000 0.000000 1489.400000 0.800000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1484.040000 0.000000 1484.340000 0.800000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1478.980000 0.000000 1479.280000 0.800000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1474.380000 0.000000 1474.680000 0.800000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1469.320000 0.000000 1469.620000 0.800000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1464.720000 0.000000 1465.020000 0.800000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1459.660000 0.000000 1459.960000 0.800000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1455.060000 0.000000 1455.360000 0.800000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1450.000000 0.000000 1450.300000 0.800000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1444.940000 0.000000 1445.240000 0.800000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1440.340000 0.000000 1440.640000 0.800000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1435.280000 0.000000 1435.580000 0.800000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1430.680000 0.000000 1430.980000 0.800000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1425.620000 0.000000 1425.920000 0.800000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1420.560000 0.000000 1420.860000 0.800000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1415.960000 0.000000 1416.260000 0.800000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1410.900000 0.000000 1411.200000 0.800000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1406.300000 0.000000 1406.600000 0.800000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1401.240000 0.000000 1401.540000 0.800000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.640000 0.000000 1396.940000 0.800000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1391.580000 0.000000 1391.880000 0.800000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1386.520000 0.000000 1386.820000 0.800000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1381.920000 0.000000 1382.220000 0.800000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1376.860000 0.000000 1377.160000 0.800000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1372.260000 0.000000 1372.560000 0.800000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1367.200000 0.000000 1367.500000 0.800000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1362.600000 0.000000 1362.900000 0.800000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1357.540000 0.000000 1357.840000 0.800000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1352.480000 0.000000 1352.780000 0.800000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1347.880000 0.000000 1348.180000 0.800000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1342.820000 0.000000 1343.120000 0.800000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1338.220000 0.000000 1338.520000 0.800000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1333.160000 0.000000 1333.460000 0.800000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1328.100000 0.000000 1328.400000 0.800000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1323.500000 0.000000 1323.800000 0.800000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1318.440000 0.000000 1318.740000 0.800000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1313.840000 0.000000 1314.140000 0.800000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1308.780000 0.000000 1309.080000 0.800000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1304.180000 0.000000 1304.480000 0.800000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1299.120000 0.000000 1299.420000 0.800000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1294.060000 0.000000 1294.360000 0.800000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1289.460000 0.000000 1289.760000 0.800000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1284.400000 0.000000 1284.700000 0.800000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1279.800000 0.000000 1280.100000 0.800000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1274.740000 0.000000 1275.040000 0.800000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1269.680000 0.000000 1269.980000 0.800000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1265.080000 0.000000 1265.380000 0.800000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1260.020000 0.000000 1260.320000 0.800000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1255.420000 0.000000 1255.720000 0.800000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1250.360000 0.000000 1250.660000 0.800000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1245.760000 0.000000 1246.060000 0.800000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1240.700000 0.000000 1241.000000 0.800000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1235.640000 0.000000 1235.940000 0.800000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1231.040000 0.000000 1231.340000 0.800000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1225.980000 0.000000 1226.280000 0.800000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1221.380000 0.000000 1221.680000 0.800000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1216.320000 0.000000 1216.620000 0.800000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1211.720000 0.000000 1212.020000 0.800000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1206.660000 0.000000 1206.960000 0.800000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1201.600000 0.000000 1201.900000 0.800000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1197.000000 0.000000 1197.300000 0.800000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1191.940000 0.000000 1192.240000 0.800000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1187.340000 0.000000 1187.640000 0.800000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1182.280000 0.000000 1182.580000 0.800000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1177.220000 0.000000 1177.520000 0.800000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1172.620000 0.000000 1172.920000 0.800000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1167.560000 0.000000 1167.860000 0.800000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1162.960000 0.000000 1163.260000 0.800000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1157.900000 0.000000 1158.200000 0.800000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1153.300000 0.000000 1153.600000 0.800000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1148.240000 0.000000 1148.540000 0.800000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1143.180000 0.000000 1143.480000 0.800000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1138.580000 0.000000 1138.880000 0.800000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2379.660000 0.000000 2379.960000 0.800000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2374.600000 0.000000 2374.900000 0.800000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2370.000000 0.000000 2370.300000 0.800000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2364.940000 0.000000 2365.240000 0.800000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2360.340000 0.000000 2360.640000 0.800000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2355.280000 0.000000 2355.580000 0.800000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2350.220000 0.000000 2350.520000 0.800000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2345.620000 0.000000 2345.920000 0.800000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2340.560000 0.000000 2340.860000 0.800000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2335.960000 0.000000 2336.260000 0.800000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2330.900000 0.000000 2331.200000 0.800000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2325.840000 0.000000 2326.140000 0.800000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2321.240000 0.000000 2321.540000 0.800000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2316.180000 0.000000 2316.480000 0.800000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2311.580000 0.000000 2311.880000 0.800000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2306.520000 0.000000 2306.820000 0.800000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2301.920000 0.000000 2302.220000 0.800000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.860000 0.000000 2297.160000 0.800000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2291.800000 0.000000 2292.100000 0.800000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2287.200000 0.000000 2287.500000 0.800000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2282.140000 0.000000 2282.440000 0.800000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2277.540000 0.000000 2277.840000 0.800000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2272.480000 0.000000 2272.780000 0.800000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2267.420000 0.000000 2267.720000 0.800000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2262.820000 0.000000 2263.120000 0.800000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2257.760000 0.000000 2258.060000 0.800000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2253.160000 0.000000 2253.460000 0.800000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2248.100000 0.000000 2248.400000 0.800000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2243.500000 0.000000 2243.800000 0.800000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.440000 0.000000 2238.740000 0.800000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2233.380000 0.000000 2233.680000 0.800000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2228.780000 0.000000 2229.080000 0.800000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2223.720000 0.000000 2224.020000 0.800000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.120000 0.000000 2219.420000 0.800000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2214.060000 0.000000 2214.360000 0.800000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2209.460000 0.000000 2209.760000 0.800000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2204.400000 0.000000 2204.700000 0.800000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2199.340000 0.000000 2199.640000 0.800000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2194.740000 0.000000 2195.040000 0.800000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2189.680000 0.000000 2189.980000 0.800000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2185.080000 0.000000 2185.380000 0.800000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2180.020000 0.000000 2180.320000 0.800000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2174.960000 0.000000 2175.260000 0.800000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2170.360000 0.000000 2170.660000 0.800000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2165.300000 0.000000 2165.600000 0.800000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2160.700000 0.000000 2161.000000 0.800000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2155.640000 0.000000 2155.940000 0.800000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2151.040000 0.000000 2151.340000 0.800000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2145.980000 0.000000 2146.280000 0.800000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2140.920000 0.000000 2141.220000 0.800000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2136.320000 0.000000 2136.620000 0.800000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2131.260000 0.000000 2131.560000 0.800000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2126.660000 0.000000 2126.960000 0.800000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2121.600000 0.000000 2121.900000 0.800000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2116.540000 0.000000 2116.840000 0.800000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2111.940000 0.000000 2112.240000 0.800000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2106.880000 0.000000 2107.180000 0.800000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2102.280000 0.000000 2102.580000 0.800000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2097.220000 0.000000 2097.520000 0.800000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2092.620000 0.000000 2092.920000 0.800000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2087.560000 0.000000 2087.860000 0.800000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2082.500000 0.000000 2082.800000 0.800000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2077.900000 0.000000 2078.200000 0.800000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2072.840000 0.000000 2073.140000 0.800000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2068.240000 0.000000 2068.540000 0.800000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2063.180000 0.000000 2063.480000 0.800000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2058.580000 0.000000 2058.880000 0.800000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2053.520000 0.000000 2053.820000 0.800000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2048.460000 0.000000 2048.760000 0.800000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2043.860000 0.000000 2044.160000 0.800000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2038.800000 0.000000 2039.100000 0.800000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2034.200000 0.000000 2034.500000 0.800000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2029.140000 0.000000 2029.440000 0.800000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2024.080000 0.000000 2024.380000 0.800000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2019.480000 0.000000 2019.780000 0.800000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2014.420000 0.000000 2014.720000 0.800000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2009.820000 0.000000 2010.120000 0.800000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2004.760000 0.000000 2005.060000 0.800000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2000.160000 0.000000 2000.460000 0.800000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1995.100000 0.000000 1995.400000 0.800000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1990.040000 0.000000 1990.340000 0.800000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1985.440000 0.000000 1985.740000 0.800000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1980.380000 0.000000 1980.680000 0.800000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1975.780000 0.000000 1976.080000 0.800000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1970.720000 0.000000 1971.020000 0.800000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1966.120000 0.000000 1966.420000 0.800000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1961.060000 0.000000 1961.360000 0.800000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1956.000000 0.000000 1956.300000 0.800000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1951.400000 0.000000 1951.700000 0.800000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.340000 0.000000 1946.640000 0.800000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1941.740000 0.000000 1942.040000 0.800000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1936.680000 0.000000 1936.980000 0.800000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1931.620000 0.000000 1931.920000 0.800000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1927.020000 0.000000 1927.320000 0.800000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1921.960000 0.000000 1922.260000 0.800000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1917.360000 0.000000 1917.660000 0.800000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1912.300000 0.000000 1912.600000 0.800000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1907.700000 0.000000 1908.000000 0.800000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1902.640000 0.000000 1902.940000 0.800000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1897.580000 0.000000 1897.880000 0.800000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1892.980000 0.000000 1893.280000 0.800000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1887.920000 0.000000 1888.220000 0.800000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1883.320000 0.000000 1883.620000 0.800000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1878.260000 0.000000 1878.560000 0.800000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1873.200000 0.000000 1873.500000 0.800000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1868.600000 0.000000 1868.900000 0.800000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1863.540000 0.000000 1863.840000 0.800000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1858.940000 0.000000 1859.240000 0.800000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1853.880000 0.000000 1854.180000 0.800000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1849.280000 0.000000 1849.580000 0.800000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1844.220000 0.000000 1844.520000 0.800000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1839.160000 0.000000 1839.460000 0.800000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1834.560000 0.000000 1834.860000 0.800000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1829.500000 0.000000 1829.800000 0.800000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1824.900000 0.000000 1825.200000 0.800000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1819.840000 0.000000 1820.140000 0.800000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1815.240000 0.000000 1815.540000 0.800000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1810.180000 0.000000 1810.480000 0.800000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1805.120000 0.000000 1805.420000 0.800000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1800.520000 0.000000 1800.820000 0.800000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1795.460000 0.000000 1795.760000 0.800000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1790.860000 0.000000 1791.160000 0.800000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1785.800000 0.000000 1786.100000 0.800000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1780.740000 0.000000 1781.040000 0.800000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1776.140000 0.000000 1776.440000 0.800000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1771.080000 0.000000 1771.380000 0.800000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1766.480000 0.000000 1766.780000 0.800000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1761.420000 0.000000 1761.720000 0.800000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1131.670000 0.800000 1131.970000 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1084.700000 0.800000 1085.000000 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1037.730000 0.800000 1038.030000 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 990.150000 0.800000 990.450000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 943.180000 0.800000 943.480000 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 896.210000 0.800000 896.510000 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 849.240000 0.800000 849.540000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 801.660000 0.800000 801.960000 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 754.690000 0.800000 754.990000 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 707.720000 0.800000 708.020000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 660.140000 0.800000 660.440000 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 613.170000 0.800000 613.470000 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 566.200000 0.800000 566.500000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 519.230000 0.800000 519.530000 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 137.160000 2499.220000 137.460000 2500.020000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 411.320000 2499.220000 411.620000 2500.020000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 685.940000 2499.220000 686.240000 2500.020000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 960.100000 2499.220000 960.400000 2500.020000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1234.260000 2499.220000 1234.560000 2500.020000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1508.420000 2499.220000 1508.720000 2500.020000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1782.580000 2499.220000 1782.880000 2500.020000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2057.200000 2499.220000 2057.500000 2500.020000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2331.360000 2499.220000 2331.660000 2500.020000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1394.580000 2399.820000 1394.880000 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1442.770000 2399.820000 1443.070000 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1490.350000 2399.820000 1490.650000 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1538.540000 2399.820000 1538.840000 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1586.730000 2399.820000 1587.030000 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1634.920000 2399.820000 1635.220000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1682.500000 2399.820000 1682.800000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1730.690000 2399.820000 1730.990000 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1778.880000 2399.820000 1779.180000 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1827.070000 2399.820000 1827.370000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1875.260000 2399.820000 1875.560000 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1922.840000 2399.820000 1923.140000 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1971.030000 2399.820000 1971.330000 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 2019.220000 2399.820000 2019.520000 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 2067.410000 2399.820000 2067.710000 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2451.710000 0.800000 2452.010000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2404.740000 0.800000 2405.040000 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2357.770000 0.800000 2358.070000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2310.190000 0.800000 2310.490000 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2263.220000 0.800000 2263.520000 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2216.250000 0.800000 2216.550000 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2169.280000 0.800000 2169.580000 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2121.700000 0.800000 2122.000000 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2074.730000 0.800000 2075.030000 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2027.760000 0.800000 2028.060000 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1980.180000 0.800000 1980.480000 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1933.210000 0.800000 1933.510000 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1886.240000 0.800000 1886.540000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1839.270000 0.800000 1839.570000 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 68.620000 2499.220000 68.920000 2500.020000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 342.780000 2499.220000 343.080000 2500.020000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 617.400000 2499.220000 617.700000 2500.020000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.560000 2499.220000 891.860000 2500.020000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1165.720000 2499.220000 1166.020000 2500.020000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1439.880000 2499.220000 1440.180000 2500.020000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1714.040000 2499.220000 1714.340000 2500.020000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1988.660000 2499.220000 1988.960000 2500.020000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2262.820000 2499.220000 2263.120000 2500.020000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 11.710000 2399.820000 12.010000 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 48.920000 2399.820000 49.220000 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 97.110000 2399.820000 97.410000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 145.300000 2399.820000 145.600000 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 193.490000 2399.820000 193.790000 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 241.070000 2399.820000 241.370000 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 289.260000 2399.820000 289.560000 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 337.450000 2399.820000 337.750000 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 385.640000 2399.820000 385.940000 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 433.220000 2399.820000 433.520000 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 481.410000 2399.820000 481.710000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 529.600000 2399.820000 529.900000 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 577.790000 2399.820000 578.090000 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 625.370000 2399.820000 625.670000 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 673.560000 2399.820000 673.860000 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.920000 0.000000 2.220000 0.800000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1791.690000 0.800000 1791.990000 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1744.720000 0.800000 1745.020000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1697.750000 0.800000 1698.050000 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1650.170000 0.800000 1650.470000 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1603.200000 0.800000 1603.500000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1556.230000 0.800000 1556.530000 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1509.260000 0.800000 1509.560000 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1461.680000 0.800000 1461.980000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1414.710000 0.800000 1415.010000 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1367.740000 0.800000 1368.040000 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1320.160000 0.800000 1320.460000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1273.190000 0.800000 1273.490000 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1226.220000 0.800000 1226.520000 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1179.250000 0.800000 1179.550000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 274.240000 2499.220000 274.540000 2500.020000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 548.400000 2499.220000 548.700000 2500.020000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 823.020000 2499.220000 823.320000 2500.020000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1097.180000 2499.220000 1097.480000 2500.020000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1371.340000 2499.220000 1371.640000 2500.020000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1645.500000 2499.220000 1645.800000 2500.020000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1920.120000 2499.220000 1920.420000 2500.020000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2194.280000 2499.220000 2194.580000 2500.020000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2394.380000 2499.220000 2394.680000 2500.020000 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 721.750000 2399.820000 722.050000 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 769.940000 2399.820000 770.240000 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 818.130000 2399.820000 818.430000 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 865.710000 2399.820000 866.010000 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 913.900000 2399.820000 914.200000 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 962.090000 2399.820000 962.390000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1010.280000 2399.820000 1010.580000 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1057.860000 2399.820000 1058.160000 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1106.050000 2399.820000 1106.350000 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1154.240000 2399.820000 1154.540000 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1202.430000 2399.820000 1202.730000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1250.620000 2399.820000 1250.920000 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1298.200000 2399.820000 1298.500000 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1346.390000 2399.820000 1346.690000 ;
    END
  END io_oeb[0]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 471.650000 0.800000 471.950000 ;
    END
  END analog_io[28]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 424.680000 0.800000 424.980000 ;
    END
  END analog_io[27]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 377.710000 0.800000 378.010000 ;
    END
  END analog_io[26]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 330.130000 0.800000 330.430000 ;
    END
  END analog_io[25]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 283.160000 0.800000 283.460000 ;
    END
  END analog_io[24]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 236.190000 0.800000 236.490000 ;
    END
  END analog_io[23]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 189.220000 0.800000 189.520000 ;
    END
  END analog_io[22]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 141.640000 0.800000 141.940000 ;
    END
  END analog_io[21]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 94.670000 0.800000 94.970000 ;
    END
  END analog_io[20]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 47.700000 0.800000 48.000000 ;
    END
  END analog_io[19]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 6.830000 0.800000 7.130000 ;
    END
  END analog_io[18]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 4.220000 2499.220000 4.520000 2500.020000 ;
    END
  END analog_io[17]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 205.700000 2499.220000 206.000000 2500.020000 ;
    END
  END analog_io[16]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 479.860000 2499.220000 480.160000 2500.020000 ;
    END
  END analog_io[15]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 754.480000 2499.220000 754.780000 2500.020000 ;
    END
  END analog_io[14]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1028.640000 2499.220000 1028.940000 2500.020000 ;
    END
  END analog_io[13]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1302.800000 2499.220000 1303.100000 2500.020000 ;
    END
  END analog_io[12]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1576.960000 2499.220000 1577.260000 2500.020000 ;
    END
  END analog_io[11]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1851.580000 2499.220000 1851.880000 2500.020000 ;
    END
  END analog_io[10]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2125.740000 2499.220000 2126.040000 2500.020000 ;
    END
  END analog_io[9]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 2114.990000 2399.820000 2115.290000 ;
    END
  END analog_io[8]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 2163.180000 2399.820000 2163.480000 ;
    END
  END analog_io[7]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 2211.370000 2399.820000 2211.670000 ;
    END
  END analog_io[6]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 2259.560000 2399.820000 2259.860000 ;
    END
  END analog_io[5]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 2307.140000 2399.820000 2307.440000 ;
    END
  END analog_io[4]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 2355.330000 2399.820000 2355.630000 ;
    END
  END analog_io[3]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 2403.520000 2399.820000 2403.820000 ;
    END
  END analog_io[2]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 2451.710000 2399.820000 2452.010000 ;
    END
  END analog_io[1]
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 2495.630000 2399.820000 2495.930000 ;
    END
  END analog_io[0]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2384.260000 0.000000 2384.560000 0.800000 ;
    END
  END user_clock2
  PIN user_irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2394.380000 0.000000 2394.680000 0.800000 ;
    END
  END user_irq[2]
  PIN user_irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2397.600000 0.000000 2397.900000 0.800000 ;
    END
  END user_irq[1]
  PIN user_irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2389.320000 0.000000 2389.620000 0.800000 ;
    END
  END user_irq[0]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2391.500000 6.260000 2393.300000 2491.380000 ;
    END
    PORT
      LAYER met4 ;
        RECT 6.520000 6.260000 8.320000 2411.380000 ;
    END

# P/G pin shape extracted from block 'azadi_soc_top'
    PORT
      LAYER met4 ;
        RECT 724.970000 383.090000 726.710000 771.070000 ;
      LAYER met4 ;
        RECT 256.450000 383.090000 258.190000 771.070000 ;
    END
    PORT
      LAYER met4 ;
        RECT 724.970000 1314.090000 726.710000 1702.070000 ;
      LAYER met4 ;
        RECT 256.450000 1314.090000 258.190000 1702.070000 ;
    END
    PORT
      LAYER met4 ;
        RECT 724.970000 1779.590000 726.710000 2167.570000 ;
      LAYER met4 ;
        RECT 256.450000 1779.590000 258.190000 2167.570000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2151.850000 377.550000 2153.590000 765.530000 ;
      LAYER met4 ;
        RECT 1683.330000 377.550000 1685.070000 765.530000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2151.850000 843.050000 2153.590000 1231.030000 ;
      LAYER met4 ;
        RECT 1683.330000 843.050000 1685.070000 1231.030000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2151.850000 1308.550000 2153.590000 1696.530000 ;
      LAYER met4 ;
        RECT 1683.330000 1308.550000 1685.070000 1696.530000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2151.850000 1774.050000 2153.590000 2162.030000 ;
      LAYER met4 ;
        RECT 1683.330000 1774.050000 1685.070000 2162.030000 ;
    END
    PORT
      LAYER met4 ;
        RECT 724.970000 848.590000 726.710000 1236.570000 ;
      LAYER met4 ;
        RECT 256.450000 848.590000 258.190000 1236.570000 ;
    END
    PORT
      LAYER met4 ;
        RECT 212.590000 328.045000 214.390000 2214.765000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2197.830000 328.045000 2199.630000 2214.765000 ;
    END
# end of P/G pin shape extracted from block 'azadi_soc_top'

  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2.920000 2.660000 4.720000 2494.980000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2395.100000 2.660000 2396.900000 2494.980000 ;
    END

# P/G pin shape extracted from block 'azadi_soc_top'
    PORT
      LAYER met4 ;
        RECT 253.050000 379.690000 254.790000 774.470000 ;
      LAYER met4 ;
        RECT 728.370000 379.690000 730.110000 774.470000 ;
    END
    PORT
      LAYER met4 ;
        RECT 253.050000 1310.690000 254.790000 1705.470000 ;
      LAYER met4 ;
        RECT 728.370000 1310.690000 730.110000 1705.470000 ;
    END
    PORT
      LAYER met4 ;
        RECT 253.050000 1776.190000 254.790000 2170.970000 ;
      LAYER met4 ;
        RECT 728.370000 1776.190000 730.110000 2170.970000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1679.930000 374.150000 1681.670000 768.930000 ;
      LAYER met4 ;
        RECT 2155.250000 374.150000 2156.990000 768.930000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1679.930000 839.650000 1681.670000 1234.430000 ;
      LAYER met4 ;
        RECT 2155.250000 839.650000 2156.990000 1234.430000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1679.930000 1305.150000 1681.670000 1699.930000 ;
      LAYER met4 ;
        RECT 2155.250000 1305.150000 2156.990000 1699.930000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1679.930000 1770.650000 1681.670000 2165.430000 ;
      LAYER met4 ;
        RECT 2155.250000 1770.650000 2156.990000 2165.430000 ;
    END
    PORT
      LAYER met4 ;
        RECT 253.050000 845.190000 254.790000 1239.970000 ;
      LAYER met4 ;
        RECT 728.370000 845.190000 730.110000 1239.970000 ;
    END
    PORT
      LAYER met4 ;
        RECT 208.990000 324.445000 210.790000 2218.365000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2201.430000 324.445000 2203.230000 2218.365000 ;
    END
# end of P/G pin shape extracted from block 'azadi_soc_top'

  END vssd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 2399.820000 2500.020000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 2399.820000 2500.020000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 2399.820000 2500.020000 ;
    LAYER met3 ;
      RECT 2394.980000 2498.920000 2399.820000 2500.020000 ;
      RECT 2331.960000 2498.920000 2394.080000 2500.020000 ;
      RECT 2263.420000 2498.920000 2331.060000 2500.020000 ;
      RECT 2194.880000 2498.920000 2262.520000 2500.020000 ;
      RECT 2126.340000 2498.920000 2193.980000 2500.020000 ;
      RECT 2057.800000 2498.920000 2125.440000 2500.020000 ;
      RECT 1989.260000 2498.920000 2056.900000 2500.020000 ;
      RECT 1920.720000 2498.920000 1988.360000 2500.020000 ;
      RECT 1852.180000 2498.920000 1919.820000 2500.020000 ;
      RECT 1783.180000 2498.920000 1851.280000 2500.020000 ;
      RECT 1714.640000 2498.920000 1782.280000 2500.020000 ;
      RECT 1646.100000 2498.920000 1713.740000 2500.020000 ;
      RECT 1577.560000 2498.920000 1645.200000 2500.020000 ;
      RECT 1509.020000 2498.920000 1576.660000 2500.020000 ;
      RECT 1440.480000 2498.920000 1508.120000 2500.020000 ;
      RECT 1371.940000 2498.920000 1439.580000 2500.020000 ;
      RECT 1303.400000 2498.920000 1371.040000 2500.020000 ;
      RECT 1234.860000 2498.920000 1302.500000 2500.020000 ;
      RECT 1166.320000 2498.920000 1233.960000 2500.020000 ;
      RECT 1097.780000 2498.920000 1165.420000 2500.020000 ;
      RECT 1029.240000 2498.920000 1096.880000 2500.020000 ;
      RECT 960.700000 2498.920000 1028.340000 2500.020000 ;
      RECT 892.160000 2498.920000 959.800000 2500.020000 ;
      RECT 823.620000 2498.920000 891.260000 2500.020000 ;
      RECT 755.080000 2498.920000 822.720000 2500.020000 ;
      RECT 686.540000 2498.920000 754.180000 2500.020000 ;
      RECT 618.000000 2498.920000 685.640000 2500.020000 ;
      RECT 549.000000 2498.920000 617.100000 2500.020000 ;
      RECT 480.460000 2498.920000 548.100000 2500.020000 ;
      RECT 411.920000 2498.920000 479.560000 2500.020000 ;
      RECT 343.380000 2498.920000 411.020000 2500.020000 ;
      RECT 274.840000 2498.920000 342.480000 2500.020000 ;
      RECT 206.300000 2498.920000 273.940000 2500.020000 ;
      RECT 137.760000 2498.920000 205.400000 2500.020000 ;
      RECT 69.220000 2498.920000 136.860000 2500.020000 ;
      RECT 4.820000 2498.920000 68.320000 2500.020000 ;
      RECT 0.000000 2498.920000 3.920000 2500.020000 ;
      RECT 0.000000 2497.450000 2399.820000 2498.920000 ;
      RECT 1.100000 2496.550000 2399.820000 2497.450000 ;
      RECT 0.000000 2496.230000 2399.820000 2496.550000 ;
      RECT 0.000000 2495.330000 2398.720000 2496.230000 ;
      RECT 0.000000 2452.310000 2399.820000 2495.330000 ;
      RECT 1.100000 2451.410000 2398.720000 2452.310000 ;
      RECT 0.000000 2405.340000 2399.820000 2451.410000 ;
      RECT 1.100000 2404.440000 2399.820000 2405.340000 ;
      RECT 0.000000 2404.120000 2399.820000 2404.440000 ;
      RECT 0.000000 2403.220000 2398.720000 2404.120000 ;
      RECT 0.000000 2358.370000 2399.820000 2403.220000 ;
      RECT 1.100000 2357.470000 2399.820000 2358.370000 ;
      RECT 0.000000 2355.930000 2399.820000 2357.470000 ;
      RECT 0.000000 2355.030000 2398.720000 2355.930000 ;
      RECT 0.000000 2310.790000 2399.820000 2355.030000 ;
      RECT 1.100000 2309.890000 2399.820000 2310.790000 ;
      RECT 0.000000 2307.740000 2399.820000 2309.890000 ;
      RECT 0.000000 2306.840000 2398.720000 2307.740000 ;
      RECT 0.000000 2263.820000 2399.820000 2306.840000 ;
      RECT 1.100000 2262.920000 2399.820000 2263.820000 ;
      RECT 0.000000 2260.160000 2399.820000 2262.920000 ;
      RECT 0.000000 2259.260000 2398.720000 2260.160000 ;
      RECT 0.000000 2216.850000 2399.820000 2259.260000 ;
      RECT 1.100000 2215.950000 2399.820000 2216.850000 ;
      RECT 0.000000 2211.970000 2399.820000 2215.950000 ;
      RECT 0.000000 2211.070000 2398.720000 2211.970000 ;
      RECT 0.000000 2169.880000 2399.820000 2211.070000 ;
      RECT 1.100000 2168.980000 2399.820000 2169.880000 ;
      RECT 0.000000 2163.780000 2399.820000 2168.980000 ;
      RECT 0.000000 2162.880000 2398.720000 2163.780000 ;
      RECT 0.000000 2122.300000 2399.820000 2162.880000 ;
      RECT 1.100000 2121.400000 2399.820000 2122.300000 ;
      RECT 0.000000 2115.590000 2399.820000 2121.400000 ;
      RECT 0.000000 2114.690000 2398.720000 2115.590000 ;
      RECT 0.000000 2075.330000 2399.820000 2114.690000 ;
      RECT 1.100000 2074.430000 2399.820000 2075.330000 ;
      RECT 0.000000 2068.010000 2399.820000 2074.430000 ;
      RECT 0.000000 2067.110000 2398.720000 2068.010000 ;
      RECT 0.000000 2028.360000 2399.820000 2067.110000 ;
      RECT 1.100000 2027.460000 2399.820000 2028.360000 ;
      RECT 0.000000 2019.820000 2399.820000 2027.460000 ;
      RECT 0.000000 2018.920000 2398.720000 2019.820000 ;
      RECT 0.000000 1980.780000 2399.820000 2018.920000 ;
      RECT 1.100000 1979.880000 2399.820000 1980.780000 ;
      RECT 0.000000 1971.630000 2399.820000 1979.880000 ;
      RECT 0.000000 1970.730000 2398.720000 1971.630000 ;
      RECT 0.000000 1933.810000 2399.820000 1970.730000 ;
      RECT 1.100000 1932.910000 2399.820000 1933.810000 ;
      RECT 0.000000 1923.440000 2399.820000 1932.910000 ;
      RECT 0.000000 1922.540000 2398.720000 1923.440000 ;
      RECT 0.000000 1886.840000 2399.820000 1922.540000 ;
      RECT 1.100000 1885.940000 2399.820000 1886.840000 ;
      RECT 0.000000 1875.860000 2399.820000 1885.940000 ;
      RECT 0.000000 1874.960000 2398.720000 1875.860000 ;
      RECT 0.000000 1839.870000 2399.820000 1874.960000 ;
      RECT 1.100000 1838.970000 2399.820000 1839.870000 ;
      RECT 0.000000 1827.670000 2399.820000 1838.970000 ;
      RECT 0.000000 1826.770000 2398.720000 1827.670000 ;
      RECT 0.000000 1792.290000 2399.820000 1826.770000 ;
      RECT 1.100000 1791.390000 2399.820000 1792.290000 ;
      RECT 0.000000 1779.480000 2399.820000 1791.390000 ;
      RECT 0.000000 1778.580000 2398.720000 1779.480000 ;
      RECT 0.000000 1745.320000 2399.820000 1778.580000 ;
      RECT 1.100000 1744.420000 2399.820000 1745.320000 ;
      RECT 0.000000 1731.290000 2399.820000 1744.420000 ;
      RECT 0.000000 1730.390000 2398.720000 1731.290000 ;
      RECT 0.000000 1698.350000 2399.820000 1730.390000 ;
      RECT 1.100000 1697.450000 2399.820000 1698.350000 ;
      RECT 0.000000 1683.100000 2399.820000 1697.450000 ;
      RECT 0.000000 1682.200000 2398.720000 1683.100000 ;
      RECT 0.000000 1650.770000 2399.820000 1682.200000 ;
      RECT 1.100000 1649.870000 2399.820000 1650.770000 ;
      RECT 0.000000 1635.520000 2399.820000 1649.870000 ;
      RECT 0.000000 1634.620000 2398.720000 1635.520000 ;
      RECT 0.000000 1603.800000 2399.820000 1634.620000 ;
      RECT 1.100000 1602.900000 2399.820000 1603.800000 ;
      RECT 0.000000 1587.330000 2399.820000 1602.900000 ;
      RECT 0.000000 1586.430000 2398.720000 1587.330000 ;
      RECT 0.000000 1556.830000 2399.820000 1586.430000 ;
      RECT 1.100000 1555.930000 2399.820000 1556.830000 ;
      RECT 0.000000 1539.140000 2399.820000 1555.930000 ;
      RECT 0.000000 1538.240000 2398.720000 1539.140000 ;
      RECT 0.000000 1509.860000 2399.820000 1538.240000 ;
      RECT 1.100000 1508.960000 2399.820000 1509.860000 ;
      RECT 0.000000 1490.950000 2399.820000 1508.960000 ;
      RECT 0.000000 1490.050000 2398.720000 1490.950000 ;
      RECT 0.000000 1462.280000 2399.820000 1490.050000 ;
      RECT 1.100000 1461.380000 2399.820000 1462.280000 ;
      RECT 0.000000 1443.370000 2399.820000 1461.380000 ;
      RECT 0.000000 1442.470000 2398.720000 1443.370000 ;
      RECT 0.000000 1415.310000 2399.820000 1442.470000 ;
      RECT 1.100000 1414.410000 2399.820000 1415.310000 ;
      RECT 0.000000 1395.180000 2399.820000 1414.410000 ;
      RECT 0.000000 1394.280000 2398.720000 1395.180000 ;
      RECT 0.000000 1368.340000 2399.820000 1394.280000 ;
      RECT 1.100000 1367.440000 2399.820000 1368.340000 ;
      RECT 0.000000 1346.990000 2399.820000 1367.440000 ;
      RECT 0.000000 1346.090000 2398.720000 1346.990000 ;
      RECT 0.000000 1320.760000 2399.820000 1346.090000 ;
      RECT 1.100000 1319.860000 2399.820000 1320.760000 ;
      RECT 0.000000 1298.800000 2399.820000 1319.860000 ;
      RECT 0.000000 1297.900000 2398.720000 1298.800000 ;
      RECT 0.000000 1273.790000 2399.820000 1297.900000 ;
      RECT 1.100000 1272.890000 2399.820000 1273.790000 ;
      RECT 0.000000 1251.220000 2399.820000 1272.890000 ;
      RECT 0.000000 1250.320000 2398.720000 1251.220000 ;
      RECT 0.000000 1226.820000 2399.820000 1250.320000 ;
      RECT 1.100000 1225.920000 2399.820000 1226.820000 ;
      RECT 0.000000 1203.030000 2399.820000 1225.920000 ;
      RECT 0.000000 1202.130000 2398.720000 1203.030000 ;
      RECT 0.000000 1179.850000 2399.820000 1202.130000 ;
      RECT 1.100000 1178.950000 2399.820000 1179.850000 ;
      RECT 0.000000 1154.840000 2399.820000 1178.950000 ;
      RECT 0.000000 1153.940000 2398.720000 1154.840000 ;
      RECT 0.000000 1132.270000 2399.820000 1153.940000 ;
      RECT 1.100000 1131.370000 2399.820000 1132.270000 ;
      RECT 0.000000 1106.650000 2399.820000 1131.370000 ;
      RECT 0.000000 1105.750000 2398.720000 1106.650000 ;
      RECT 0.000000 1085.300000 2399.820000 1105.750000 ;
      RECT 1.100000 1084.400000 2399.820000 1085.300000 ;
      RECT 0.000000 1058.460000 2399.820000 1084.400000 ;
      RECT 0.000000 1057.560000 2398.720000 1058.460000 ;
      RECT 0.000000 1038.330000 2399.820000 1057.560000 ;
      RECT 1.100000 1037.430000 2399.820000 1038.330000 ;
      RECT 0.000000 1010.880000 2399.820000 1037.430000 ;
      RECT 0.000000 1009.980000 2398.720000 1010.880000 ;
      RECT 0.000000 990.750000 2399.820000 1009.980000 ;
      RECT 1.100000 989.850000 2399.820000 990.750000 ;
      RECT 0.000000 962.690000 2399.820000 989.850000 ;
      RECT 0.000000 961.790000 2398.720000 962.690000 ;
      RECT 0.000000 943.780000 2399.820000 961.790000 ;
      RECT 1.100000 942.880000 2399.820000 943.780000 ;
      RECT 0.000000 914.500000 2399.820000 942.880000 ;
      RECT 0.000000 913.600000 2398.720000 914.500000 ;
      RECT 0.000000 896.810000 2399.820000 913.600000 ;
      RECT 1.100000 895.910000 2399.820000 896.810000 ;
      RECT 0.000000 866.310000 2399.820000 895.910000 ;
      RECT 0.000000 865.410000 2398.720000 866.310000 ;
      RECT 0.000000 849.840000 2399.820000 865.410000 ;
      RECT 1.100000 848.940000 2399.820000 849.840000 ;
      RECT 0.000000 818.730000 2399.820000 848.940000 ;
      RECT 0.000000 817.830000 2398.720000 818.730000 ;
      RECT 0.000000 802.260000 2399.820000 817.830000 ;
      RECT 1.100000 801.360000 2399.820000 802.260000 ;
      RECT 0.000000 770.540000 2399.820000 801.360000 ;
      RECT 0.000000 769.640000 2398.720000 770.540000 ;
      RECT 0.000000 755.290000 2399.820000 769.640000 ;
      RECT 1.100000 754.390000 2399.820000 755.290000 ;
      RECT 0.000000 722.350000 2399.820000 754.390000 ;
      RECT 0.000000 721.450000 2398.720000 722.350000 ;
      RECT 0.000000 708.320000 2399.820000 721.450000 ;
      RECT 1.100000 707.420000 2399.820000 708.320000 ;
      RECT 0.000000 674.160000 2399.820000 707.420000 ;
      RECT 0.000000 673.260000 2398.720000 674.160000 ;
      RECT 0.000000 660.740000 2399.820000 673.260000 ;
      RECT 1.100000 659.840000 2399.820000 660.740000 ;
      RECT 0.000000 625.970000 2399.820000 659.840000 ;
      RECT 0.000000 625.070000 2398.720000 625.970000 ;
      RECT 0.000000 613.770000 2399.820000 625.070000 ;
      RECT 1.100000 612.870000 2399.820000 613.770000 ;
      RECT 0.000000 578.390000 2399.820000 612.870000 ;
      RECT 0.000000 577.490000 2398.720000 578.390000 ;
      RECT 0.000000 566.800000 2399.820000 577.490000 ;
      RECT 1.100000 565.900000 2399.820000 566.800000 ;
      RECT 0.000000 530.200000 2399.820000 565.900000 ;
      RECT 0.000000 529.300000 2398.720000 530.200000 ;
      RECT 0.000000 519.830000 2399.820000 529.300000 ;
      RECT 1.100000 518.930000 2399.820000 519.830000 ;
      RECT 0.000000 482.010000 2399.820000 518.930000 ;
      RECT 0.000000 481.110000 2398.720000 482.010000 ;
      RECT 0.000000 472.250000 2399.820000 481.110000 ;
      RECT 1.100000 471.350000 2399.820000 472.250000 ;
      RECT 0.000000 433.820000 2399.820000 471.350000 ;
      RECT 0.000000 432.920000 2398.720000 433.820000 ;
      RECT 0.000000 425.280000 2399.820000 432.920000 ;
      RECT 1.100000 424.380000 2399.820000 425.280000 ;
      RECT 0.000000 386.240000 2399.820000 424.380000 ;
      RECT 0.000000 385.340000 2398.720000 386.240000 ;
      RECT 0.000000 378.310000 2399.820000 385.340000 ;
      RECT 1.100000 377.410000 2399.820000 378.310000 ;
      RECT 0.000000 338.050000 2399.820000 377.410000 ;
      RECT 0.000000 337.150000 2398.720000 338.050000 ;
      RECT 0.000000 330.730000 2399.820000 337.150000 ;
      RECT 1.100000 329.830000 2399.820000 330.730000 ;
      RECT 0.000000 289.860000 2399.820000 329.830000 ;
      RECT 0.000000 288.960000 2398.720000 289.860000 ;
      RECT 0.000000 283.760000 2399.820000 288.960000 ;
      RECT 1.100000 282.860000 2399.820000 283.760000 ;
      RECT 0.000000 241.670000 2399.820000 282.860000 ;
      RECT 0.000000 240.770000 2398.720000 241.670000 ;
      RECT 0.000000 236.790000 2399.820000 240.770000 ;
      RECT 1.100000 235.890000 2399.820000 236.790000 ;
      RECT 0.000000 194.090000 2399.820000 235.890000 ;
      RECT 0.000000 193.190000 2398.720000 194.090000 ;
      RECT 0.000000 189.820000 2399.820000 193.190000 ;
      RECT 1.100000 188.920000 2399.820000 189.820000 ;
      RECT 0.000000 145.900000 2399.820000 188.920000 ;
      RECT 0.000000 145.000000 2398.720000 145.900000 ;
      RECT 0.000000 142.240000 2399.820000 145.000000 ;
      RECT 1.100000 141.340000 2399.820000 142.240000 ;
      RECT 0.000000 97.710000 2399.820000 141.340000 ;
      RECT 0.000000 96.810000 2398.720000 97.710000 ;
      RECT 0.000000 95.270000 2399.820000 96.810000 ;
      RECT 1.100000 94.370000 2399.820000 95.270000 ;
      RECT 0.000000 49.520000 2399.820000 94.370000 ;
      RECT 0.000000 48.620000 2398.720000 49.520000 ;
      RECT 0.000000 48.300000 2399.820000 48.620000 ;
      RECT 1.100000 47.400000 2399.820000 48.300000 ;
      RECT 0.000000 12.310000 2399.820000 47.400000 ;
      RECT 0.000000 11.410000 2398.720000 12.310000 ;
      RECT 0.000000 7.430000 2399.820000 11.410000 ;
      RECT 1.100000 6.530000 2399.820000 7.430000 ;
      RECT 0.000000 1.100000 2399.820000 6.530000 ;
      RECT 2398.200000 0.000000 2399.820000 1.100000 ;
      RECT 2394.980000 0.000000 2397.300000 1.100000 ;
      RECT 2389.920000 0.000000 2394.080000 1.100000 ;
      RECT 2384.860000 0.000000 2389.020000 1.100000 ;
      RECT 2380.260000 0.000000 2383.960000 1.100000 ;
      RECT 2375.200000 0.000000 2379.360000 1.100000 ;
      RECT 2370.600000 0.000000 2374.300000 1.100000 ;
      RECT 2365.540000 0.000000 2369.700000 1.100000 ;
      RECT 2360.940000 0.000000 2364.640000 1.100000 ;
      RECT 2355.880000 0.000000 2360.040000 1.100000 ;
      RECT 2350.820000 0.000000 2354.980000 1.100000 ;
      RECT 2346.220000 0.000000 2349.920000 1.100000 ;
      RECT 2341.160000 0.000000 2345.320000 1.100000 ;
      RECT 2336.560000 0.000000 2340.260000 1.100000 ;
      RECT 2331.500000 0.000000 2335.660000 1.100000 ;
      RECT 2326.440000 0.000000 2330.600000 1.100000 ;
      RECT 2321.840000 0.000000 2325.540000 1.100000 ;
      RECT 2316.780000 0.000000 2320.940000 1.100000 ;
      RECT 2312.180000 0.000000 2315.880000 1.100000 ;
      RECT 2307.120000 0.000000 2311.280000 1.100000 ;
      RECT 2302.520000 0.000000 2306.220000 1.100000 ;
      RECT 2297.460000 0.000000 2301.620000 1.100000 ;
      RECT 2292.400000 0.000000 2296.560000 1.100000 ;
      RECT 2287.800000 0.000000 2291.500000 1.100000 ;
      RECT 2282.740000 0.000000 2286.900000 1.100000 ;
      RECT 2278.140000 0.000000 2281.840000 1.100000 ;
      RECT 2273.080000 0.000000 2277.240000 1.100000 ;
      RECT 2268.020000 0.000000 2272.180000 1.100000 ;
      RECT 2263.420000 0.000000 2267.120000 1.100000 ;
      RECT 2258.360000 0.000000 2262.520000 1.100000 ;
      RECT 2253.760000 0.000000 2257.460000 1.100000 ;
      RECT 2248.700000 0.000000 2252.860000 1.100000 ;
      RECT 2244.100000 0.000000 2247.800000 1.100000 ;
      RECT 2239.040000 0.000000 2243.200000 1.100000 ;
      RECT 2233.980000 0.000000 2238.140000 1.100000 ;
      RECT 2229.380000 0.000000 2233.080000 1.100000 ;
      RECT 2224.320000 0.000000 2228.480000 1.100000 ;
      RECT 2219.720000 0.000000 2223.420000 1.100000 ;
      RECT 2214.660000 0.000000 2218.820000 1.100000 ;
      RECT 2210.060000 0.000000 2213.760000 1.100000 ;
      RECT 2205.000000 0.000000 2209.160000 1.100000 ;
      RECT 2199.940000 0.000000 2204.100000 1.100000 ;
      RECT 2195.340000 0.000000 2199.040000 1.100000 ;
      RECT 2190.280000 0.000000 2194.440000 1.100000 ;
      RECT 2185.680000 0.000000 2189.380000 1.100000 ;
      RECT 2180.620000 0.000000 2184.780000 1.100000 ;
      RECT 2175.560000 0.000000 2179.720000 1.100000 ;
      RECT 2170.960000 0.000000 2174.660000 1.100000 ;
      RECT 2165.900000 0.000000 2170.060000 1.100000 ;
      RECT 2161.300000 0.000000 2165.000000 1.100000 ;
      RECT 2156.240000 0.000000 2160.400000 1.100000 ;
      RECT 2151.640000 0.000000 2155.340000 1.100000 ;
      RECT 2146.580000 0.000000 2150.740000 1.100000 ;
      RECT 2141.520000 0.000000 2145.680000 1.100000 ;
      RECT 2136.920000 0.000000 2140.620000 1.100000 ;
      RECT 2131.860000 0.000000 2136.020000 1.100000 ;
      RECT 2127.260000 0.000000 2130.960000 1.100000 ;
      RECT 2122.200000 0.000000 2126.360000 1.100000 ;
      RECT 2117.140000 0.000000 2121.300000 1.100000 ;
      RECT 2112.540000 0.000000 2116.240000 1.100000 ;
      RECT 2107.480000 0.000000 2111.640000 1.100000 ;
      RECT 2102.880000 0.000000 2106.580000 1.100000 ;
      RECT 2097.820000 0.000000 2101.980000 1.100000 ;
      RECT 2093.220000 0.000000 2096.920000 1.100000 ;
      RECT 2088.160000 0.000000 2092.320000 1.100000 ;
      RECT 2083.100000 0.000000 2087.260000 1.100000 ;
      RECT 2078.500000 0.000000 2082.200000 1.100000 ;
      RECT 2073.440000 0.000000 2077.600000 1.100000 ;
      RECT 2068.840000 0.000000 2072.540000 1.100000 ;
      RECT 2063.780000 0.000000 2067.940000 1.100000 ;
      RECT 2059.180000 0.000000 2062.880000 1.100000 ;
      RECT 2054.120000 0.000000 2058.280000 1.100000 ;
      RECT 2049.060000 0.000000 2053.220000 1.100000 ;
      RECT 2044.460000 0.000000 2048.160000 1.100000 ;
      RECT 2039.400000 0.000000 2043.560000 1.100000 ;
      RECT 2034.800000 0.000000 2038.500000 1.100000 ;
      RECT 2029.740000 0.000000 2033.900000 1.100000 ;
      RECT 2024.680000 0.000000 2028.840000 1.100000 ;
      RECT 2020.080000 0.000000 2023.780000 1.100000 ;
      RECT 2015.020000 0.000000 2019.180000 1.100000 ;
      RECT 2010.420000 0.000000 2014.120000 1.100000 ;
      RECT 2005.360000 0.000000 2009.520000 1.100000 ;
      RECT 2000.760000 0.000000 2004.460000 1.100000 ;
      RECT 1995.700000 0.000000 1999.860000 1.100000 ;
      RECT 1990.640000 0.000000 1994.800000 1.100000 ;
      RECT 1986.040000 0.000000 1989.740000 1.100000 ;
      RECT 1980.980000 0.000000 1985.140000 1.100000 ;
      RECT 1976.380000 0.000000 1980.080000 1.100000 ;
      RECT 1971.320000 0.000000 1975.480000 1.100000 ;
      RECT 1966.720000 0.000000 1970.420000 1.100000 ;
      RECT 1961.660000 0.000000 1965.820000 1.100000 ;
      RECT 1956.600000 0.000000 1960.760000 1.100000 ;
      RECT 1952.000000 0.000000 1955.700000 1.100000 ;
      RECT 1946.940000 0.000000 1951.100000 1.100000 ;
      RECT 1942.340000 0.000000 1946.040000 1.100000 ;
      RECT 1937.280000 0.000000 1941.440000 1.100000 ;
      RECT 1932.220000 0.000000 1936.380000 1.100000 ;
      RECT 1927.620000 0.000000 1931.320000 1.100000 ;
      RECT 1922.560000 0.000000 1926.720000 1.100000 ;
      RECT 1917.960000 0.000000 1921.660000 1.100000 ;
      RECT 1912.900000 0.000000 1917.060000 1.100000 ;
      RECT 1908.300000 0.000000 1912.000000 1.100000 ;
      RECT 1903.240000 0.000000 1907.400000 1.100000 ;
      RECT 1898.180000 0.000000 1902.340000 1.100000 ;
      RECT 1893.580000 0.000000 1897.280000 1.100000 ;
      RECT 1888.520000 0.000000 1892.680000 1.100000 ;
      RECT 1883.920000 0.000000 1887.620000 1.100000 ;
      RECT 1878.860000 0.000000 1883.020000 1.100000 ;
      RECT 1873.800000 0.000000 1877.960000 1.100000 ;
      RECT 1869.200000 0.000000 1872.900000 1.100000 ;
      RECT 1864.140000 0.000000 1868.300000 1.100000 ;
      RECT 1859.540000 0.000000 1863.240000 1.100000 ;
      RECT 1854.480000 0.000000 1858.640000 1.100000 ;
      RECT 1849.880000 0.000000 1853.580000 1.100000 ;
      RECT 1844.820000 0.000000 1848.980000 1.100000 ;
      RECT 1839.760000 0.000000 1843.920000 1.100000 ;
      RECT 1835.160000 0.000000 1838.860000 1.100000 ;
      RECT 1830.100000 0.000000 1834.260000 1.100000 ;
      RECT 1825.500000 0.000000 1829.200000 1.100000 ;
      RECT 1820.440000 0.000000 1824.600000 1.100000 ;
      RECT 1815.840000 0.000000 1819.540000 1.100000 ;
      RECT 1810.780000 0.000000 1814.940000 1.100000 ;
      RECT 1805.720000 0.000000 1809.880000 1.100000 ;
      RECT 1801.120000 0.000000 1804.820000 1.100000 ;
      RECT 1796.060000 0.000000 1800.220000 1.100000 ;
      RECT 1791.460000 0.000000 1795.160000 1.100000 ;
      RECT 1786.400000 0.000000 1790.560000 1.100000 ;
      RECT 1781.340000 0.000000 1785.500000 1.100000 ;
      RECT 1776.740000 0.000000 1780.440000 1.100000 ;
      RECT 1771.680000 0.000000 1775.840000 1.100000 ;
      RECT 1767.080000 0.000000 1770.780000 1.100000 ;
      RECT 1762.020000 0.000000 1766.180000 1.100000 ;
      RECT 1757.420000 0.000000 1761.120000 1.100000 ;
      RECT 1752.360000 0.000000 1756.520000 1.100000 ;
      RECT 1747.300000 0.000000 1751.460000 1.100000 ;
      RECT 1742.700000 0.000000 1746.400000 1.100000 ;
      RECT 1737.640000 0.000000 1741.800000 1.100000 ;
      RECT 1733.040000 0.000000 1736.740000 1.100000 ;
      RECT 1727.980000 0.000000 1732.140000 1.100000 ;
      RECT 1722.920000 0.000000 1727.080000 1.100000 ;
      RECT 1718.320000 0.000000 1722.020000 1.100000 ;
      RECT 1713.260000 0.000000 1717.420000 1.100000 ;
      RECT 1708.660000 0.000000 1712.360000 1.100000 ;
      RECT 1703.600000 0.000000 1707.760000 1.100000 ;
      RECT 1699.000000 0.000000 1702.700000 1.100000 ;
      RECT 1693.940000 0.000000 1698.100000 1.100000 ;
      RECT 1688.880000 0.000000 1693.040000 1.100000 ;
      RECT 1684.280000 0.000000 1687.980000 1.100000 ;
      RECT 1679.220000 0.000000 1683.380000 1.100000 ;
      RECT 1674.620000 0.000000 1678.320000 1.100000 ;
      RECT 1669.560000 0.000000 1673.720000 1.100000 ;
      RECT 1664.960000 0.000000 1668.660000 1.100000 ;
      RECT 1659.900000 0.000000 1664.060000 1.100000 ;
      RECT 1654.840000 0.000000 1659.000000 1.100000 ;
      RECT 1650.240000 0.000000 1653.940000 1.100000 ;
      RECT 1645.180000 0.000000 1649.340000 1.100000 ;
      RECT 1640.580000 0.000000 1644.280000 1.100000 ;
      RECT 1635.520000 0.000000 1639.680000 1.100000 ;
      RECT 1630.460000 0.000000 1634.620000 1.100000 ;
      RECT 1625.860000 0.000000 1629.560000 1.100000 ;
      RECT 1620.800000 0.000000 1624.960000 1.100000 ;
      RECT 1616.200000 0.000000 1619.900000 1.100000 ;
      RECT 1611.140000 0.000000 1615.300000 1.100000 ;
      RECT 1606.540000 0.000000 1610.240000 1.100000 ;
      RECT 1601.480000 0.000000 1605.640000 1.100000 ;
      RECT 1596.420000 0.000000 1600.580000 1.100000 ;
      RECT 1591.820000 0.000000 1595.520000 1.100000 ;
      RECT 1586.760000 0.000000 1590.920000 1.100000 ;
      RECT 1582.160000 0.000000 1585.860000 1.100000 ;
      RECT 1577.100000 0.000000 1581.260000 1.100000 ;
      RECT 1572.040000 0.000000 1576.200000 1.100000 ;
      RECT 1567.440000 0.000000 1571.140000 1.100000 ;
      RECT 1562.380000 0.000000 1566.540000 1.100000 ;
      RECT 1557.780000 0.000000 1561.480000 1.100000 ;
      RECT 1552.720000 0.000000 1556.880000 1.100000 ;
      RECT 1548.120000 0.000000 1551.820000 1.100000 ;
      RECT 1543.060000 0.000000 1547.220000 1.100000 ;
      RECT 1538.000000 0.000000 1542.160000 1.100000 ;
      RECT 1533.400000 0.000000 1537.100000 1.100000 ;
      RECT 1528.340000 0.000000 1532.500000 1.100000 ;
      RECT 1523.740000 0.000000 1527.440000 1.100000 ;
      RECT 1518.680000 0.000000 1522.840000 1.100000 ;
      RECT 1514.080000 0.000000 1517.780000 1.100000 ;
      RECT 1509.020000 0.000000 1513.180000 1.100000 ;
      RECT 1503.960000 0.000000 1508.120000 1.100000 ;
      RECT 1499.360000 0.000000 1503.060000 1.100000 ;
      RECT 1494.300000 0.000000 1498.460000 1.100000 ;
      RECT 1489.700000 0.000000 1493.400000 1.100000 ;
      RECT 1484.640000 0.000000 1488.800000 1.100000 ;
      RECT 1479.580000 0.000000 1483.740000 1.100000 ;
      RECT 1474.980000 0.000000 1478.680000 1.100000 ;
      RECT 1469.920000 0.000000 1474.080000 1.100000 ;
      RECT 1465.320000 0.000000 1469.020000 1.100000 ;
      RECT 1460.260000 0.000000 1464.420000 1.100000 ;
      RECT 1455.660000 0.000000 1459.360000 1.100000 ;
      RECT 1450.600000 0.000000 1454.760000 1.100000 ;
      RECT 1445.540000 0.000000 1449.700000 1.100000 ;
      RECT 1440.940000 0.000000 1444.640000 1.100000 ;
      RECT 1435.880000 0.000000 1440.040000 1.100000 ;
      RECT 1431.280000 0.000000 1434.980000 1.100000 ;
      RECT 1426.220000 0.000000 1430.380000 1.100000 ;
      RECT 1421.160000 0.000000 1425.320000 1.100000 ;
      RECT 1416.560000 0.000000 1420.260000 1.100000 ;
      RECT 1411.500000 0.000000 1415.660000 1.100000 ;
      RECT 1406.900000 0.000000 1410.600000 1.100000 ;
      RECT 1401.840000 0.000000 1406.000000 1.100000 ;
      RECT 1397.240000 0.000000 1400.940000 1.100000 ;
      RECT 1392.180000 0.000000 1396.340000 1.100000 ;
      RECT 1387.120000 0.000000 1391.280000 1.100000 ;
      RECT 1382.520000 0.000000 1386.220000 1.100000 ;
      RECT 1377.460000 0.000000 1381.620000 1.100000 ;
      RECT 1372.860000 0.000000 1376.560000 1.100000 ;
      RECT 1367.800000 0.000000 1371.960000 1.100000 ;
      RECT 1363.200000 0.000000 1366.900000 1.100000 ;
      RECT 1358.140000 0.000000 1362.300000 1.100000 ;
      RECT 1353.080000 0.000000 1357.240000 1.100000 ;
      RECT 1348.480000 0.000000 1352.180000 1.100000 ;
      RECT 1343.420000 0.000000 1347.580000 1.100000 ;
      RECT 1338.820000 0.000000 1342.520000 1.100000 ;
      RECT 1333.760000 0.000000 1337.920000 1.100000 ;
      RECT 1328.700000 0.000000 1332.860000 1.100000 ;
      RECT 1324.100000 0.000000 1327.800000 1.100000 ;
      RECT 1319.040000 0.000000 1323.200000 1.100000 ;
      RECT 1314.440000 0.000000 1318.140000 1.100000 ;
      RECT 1309.380000 0.000000 1313.540000 1.100000 ;
      RECT 1304.780000 0.000000 1308.480000 1.100000 ;
      RECT 1299.720000 0.000000 1303.880000 1.100000 ;
      RECT 1294.660000 0.000000 1298.820000 1.100000 ;
      RECT 1290.060000 0.000000 1293.760000 1.100000 ;
      RECT 1285.000000 0.000000 1289.160000 1.100000 ;
      RECT 1280.400000 0.000000 1284.100000 1.100000 ;
      RECT 1275.340000 0.000000 1279.500000 1.100000 ;
      RECT 1270.280000 0.000000 1274.440000 1.100000 ;
      RECT 1265.680000 0.000000 1269.380000 1.100000 ;
      RECT 1260.620000 0.000000 1264.780000 1.100000 ;
      RECT 1256.020000 0.000000 1259.720000 1.100000 ;
      RECT 1250.960000 0.000000 1255.120000 1.100000 ;
      RECT 1246.360000 0.000000 1250.060000 1.100000 ;
      RECT 1241.300000 0.000000 1245.460000 1.100000 ;
      RECT 1236.240000 0.000000 1240.400000 1.100000 ;
      RECT 1231.640000 0.000000 1235.340000 1.100000 ;
      RECT 1226.580000 0.000000 1230.740000 1.100000 ;
      RECT 1221.980000 0.000000 1225.680000 1.100000 ;
      RECT 1216.920000 0.000000 1221.080000 1.100000 ;
      RECT 1212.320000 0.000000 1216.020000 1.100000 ;
      RECT 1207.260000 0.000000 1211.420000 1.100000 ;
      RECT 1202.200000 0.000000 1206.360000 1.100000 ;
      RECT 1197.600000 0.000000 1201.300000 1.100000 ;
      RECT 1192.540000 0.000000 1196.700000 1.100000 ;
      RECT 1187.940000 0.000000 1191.640000 1.100000 ;
      RECT 1182.880000 0.000000 1187.040000 1.100000 ;
      RECT 1177.820000 0.000000 1181.980000 1.100000 ;
      RECT 1173.220000 0.000000 1176.920000 1.100000 ;
      RECT 1168.160000 0.000000 1172.320000 1.100000 ;
      RECT 1163.560000 0.000000 1167.260000 1.100000 ;
      RECT 1158.500000 0.000000 1162.660000 1.100000 ;
      RECT 1153.900000 0.000000 1157.600000 1.100000 ;
      RECT 1148.840000 0.000000 1153.000000 1.100000 ;
      RECT 1143.780000 0.000000 1147.940000 1.100000 ;
      RECT 1139.180000 0.000000 1142.880000 1.100000 ;
      RECT 1134.120000 0.000000 1138.280000 1.100000 ;
      RECT 1129.520000 0.000000 1133.220000 1.100000 ;
      RECT 1124.460000 0.000000 1128.620000 1.100000 ;
      RECT 1119.860000 0.000000 1123.560000 1.100000 ;
      RECT 1114.800000 0.000000 1118.960000 1.100000 ;
      RECT 1109.740000 0.000000 1113.900000 1.100000 ;
      RECT 1105.140000 0.000000 1108.840000 1.100000 ;
      RECT 1100.080000 0.000000 1104.240000 1.100000 ;
      RECT 1095.480000 0.000000 1099.180000 1.100000 ;
      RECT 1090.420000 0.000000 1094.580000 1.100000 ;
      RECT 1085.360000 0.000000 1089.520000 1.100000 ;
      RECT 1080.760000 0.000000 1084.460000 1.100000 ;
      RECT 1075.700000 0.000000 1079.860000 1.100000 ;
      RECT 1071.100000 0.000000 1074.800000 1.100000 ;
      RECT 1066.040000 0.000000 1070.200000 1.100000 ;
      RECT 1061.440000 0.000000 1065.140000 1.100000 ;
      RECT 1056.380000 0.000000 1060.540000 1.100000 ;
      RECT 1051.320000 0.000000 1055.480000 1.100000 ;
      RECT 1046.720000 0.000000 1050.420000 1.100000 ;
      RECT 1041.660000 0.000000 1045.820000 1.100000 ;
      RECT 1037.060000 0.000000 1040.760000 1.100000 ;
      RECT 1032.000000 0.000000 1036.160000 1.100000 ;
      RECT 1026.940000 0.000000 1031.100000 1.100000 ;
      RECT 1022.340000 0.000000 1026.040000 1.100000 ;
      RECT 1017.280000 0.000000 1021.440000 1.100000 ;
      RECT 1012.680000 0.000000 1016.380000 1.100000 ;
      RECT 1007.620000 0.000000 1011.780000 1.100000 ;
      RECT 1003.020000 0.000000 1006.720000 1.100000 ;
      RECT 997.960000 0.000000 1002.120000 1.100000 ;
      RECT 992.900000 0.000000 997.060000 1.100000 ;
      RECT 988.300000 0.000000 992.000000 1.100000 ;
      RECT 983.240000 0.000000 987.400000 1.100000 ;
      RECT 978.640000 0.000000 982.340000 1.100000 ;
      RECT 973.580000 0.000000 977.740000 1.100000 ;
      RECT 968.980000 0.000000 972.680000 1.100000 ;
      RECT 963.920000 0.000000 968.080000 1.100000 ;
      RECT 958.860000 0.000000 963.020000 1.100000 ;
      RECT 954.260000 0.000000 957.960000 1.100000 ;
      RECT 949.200000 0.000000 953.360000 1.100000 ;
      RECT 944.600000 0.000000 948.300000 1.100000 ;
      RECT 939.540000 0.000000 943.700000 1.100000 ;
      RECT 934.480000 0.000000 938.640000 1.100000 ;
      RECT 929.880000 0.000000 933.580000 1.100000 ;
      RECT 924.820000 0.000000 928.980000 1.100000 ;
      RECT 920.220000 0.000000 923.920000 1.100000 ;
      RECT 915.160000 0.000000 919.320000 1.100000 ;
      RECT 910.560000 0.000000 914.260000 1.100000 ;
      RECT 905.500000 0.000000 909.660000 1.100000 ;
      RECT 900.440000 0.000000 904.600000 1.100000 ;
      RECT 895.840000 0.000000 899.540000 1.100000 ;
      RECT 890.780000 0.000000 894.940000 1.100000 ;
      RECT 886.180000 0.000000 889.880000 1.100000 ;
      RECT 881.120000 0.000000 885.280000 1.100000 ;
      RECT 876.060000 0.000000 880.220000 1.100000 ;
      RECT 871.460000 0.000000 875.160000 1.100000 ;
      RECT 866.400000 0.000000 870.560000 1.100000 ;
      RECT 861.800000 0.000000 865.500000 1.100000 ;
      RECT 856.740000 0.000000 860.900000 1.100000 ;
      RECT 852.140000 0.000000 855.840000 1.100000 ;
      RECT 847.080000 0.000000 851.240000 1.100000 ;
      RECT 842.020000 0.000000 846.180000 1.100000 ;
      RECT 837.420000 0.000000 841.120000 1.100000 ;
      RECT 832.360000 0.000000 836.520000 1.100000 ;
      RECT 827.760000 0.000000 831.460000 1.100000 ;
      RECT 822.700000 0.000000 826.860000 1.100000 ;
      RECT 818.100000 0.000000 821.800000 1.100000 ;
      RECT 813.040000 0.000000 817.200000 1.100000 ;
      RECT 807.980000 0.000000 812.140000 1.100000 ;
      RECT 803.380000 0.000000 807.080000 1.100000 ;
      RECT 798.320000 0.000000 802.480000 1.100000 ;
      RECT 793.720000 0.000000 797.420000 1.100000 ;
      RECT 788.660000 0.000000 792.820000 1.100000 ;
      RECT 783.600000 0.000000 787.760000 1.100000 ;
      RECT 779.000000 0.000000 782.700000 1.100000 ;
      RECT 773.940000 0.000000 778.100000 1.100000 ;
      RECT 769.340000 0.000000 773.040000 1.100000 ;
      RECT 764.280000 0.000000 768.440000 1.100000 ;
      RECT 759.680000 0.000000 763.380000 1.100000 ;
      RECT 754.620000 0.000000 758.780000 1.100000 ;
      RECT 749.560000 0.000000 753.720000 1.100000 ;
      RECT 744.960000 0.000000 748.660000 1.100000 ;
      RECT 739.900000 0.000000 744.060000 1.100000 ;
      RECT 735.300000 0.000000 739.000000 1.100000 ;
      RECT 730.240000 0.000000 734.400000 1.100000 ;
      RECT 725.180000 0.000000 729.340000 1.100000 ;
      RECT 720.580000 0.000000 724.280000 1.100000 ;
      RECT 715.520000 0.000000 719.680000 1.100000 ;
      RECT 710.920000 0.000000 714.620000 1.100000 ;
      RECT 705.860000 0.000000 710.020000 1.100000 ;
      RECT 701.260000 0.000000 704.960000 1.100000 ;
      RECT 696.200000 0.000000 700.360000 1.100000 ;
      RECT 691.140000 0.000000 695.300000 1.100000 ;
      RECT 686.540000 0.000000 690.240000 1.100000 ;
      RECT 681.480000 0.000000 685.640000 1.100000 ;
      RECT 676.880000 0.000000 680.580000 1.100000 ;
      RECT 671.820000 0.000000 675.980000 1.100000 ;
      RECT 667.220000 0.000000 670.920000 1.100000 ;
      RECT 662.160000 0.000000 666.320000 1.100000 ;
      RECT 657.100000 0.000000 661.260000 1.100000 ;
      RECT 652.500000 0.000000 656.200000 1.100000 ;
      RECT 647.440000 0.000000 651.600000 1.100000 ;
      RECT 642.840000 0.000000 646.540000 1.100000 ;
      RECT 637.780000 0.000000 641.940000 1.100000 ;
      RECT 632.720000 0.000000 636.880000 1.100000 ;
      RECT 628.120000 0.000000 631.820000 1.100000 ;
      RECT 623.060000 0.000000 627.220000 1.100000 ;
      RECT 618.460000 0.000000 622.160000 1.100000 ;
      RECT 613.400000 0.000000 617.560000 1.100000 ;
      RECT 608.800000 0.000000 612.500000 1.100000 ;
      RECT 603.740000 0.000000 607.900000 1.100000 ;
      RECT 598.680000 0.000000 602.840000 1.100000 ;
      RECT 594.080000 0.000000 597.780000 1.100000 ;
      RECT 589.020000 0.000000 593.180000 1.100000 ;
      RECT 584.420000 0.000000 588.120000 1.100000 ;
      RECT 579.360000 0.000000 583.520000 1.100000 ;
      RECT 574.300000 0.000000 578.460000 1.100000 ;
      RECT 569.700000 0.000000 573.400000 1.100000 ;
      RECT 564.640000 0.000000 568.800000 1.100000 ;
      RECT 560.040000 0.000000 563.740000 1.100000 ;
      RECT 554.980000 0.000000 559.140000 1.100000 ;
      RECT 550.380000 0.000000 554.080000 1.100000 ;
      RECT 545.320000 0.000000 549.480000 1.100000 ;
      RECT 540.260000 0.000000 544.420000 1.100000 ;
      RECT 535.660000 0.000000 539.360000 1.100000 ;
      RECT 530.600000 0.000000 534.760000 1.100000 ;
      RECT 526.000000 0.000000 529.700000 1.100000 ;
      RECT 520.940000 0.000000 525.100000 1.100000 ;
      RECT 516.340000 0.000000 520.040000 1.100000 ;
      RECT 511.280000 0.000000 515.440000 1.100000 ;
      RECT 506.220000 0.000000 510.380000 1.100000 ;
      RECT 501.620000 0.000000 505.320000 1.100000 ;
      RECT 496.560000 0.000000 500.720000 1.100000 ;
      RECT 491.960000 0.000000 495.660000 1.100000 ;
      RECT 486.900000 0.000000 491.060000 1.100000 ;
      RECT 481.840000 0.000000 486.000000 1.100000 ;
      RECT 477.240000 0.000000 480.940000 1.100000 ;
      RECT 472.180000 0.000000 476.340000 1.100000 ;
      RECT 467.580000 0.000000 471.280000 1.100000 ;
      RECT 462.520000 0.000000 466.680000 1.100000 ;
      RECT 457.920000 0.000000 461.620000 1.100000 ;
      RECT 452.860000 0.000000 457.020000 1.100000 ;
      RECT 447.800000 0.000000 451.960000 1.100000 ;
      RECT 443.200000 0.000000 446.900000 1.100000 ;
      RECT 438.140000 0.000000 442.300000 1.100000 ;
      RECT 433.540000 0.000000 437.240000 1.100000 ;
      RECT 428.480000 0.000000 432.640000 1.100000 ;
      RECT 423.880000 0.000000 427.580000 1.100000 ;
      RECT 418.820000 0.000000 422.980000 1.100000 ;
      RECT 413.760000 0.000000 417.920000 1.100000 ;
      RECT 409.160000 0.000000 412.860000 1.100000 ;
      RECT 404.100000 0.000000 408.260000 1.100000 ;
      RECT 399.500000 0.000000 403.200000 1.100000 ;
      RECT 394.440000 0.000000 398.600000 1.100000 ;
      RECT 389.380000 0.000000 393.540000 1.100000 ;
      RECT 384.780000 0.000000 388.480000 1.100000 ;
      RECT 379.720000 0.000000 383.880000 1.100000 ;
      RECT 375.120000 0.000000 378.820000 1.100000 ;
      RECT 370.060000 0.000000 374.220000 1.100000 ;
      RECT 365.460000 0.000000 369.160000 1.100000 ;
      RECT 360.400000 0.000000 364.560000 1.100000 ;
      RECT 355.340000 0.000000 359.500000 1.100000 ;
      RECT 350.740000 0.000000 354.440000 1.100000 ;
      RECT 345.680000 0.000000 349.840000 1.100000 ;
      RECT 341.080000 0.000000 344.780000 1.100000 ;
      RECT 336.020000 0.000000 340.180000 1.100000 ;
      RECT 330.960000 0.000000 335.120000 1.100000 ;
      RECT 326.360000 0.000000 330.060000 1.100000 ;
      RECT 321.300000 0.000000 325.460000 1.100000 ;
      RECT 316.700000 0.000000 320.400000 1.100000 ;
      RECT 311.640000 0.000000 315.800000 1.100000 ;
      RECT 307.040000 0.000000 310.740000 1.100000 ;
      RECT 301.980000 0.000000 306.140000 1.100000 ;
      RECT 296.920000 0.000000 301.080000 1.100000 ;
      RECT 292.320000 0.000000 296.020000 1.100000 ;
      RECT 287.260000 0.000000 291.420000 1.100000 ;
      RECT 282.660000 0.000000 286.360000 1.100000 ;
      RECT 277.600000 0.000000 281.760000 1.100000 ;
      RECT 273.000000 0.000000 276.700000 1.100000 ;
      RECT 267.940000 0.000000 272.100000 1.100000 ;
      RECT 262.880000 0.000000 267.040000 1.100000 ;
      RECT 258.280000 0.000000 261.980000 1.100000 ;
      RECT 253.220000 0.000000 257.380000 1.100000 ;
      RECT 248.620000 0.000000 252.320000 1.100000 ;
      RECT 243.560000 0.000000 247.720000 1.100000 ;
      RECT 238.500000 0.000000 242.660000 1.100000 ;
      RECT 233.900000 0.000000 237.600000 1.100000 ;
      RECT 228.840000 0.000000 233.000000 1.100000 ;
      RECT 224.240000 0.000000 227.940000 1.100000 ;
      RECT 219.180000 0.000000 223.340000 1.100000 ;
      RECT 214.580000 0.000000 218.280000 1.100000 ;
      RECT 209.520000 0.000000 213.680000 1.100000 ;
      RECT 204.460000 0.000000 208.620000 1.100000 ;
      RECT 199.860000 0.000000 203.560000 1.100000 ;
      RECT 194.800000 0.000000 198.960000 1.100000 ;
      RECT 190.200000 0.000000 193.900000 1.100000 ;
      RECT 185.140000 0.000000 189.300000 1.100000 ;
      RECT 180.080000 0.000000 184.240000 1.100000 ;
      RECT 175.480000 0.000000 179.180000 1.100000 ;
      RECT 170.420000 0.000000 174.580000 1.100000 ;
      RECT 165.820000 0.000000 169.520000 1.100000 ;
      RECT 160.760000 0.000000 164.920000 1.100000 ;
      RECT 156.160000 0.000000 159.860000 1.100000 ;
      RECT 151.100000 0.000000 155.260000 1.100000 ;
      RECT 146.040000 0.000000 150.200000 1.100000 ;
      RECT 141.440000 0.000000 145.140000 1.100000 ;
      RECT 136.380000 0.000000 140.540000 1.100000 ;
      RECT 131.780000 0.000000 135.480000 1.100000 ;
      RECT 126.720000 0.000000 130.880000 1.100000 ;
      RECT 122.120000 0.000000 125.820000 1.100000 ;
      RECT 117.060000 0.000000 121.220000 1.100000 ;
      RECT 112.000000 0.000000 116.160000 1.100000 ;
      RECT 107.400000 0.000000 111.100000 1.100000 ;
      RECT 102.340000 0.000000 106.500000 1.100000 ;
      RECT 97.740000 0.000000 101.440000 1.100000 ;
      RECT 92.680000 0.000000 96.840000 1.100000 ;
      RECT 87.620000 0.000000 91.780000 1.100000 ;
      RECT 83.020000 0.000000 86.720000 1.100000 ;
      RECT 77.960000 0.000000 82.120000 1.100000 ;
      RECT 73.360000 0.000000 77.060000 1.100000 ;
      RECT 68.300000 0.000000 72.460000 1.100000 ;
      RECT 63.700000 0.000000 67.400000 1.100000 ;
      RECT 58.640000 0.000000 62.800000 1.100000 ;
      RECT 53.580000 0.000000 57.740000 1.100000 ;
      RECT 48.980000 0.000000 52.680000 1.100000 ;
      RECT 43.920000 0.000000 48.080000 1.100000 ;
      RECT 39.320000 0.000000 43.020000 1.100000 ;
      RECT 34.260000 0.000000 38.420000 1.100000 ;
      RECT 29.200000 0.000000 33.360000 1.100000 ;
      RECT 24.600000 0.000000 28.300000 1.100000 ;
      RECT 19.540000 0.000000 23.700000 1.100000 ;
      RECT 14.940000 0.000000 18.640000 1.100000 ;
      RECT 9.880000 0.000000 14.040000 1.100000 ;
      RECT 5.280000 0.000000 8.980000 1.100000 ;
      RECT 2.520000 0.000000 4.380000 1.100000 ;
      RECT 0.000000 0.000000 1.620000 1.100000 ;
    LAYER met4 ;
      RECT 0.000000 2495.280000 2399.820000 2500.020000 ;
      RECT 5.020000 2491.680000 2394.800000 2495.280000 ;
      RECT 5.020000 2411.680000 2391.200000 2491.680000 ;
      RECT 2393.600000 5.960000 2394.800000 2491.680000 ;
      RECT 8.620000 5.960000 2391.200000 2411.680000 ;
      RECT 5.020000 5.960000 6.220000 2411.680000 ;
      RECT 2397.200000 2.360000 2399.820000 2495.280000 ;
      RECT 5.020000 2.360000 2394.800000 5.960000 ;
      RECT 0.000000 2.360000 2.620000 2495.280000 ;
      RECT 0.000000 0.000000 2399.820000 2.360000 ;
    LAYER met5 ;
      RECT 0.000000 0.000000 2399.820000 2500.020000 ;
  END
END azadi_soc_top_caravel

END LIBRARY
