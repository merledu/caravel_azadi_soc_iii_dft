magic
tech sky130A
magscale 1 2
timestamp 1653864141
<< metal1 >>
rect 10318 558900 10324 558952
rect 10376 558940 10382 558952
rect 57422 558940 57428 558952
rect 10376 558912 57428 558940
rect 10376 558900 10382 558912
rect 57422 558900 57428 558912
rect 57480 558900 57486 558952
rect 381906 59780 381912 59832
rect 381964 59820 381970 59832
rect 383286 59820 383292 59832
rect 381964 59792 383292 59820
rect 381964 59780 381970 59792
rect 383286 59780 383292 59792
rect 383344 59780 383350 59832
rect 64782 59712 64788 59764
rect 64840 59752 64846 59764
rect 65886 59752 65892 59764
rect 64840 59724 65892 59752
rect 64840 59712 64846 59724
rect 65886 59712 65892 59724
rect 65944 59712 65950 59764
rect 94498 59712 94504 59764
rect 94556 59752 94562 59764
rect 97074 59752 97080 59764
rect 94556 59724 97080 59752
rect 94556 59712 94562 59724
rect 97074 59712 97080 59724
rect 97132 59712 97138 59764
rect 98822 59712 98828 59764
rect 98880 59752 98886 59764
rect 100938 59752 100944 59764
rect 98880 59724 100944 59752
rect 98880 59712 98886 59724
rect 100938 59712 100944 59724
rect 100996 59712 101002 59764
rect 105538 59712 105544 59764
rect 105596 59752 105602 59764
rect 107746 59752 107752 59764
rect 105596 59724 107752 59752
rect 105596 59712 105602 59724
rect 107746 59712 107752 59724
rect 107804 59712 107810 59764
rect 108482 59712 108488 59764
rect 108540 59752 108546 59764
rect 110690 59752 110696 59764
rect 108540 59724 110696 59752
rect 108540 59712 108546 59724
rect 110690 59712 110696 59724
rect 110748 59712 110754 59764
rect 113818 59712 113824 59764
rect 113876 59752 113882 59764
rect 115566 59752 115572 59764
rect 113876 59724 115572 59752
rect 113876 59712 113882 59724
rect 115566 59712 115572 59724
rect 115624 59712 115630 59764
rect 124858 59712 124864 59764
rect 124916 59752 124922 59764
rect 127250 59752 127256 59764
rect 124916 59724 127256 59752
rect 124916 59712 124922 59724
rect 127250 59712 127256 59724
rect 127308 59712 127314 59764
rect 128998 59712 129004 59764
rect 129056 59752 129062 59764
rect 131114 59752 131120 59764
rect 129056 59724 131120 59752
rect 129056 59712 129062 59724
rect 131114 59712 131120 59724
rect 131172 59712 131178 59764
rect 131758 59712 131764 59764
rect 131816 59752 131822 59764
rect 134058 59752 134064 59764
rect 131816 59724 134064 59752
rect 131816 59712 131822 59724
rect 134058 59712 134064 59724
rect 134116 59712 134122 59764
rect 135162 59712 135168 59764
rect 135220 59752 135226 59764
rect 137002 59752 137008 59764
rect 135220 59724 137008 59752
rect 135220 59712 135226 59724
rect 137002 59712 137008 59724
rect 137060 59712 137066 59764
rect 141418 59712 141424 59764
rect 141476 59752 141482 59764
rect 143810 59752 143816 59764
rect 141476 59724 143816 59752
rect 141476 59712 141482 59724
rect 143810 59712 143816 59724
rect 143868 59712 143874 59764
rect 145558 59712 145564 59764
rect 145616 59752 145622 59764
rect 147674 59752 147680 59764
rect 145616 59724 147680 59752
rect 145616 59712 145622 59724
rect 147674 59712 147680 59724
rect 147732 59712 147738 59764
rect 148318 59712 148324 59764
rect 148376 59752 148382 59764
rect 150618 59752 150624 59764
rect 148376 59724 150624 59752
rect 148376 59712 148382 59724
rect 150618 59712 150624 59724
rect 150676 59712 150682 59764
rect 155218 59712 155224 59764
rect 155276 59752 155282 59764
rect 157426 59752 157432 59764
rect 155276 59724 157432 59752
rect 155276 59712 155282 59724
rect 157426 59712 157432 59724
rect 157484 59712 157490 59764
rect 160738 59712 160744 59764
rect 160796 59752 160802 59764
rect 163314 59752 163320 59764
rect 160796 59724 163320 59752
rect 160796 59712 160802 59724
rect 163314 59712 163320 59724
rect 163372 59712 163378 59764
rect 179322 59712 179328 59764
rect 179380 59752 179386 59764
rect 180794 59752 180800 59764
rect 179380 59724 180800 59752
rect 179380 59712 179386 59724
rect 180794 59712 180800 59724
rect 180852 59712 180858 59764
rect 184750 59712 184756 59764
rect 184808 59752 184814 59764
rect 186590 59752 186596 59764
rect 184808 59724 186596 59752
rect 184808 59712 184814 59724
rect 186590 59712 186596 59724
rect 186648 59712 186654 59764
rect 193214 59712 193220 59764
rect 193272 59752 193278 59764
rect 193766 59752 193772 59764
rect 193272 59724 193772 59752
rect 193272 59712 193278 59724
rect 193766 59712 193772 59724
rect 193824 59712 193830 59764
rect 202782 59712 202788 59764
rect 202840 59752 202846 59764
rect 204162 59752 204168 59764
rect 202840 59724 204168 59752
rect 202840 59712 202846 59724
rect 204162 59712 204168 59724
rect 204220 59712 204226 59764
rect 208026 59712 208032 59764
rect 208084 59752 208090 59764
rect 209682 59752 209688 59764
rect 208084 59724 209688 59752
rect 208084 59712 208090 59724
rect 209682 59712 209688 59724
rect 209740 59712 209746 59764
rect 210970 59712 210976 59764
rect 211028 59752 211034 59764
rect 212902 59752 212908 59764
rect 211028 59724 212908 59752
rect 211028 59712 211034 59724
rect 212902 59712 212908 59724
rect 212960 59712 212966 59764
rect 220538 59712 220544 59764
rect 220596 59752 220602 59764
rect 222654 59752 222660 59764
rect 220596 59724 222660 59752
rect 220596 59712 220602 59724
rect 222654 59712 222660 59724
rect 222712 59712 222718 59764
rect 227530 59712 227536 59764
rect 227588 59752 227594 59764
rect 229462 59752 229468 59764
rect 227588 59724 229468 59752
rect 227588 59712 227594 59724
rect 229462 59712 229468 59724
rect 229520 59712 229526 59764
rect 230106 59712 230112 59764
rect 230164 59752 230170 59764
rect 232406 59752 232412 59764
rect 230164 59724 232412 59752
rect 230164 59712 230170 59724
rect 232406 59712 232412 59724
rect 232464 59712 232470 59764
rect 238662 59712 238668 59764
rect 238720 59752 238726 59764
rect 240134 59752 240140 59764
rect 238720 59724 240140 59752
rect 238720 59712 238726 59724
rect 240134 59712 240140 59724
rect 240192 59712 240198 59764
rect 246666 59712 246672 59764
rect 246724 59752 246730 59764
rect 248966 59752 248972 59764
rect 246724 59724 248972 59752
rect 246724 59712 246730 59724
rect 248966 59712 248972 59724
rect 249024 59712 249030 59764
rect 250990 59712 250996 59764
rect 251048 59752 251054 59764
rect 252830 59752 252836 59764
rect 251048 59724 252836 59752
rect 251048 59712 251054 59724
rect 252830 59712 252836 59724
rect 252888 59712 252894 59764
rect 271782 59712 271788 59764
rect 271840 59752 271846 59764
rect 273254 59752 273260 59764
rect 271840 59724 273260 59752
rect 271840 59712 271846 59724
rect 273254 59712 273260 59724
rect 273312 59712 273318 59764
rect 278682 59712 278688 59764
rect 278740 59752 278746 59764
rect 280062 59752 280068 59764
rect 278740 59724 280068 59752
rect 278740 59712 278746 59724
rect 280062 59712 280068 59724
rect 280120 59712 280126 59764
rect 287698 59712 287704 59764
rect 287756 59752 287762 59764
rect 289814 59752 289820 59764
rect 287756 59724 289820 59752
rect 287756 59712 287762 59724
rect 289814 59712 289820 59724
rect 289872 59712 289878 59764
rect 290458 59712 290464 59764
rect 290516 59752 290522 59764
rect 292758 59752 292764 59764
rect 290516 59724 292764 59752
rect 290516 59712 290522 59724
rect 292758 59712 292764 59724
rect 292816 59712 292822 59764
rect 315758 59712 315764 59764
rect 315816 59752 315822 59764
rect 317598 59752 317604 59764
rect 315816 59724 317604 59752
rect 315816 59712 315822 59724
rect 317598 59712 317604 59724
rect 317656 59712 317662 59764
rect 322566 59712 322572 59764
rect 322624 59752 322630 59764
rect 324682 59752 324688 59764
rect 322624 59724 324688 59752
rect 322624 59712 322630 59724
rect 324682 59712 324688 59724
rect 324740 59712 324746 59764
rect 334342 59712 334348 59764
rect 334400 59752 334406 59764
rect 335262 59752 335268 59764
rect 334400 59724 335268 59752
rect 334400 59712 334406 59724
rect 335262 59712 335268 59724
rect 335320 59712 335326 59764
rect 339126 59712 339132 59764
rect 339184 59752 339190 59764
rect 340966 59752 340972 59764
rect 339184 59724 340972 59752
rect 339184 59712 339190 59724
rect 340966 59712 340972 59724
rect 341024 59712 341030 59764
rect 355594 59712 355600 59764
rect 355652 59752 355658 59764
rect 358262 59752 358268 59764
rect 355652 59724 358268 59752
rect 355652 59712 355658 59724
rect 358262 59712 358268 59724
rect 358320 59712 358326 59764
rect 365346 59712 365352 59764
rect 365404 59752 365410 59764
rect 367738 59752 367744 59764
rect 365404 59724 367744 59752
rect 365404 59712 365410 59724
rect 367738 59712 367744 59724
rect 367796 59712 367802 59764
rect 369302 59712 369308 59764
rect 369360 59752 369366 59764
rect 371970 59752 371976 59764
rect 369360 59724 371976 59752
rect 369360 59712 369366 59724
rect 371970 59712 371976 59724
rect 372028 59712 372034 59764
rect 385954 59712 385960 59764
rect 386012 59752 386018 59764
rect 388622 59752 388628 59764
rect 386012 59724 388628 59752
rect 386012 59712 386018 59724
rect 388622 59712 388628 59724
rect 388680 59712 388686 59764
rect 388714 59712 388720 59764
rect 388772 59752 388778 59764
rect 391382 59752 391388 59764
rect 388772 59724 391388 59752
rect 388772 59712 388778 59724
rect 391382 59712 391388 59724
rect 391440 59712 391446 59764
rect 391658 59712 391664 59764
rect 391716 59752 391722 59764
rect 394142 59752 394148 59764
rect 391716 59724 394148 59752
rect 391716 59712 391722 59724
rect 394142 59712 394148 59724
rect 394200 59712 394206 59764
rect 395706 59712 395712 59764
rect 395764 59752 395770 59764
rect 398098 59752 398104 59764
rect 395764 59724 398104 59752
rect 395764 59712 395770 59724
rect 398098 59712 398104 59724
rect 398156 59712 398162 59764
rect 398466 59712 398472 59764
rect 398524 59752 398530 59764
rect 401042 59752 401048 59764
rect 398524 59724 401048 59752
rect 398524 59712 398530 59724
rect 401042 59712 401048 59724
rect 401100 59712 401106 59764
rect 402422 59712 402428 59764
rect 402480 59752 402486 59764
rect 405182 59752 405188 59764
rect 402480 59724 405188 59752
rect 402480 59712 402486 59724
rect 405182 59712 405188 59724
rect 405240 59712 405246 59764
rect 405274 59712 405280 59764
rect 405332 59752 405338 59764
rect 407942 59752 407948 59764
rect 405332 59724 407948 59752
rect 405332 59712 405338 59724
rect 407942 59712 407948 59724
rect 408000 59712 408006 59764
rect 410150 59712 410156 59764
rect 410208 59752 410214 59764
rect 411898 59752 411904 59764
rect 410208 59724 411904 59752
rect 410208 59712 410214 59724
rect 411898 59712 411904 59724
rect 411956 59712 411962 59764
rect 413094 59712 413100 59764
rect 413152 59752 413158 59764
rect 414658 59752 414664 59764
rect 413152 59724 414664 59752
rect 413152 59712 413158 59724
rect 414658 59712 414664 59724
rect 414716 59712 414722 59764
rect 438026 59712 438032 59764
rect 438084 59752 438090 59764
rect 438854 59752 438860 59764
rect 438084 59724 438860 59752
rect 438084 59712 438090 59724
rect 438854 59712 438860 59724
rect 438912 59712 438918 59764
rect 456610 59712 456616 59764
rect 456668 59752 456674 59764
rect 457070 59752 457076 59764
rect 456668 59724 457076 59752
rect 456668 59712 456674 59724
rect 457070 59712 457076 59724
rect 457128 59712 457134 59764
rect 461578 59712 461584 59764
rect 461636 59752 461642 59764
rect 462406 59752 462412 59764
rect 461636 59724 462412 59752
rect 461636 59712 461642 59724
rect 462406 59712 462412 59724
rect 462464 59712 462470 59764
rect 470594 59712 470600 59764
rect 470652 59752 470658 59764
rect 471974 59752 471980 59764
rect 470652 59724 471980 59752
rect 470652 59712 470658 59724
rect 471974 59712 471980 59724
rect 472032 59712 472038 59764
rect 474366 59712 474372 59764
rect 474424 59752 474430 59764
rect 476390 59752 476396 59764
rect 474424 59724 476396 59752
rect 474424 59712 474430 59724
rect 476390 59712 476396 59724
rect 476448 59712 476454 59764
rect 480254 59712 480260 59764
rect 480312 59752 480318 59764
rect 481634 59752 481640 59764
rect 480312 59724 481640 59752
rect 480312 59712 480318 59724
rect 481634 59712 481640 59724
rect 481692 59712 481698 59764
rect 495894 59712 495900 59764
rect 495952 59752 495958 59764
rect 496906 59752 496912 59764
rect 495952 59724 496912 59752
rect 495952 59712 495958 59724
rect 496906 59712 496912 59724
rect 496964 59712 496970 59764
rect 500678 59712 500684 59764
rect 500736 59752 500742 59764
rect 502610 59752 502616 59764
rect 500736 59724 502616 59752
rect 500736 59712 500742 59724
rect 502610 59712 502616 59724
rect 502668 59712 502674 59764
rect 503622 59712 503628 59764
rect 503680 59752 503686 59764
rect 505186 59752 505192 59764
rect 503680 59724 505192 59752
rect 503680 59712 503686 59724
rect 505186 59712 505192 59724
rect 505244 59712 505250 59764
rect 517238 59712 517244 59764
rect 517296 59752 517302 59764
rect 519170 59752 519176 59764
rect 517296 59724 519176 59752
rect 517296 59712 517302 59724
rect 519170 59712 519176 59724
rect 519228 59712 519234 59764
rect 522114 59712 522120 59764
rect 522172 59752 522178 59764
rect 523678 59752 523684 59764
rect 522172 59724 523684 59752
rect 522172 59712 522178 59724
rect 523678 59712 523684 59724
rect 523736 59712 523742 59764
rect 524046 59712 524052 59764
rect 524104 59752 524110 59764
rect 526438 59752 526444 59764
rect 524104 59724 526444 59752
rect 524104 59712 524110 59724
rect 526438 59712 526444 59724
rect 526496 59712 526502 59764
rect 526990 59712 526996 59764
rect 527048 59752 527054 59764
rect 529198 59752 529204 59764
rect 527048 59724 529204 59752
rect 527048 59712 527054 59724
rect 529198 59712 529204 59724
rect 529256 59712 529262 59764
rect 530854 59712 530860 59764
rect 530912 59752 530918 59764
rect 533522 59752 533528 59764
rect 530912 59724 533528 59752
rect 530912 59712 530918 59724
rect 533522 59712 533528 59724
rect 533580 59712 533586 59764
rect 533798 59712 533804 59764
rect 533856 59752 533862 59764
rect 536282 59752 536288 59764
rect 533856 59724 536288 59752
rect 533856 59712 533862 59724
rect 536282 59712 536288 59724
rect 536340 59712 536346 59764
rect 123478 59576 123484 59628
rect 123536 59616 123542 59628
rect 125318 59616 125324 59628
rect 123536 59588 125324 59616
rect 123536 59576 123542 59588
rect 125318 59576 125324 59588
rect 125376 59576 125382 59628
rect 159358 59576 159364 59628
rect 159416 59616 159422 59628
rect 161290 59616 161296 59628
rect 159416 59588 161296 59616
rect 159416 59576 159422 59588
rect 161290 59576 161296 59588
rect 161348 59576 161354 59628
rect 198366 59576 198372 59628
rect 198424 59616 198430 59628
rect 200022 59616 200028 59628
rect 198424 59588 200028 59616
rect 198424 59576 198430 59588
rect 200022 59576 200028 59588
rect 200080 59576 200086 59628
rect 242802 59576 242808 59628
rect 242860 59616 242866 59628
rect 244090 59616 244096 59628
rect 242860 59588 244096 59616
rect 242860 59576 242866 59588
rect 244090 59576 244096 59588
rect 244148 59576 244154 59628
rect 269022 59576 269028 59628
rect 269080 59616 269086 59628
rect 270310 59616 270316 59628
rect 269080 59588 270316 59616
rect 269080 59576 269086 59588
rect 270310 59576 270316 59588
rect 270368 59576 270374 59628
rect 275922 59576 275928 59628
rect 275980 59616 275986 59628
rect 277118 59616 277124 59628
rect 275980 59588 277124 59616
rect 275980 59576 275986 59588
rect 277118 59576 277124 59588
rect 277176 59576 277182 59628
rect 284938 59576 284944 59628
rect 284996 59616 285002 59628
rect 286870 59616 286876 59628
rect 284996 59588 286876 59616
rect 284996 59576 285002 59588
rect 286870 59576 286876 59588
rect 286928 59576 286934 59628
rect 295242 59576 295248 59628
rect 295300 59616 295306 59628
rect 296622 59616 296628 59628
rect 295300 59588 296628 59616
rect 295300 59576 295306 59588
rect 296622 59576 296628 59588
rect 296680 59576 296686 59628
rect 324498 59576 324504 59628
rect 324556 59616 324562 59628
rect 325694 59616 325700 59628
rect 324556 59588 325700 59616
rect 324556 59576 324562 59588
rect 325694 59576 325700 59588
rect 325752 59576 325758 59628
rect 374086 59576 374092 59628
rect 374144 59616 374150 59628
rect 376018 59616 376024 59628
rect 374144 59588 376024 59616
rect 374144 59576 374150 59588
rect 376018 59576 376024 59588
rect 376076 59576 376082 59628
rect 419810 59576 419816 59628
rect 419868 59616 419874 59628
rect 421098 59616 421104 59628
rect 419868 59588 421104 59616
rect 419868 59576 419874 59588
rect 421098 59576 421104 59588
rect 421156 59576 421162 59628
rect 456886 59576 456892 59628
rect 456944 59616 456950 59628
rect 458266 59616 458272 59628
rect 456944 59588 458272 59616
rect 456944 59576 456950 59588
rect 458266 59576 458272 59588
rect 458324 59576 458330 59628
rect 492858 59576 492864 59628
rect 492916 59616 492922 59628
rect 494146 59616 494152 59628
rect 492916 59588 494152 59616
rect 492916 59576 492922 59588
rect 494146 59576 494152 59588
rect 494204 59576 494210 59628
rect 61930 59440 61936 59492
rect 61988 59480 61994 59492
rect 63954 59480 63960 59492
rect 61988 59452 63960 59480
rect 61988 59440 61994 59452
rect 63954 59440 63960 59452
rect 64012 59440 64018 59492
rect 113266 59440 113272 59492
rect 113324 59480 113330 59492
rect 114646 59480 114652 59492
rect 113324 59452 114652 59480
rect 113324 59440 113330 59452
rect 114646 59440 114652 59452
rect 114704 59440 114710 59492
rect 152458 59440 152464 59492
rect 152516 59480 152522 59492
rect 154482 59480 154488 59492
rect 152516 59452 154488 59480
rect 152516 59440 152522 59452
rect 154482 59440 154488 59452
rect 154540 59440 154546 59492
rect 165062 59440 165068 59492
rect 165120 59480 165126 59492
rect 167178 59480 167184 59492
rect 165120 59452 167184 59480
rect 165120 59440 165126 59452
rect 167178 59440 167184 59452
rect 167236 59440 167242 59492
rect 235902 59440 235908 59492
rect 235960 59480 235966 59492
rect 237374 59480 237380 59492
rect 235960 59452 237380 59480
rect 235960 59440 235966 59452
rect 237374 59440 237380 59452
rect 237432 59440 237438 59492
rect 244182 59440 244188 59492
rect 244240 59480 244246 59492
rect 246022 59480 246028 59492
rect 244240 59452 246028 59480
rect 244240 59440 244246 59452
rect 246022 59440 246028 59452
rect 246080 59440 246086 59492
rect 352742 59440 352748 59492
rect 352800 59480 352806 59492
rect 354674 59480 354680 59492
rect 352800 59452 354680 59480
rect 352800 59440 352806 59452
rect 354674 59440 354680 59452
rect 354732 59440 354738 59492
rect 497734 59440 497740 59492
rect 497792 59480 497798 59492
rect 499666 59480 499672 59492
rect 497792 59452 499672 59480
rect 497792 59440 497798 59452
rect 499666 59440 499672 59452
rect 499724 59440 499730 59492
rect 507486 59440 507492 59492
rect 507544 59480 507550 59492
rect 509418 59480 509424 59492
rect 507544 59452 509424 59480
rect 507544 59440 507550 59452
rect 509418 59440 509424 59452
rect 509476 59440 509482 59492
rect 11698 59372 11704 59424
rect 11756 59412 11762 59424
rect 59354 59412 59360 59424
rect 11756 59384 59360 59412
rect 11756 59372 11762 59384
rect 59354 59372 59360 59384
rect 59412 59372 59418 59424
rect 103514 59372 103520 59424
rect 103572 59412 103578 59424
rect 104894 59412 104900 59424
rect 103572 59384 104900 59412
rect 103572 59372 103578 59384
rect 104894 59372 104900 59384
rect 104952 59372 104958 59424
rect 542262 59372 542268 59424
rect 542320 59412 542326 59424
rect 582374 59412 582380 59424
rect 542320 59384 582380 59412
rect 542320 59372 542326 59384
rect 582374 59372 582380 59384
rect 582432 59372 582438 59424
rect 85022 59304 85028 59356
rect 85080 59344 85086 59356
rect 89714 59344 89720 59356
rect 85080 59316 89720 59344
rect 85080 59304 85086 59316
rect 89714 59304 89720 59316
rect 89772 59304 89778 59356
rect 168374 59304 168380 59356
rect 168432 59344 168438 59356
rect 173986 59344 173992 59356
rect 168432 59316 173992 59344
rect 168432 59304 168438 59316
rect 173986 59304 173992 59316
rect 174044 59304 174050 59356
rect 346394 59304 346400 59356
rect 346452 59344 346458 59356
rect 347774 59344 347780 59356
rect 346452 59316 347780 59344
rect 346452 59304 346458 59316
rect 347774 59304 347780 59316
rect 347832 59304 347838 59356
rect 447134 58896 447140 58948
rect 447192 58936 447198 58948
rect 448514 58936 448520 58948
rect 447192 58908 448520 58936
rect 447192 58896 447198 58908
rect 448514 58896 448520 58908
rect 448572 58896 448578 58948
rect 267734 58828 267740 58880
rect 267792 58868 267798 58880
rect 326154 58868 326160 58880
rect 267792 58840 326160 58868
rect 267792 58828 267798 58840
rect 326154 58828 326160 58840
rect 326212 58828 326218 58880
rect 371142 58828 371148 58880
rect 371200 58868 371206 58880
rect 427814 58868 427820 58880
rect 371200 58840 427820 58868
rect 371200 58828 371206 58840
rect 427814 58828 427820 58840
rect 427872 58828 427878 58880
rect 91002 58760 91008 58812
rect 91060 58800 91066 58812
rect 92290 58800 92296 58812
rect 91060 58772 92296 58800
rect 91060 58760 91066 58772
rect 92290 58760 92296 58772
rect 92348 58760 92354 58812
rect 190454 58760 190460 58812
rect 190512 58800 190518 58812
rect 304994 58800 305000 58812
rect 190512 58772 305000 58800
rect 190512 58760 190518 58772
rect 304994 58760 305000 58772
rect 305052 58760 305058 58812
rect 319622 58760 319628 58812
rect 319680 58800 319686 58812
rect 321738 58800 321744 58812
rect 319680 58772 321744 58800
rect 319680 58760 319686 58772
rect 321738 58760 321744 58772
rect 321796 58760 321802 58812
rect 335354 58760 335360 58812
rect 335412 58800 335418 58812
rect 345382 58800 345388 58812
rect 335412 58772 345388 58800
rect 335412 58760 335418 58772
rect 345382 58760 345388 58772
rect 345440 58760 345446 58812
rect 392578 58760 392584 58812
rect 392636 58800 392642 58812
rect 483474 58800 483480 58812
rect 392636 58772 483480 58800
rect 392636 58760 392642 58772
rect 483474 58760 483480 58772
rect 483532 58760 483538 58812
rect 237374 58692 237380 58744
rect 237432 58732 237438 58744
rect 441982 58732 441988 58744
rect 237432 58704 441988 58732
rect 237432 58692 237438 58704
rect 441982 58692 441988 58704
rect 442040 58692 442046 58744
rect 3418 58624 3424 58676
rect 3476 58664 3482 58676
rect 57974 58664 57980 58676
rect 3476 58636 57980 58664
rect 3476 58624 3482 58636
rect 57974 58624 57980 58636
rect 58032 58624 58038 58676
rect 104894 58624 104900 58676
rect 104952 58664 104958 58676
rect 118602 58664 118608 58676
rect 104952 58636 118608 58664
rect 104952 58624 104958 58636
rect 118602 58624 118608 58636
rect 118660 58624 118666 58676
rect 150434 58624 150440 58676
rect 150492 58664 150498 58676
rect 168282 58664 168288 58676
rect 150492 58636 168288 58664
rect 150492 58624 150498 58636
rect 168282 58624 168288 58636
rect 168340 58624 168346 58676
rect 193030 58624 193036 58676
rect 193088 58664 193094 58676
rect 231854 58664 231860 58676
rect 193088 58636 231860 58664
rect 193088 58624 193094 58636
rect 231854 58624 231860 58636
rect 231912 58624 231918 58676
rect 264790 58624 264796 58676
rect 264848 58664 264854 58676
rect 494054 58664 494060 58676
rect 264848 58636 494060 58664
rect 264848 58624 264854 58636
rect 494054 58624 494060 58636
rect 494112 58624 494118 58676
rect 91738 58488 91744 58540
rect 91796 58528 91802 58540
rect 94130 58528 94136 58540
rect 91796 58500 94136 58528
rect 91796 58488 91802 58500
rect 94130 58488 94136 58500
rect 94188 58488 94194 58540
rect 253566 58488 253572 58540
rect 253624 58528 253630 58540
rect 254302 58528 254308 58540
rect 253624 58500 254308 58528
rect 253624 58488 253630 58500
rect 254302 58488 254308 58500
rect 254360 58488 254366 58540
rect 320450 58488 320456 58540
rect 320508 58528 320514 58540
rect 321922 58528 321928 58540
rect 320508 58500 321928 58528
rect 320508 58488 320514 58500
rect 321922 58488 321928 58500
rect 321980 58488 321986 58540
rect 448146 58352 448152 58404
rect 448204 58392 448210 58404
rect 450170 58392 450176 58404
rect 448204 58364 450176 58392
rect 448204 58352 448210 58364
rect 450170 58352 450176 58364
rect 450228 58352 450234 58404
rect 446398 58080 446404 58132
rect 446456 58120 446462 58132
rect 447410 58120 447416 58132
rect 446456 58092 447416 58120
rect 446456 58080 446462 58092
rect 447410 58080 447416 58092
rect 447468 58080 447474 58132
rect 75914 57944 75920 57996
rect 75972 57984 75978 57996
rect 78490 57984 78496 57996
rect 75972 57956 78496 57984
rect 75972 57944 75978 57956
rect 78490 57944 78496 57956
rect 78548 57944 78554 57996
rect 354674 57944 354680 57996
rect 354732 57984 354738 57996
rect 360194 57984 360200 57996
rect 354732 57956 360200 57984
rect 354732 57944 354738 57956
rect 360194 57944 360200 57956
rect 360252 57944 360258 57996
rect 215294 57400 215300 57452
rect 215352 57440 215358 57452
rect 311986 57440 311992 57452
rect 215352 57412 311992 57440
rect 215352 57400 215358 57412
rect 311986 57400 311992 57412
rect 312044 57400 312050 57452
rect 161474 57332 161480 57384
rect 161532 57372 161538 57384
rect 295242 57372 295248 57384
rect 161532 57344 295248 57372
rect 161532 57332 161538 57344
rect 295242 57332 295248 57344
rect 295300 57332 295306 57384
rect 321554 57332 321560 57384
rect 321612 57372 321618 57384
rect 340874 57372 340880 57384
rect 321612 57344 340880 57372
rect 321612 57332 321618 57344
rect 340874 57332 340880 57344
rect 340932 57332 340938 57384
rect 383838 57332 383844 57384
rect 383896 57372 383902 57384
rect 470594 57372 470600 57384
rect 383896 57344 470600 57372
rect 383896 57332 383902 57344
rect 470594 57332 470600 57344
rect 470652 57332 470658 57384
rect 194594 57264 194600 57316
rect 194652 57304 194658 57316
rect 430574 57304 430580 57316
rect 194652 57276 430580 57304
rect 194652 57264 194658 57276
rect 430574 57264 430580 57276
rect 430632 57264 430638 57316
rect 53834 57196 53840 57248
rect 53892 57236 53898 57248
rect 71774 57236 71780 57248
rect 53892 57208 71780 57236
rect 53892 57196 53898 57208
rect 71774 57196 71780 57208
rect 71832 57196 71838 57248
rect 87966 57196 87972 57248
rect 88024 57236 88030 57248
rect 100754 57236 100760 57248
rect 88024 57208 100760 57236
rect 88024 57196 88030 57208
rect 100754 57196 100760 57208
rect 100812 57196 100818 57248
rect 267642 57196 267648 57248
rect 267700 57236 267706 57248
rect 507854 57236 507860 57248
rect 267700 57208 507860 57236
rect 267700 57196 267706 57208
rect 507854 57196 507860 57208
rect 507912 57196 507918 57248
rect 276014 56108 276020 56160
rect 276072 56148 276078 56160
rect 328546 56148 328552 56160
rect 276072 56120 328552 56148
rect 276072 56108 276078 56120
rect 328546 56108 328552 56120
rect 328604 56108 328610 56160
rect 206738 56040 206744 56092
rect 206796 56080 206802 56092
rect 281534 56080 281540 56092
rect 206796 56052 281540 56080
rect 206796 56040 206802 56052
rect 281534 56040 281540 56052
rect 281592 56040 281598 56092
rect 204254 55972 204260 56024
rect 204312 56012 204318 56024
rect 308950 56012 308956 56024
rect 204312 55984 308956 56012
rect 204312 55972 204318 55984
rect 308950 55972 308956 55984
rect 309008 55972 309014 56024
rect 316034 55972 316040 56024
rect 316092 56012 316098 56024
rect 463602 56012 463608 56024
rect 316092 55984 463608 56012
rect 316092 55972 316098 55984
rect 463602 55972 463608 55984
rect 463660 55972 463666 56024
rect 16574 55904 16580 55956
rect 16632 55944 16638 55956
rect 61930 55944 61936 55956
rect 16632 55916 61936 55944
rect 16632 55904 16638 55916
rect 61930 55904 61936 55916
rect 61988 55904 61994 55956
rect 186958 55904 186964 55956
rect 187016 55944 187022 55956
rect 427630 55944 427636 55956
rect 187016 55916 427636 55944
rect 187016 55904 187022 55916
rect 427630 55904 427636 55916
rect 427688 55904 427694 55956
rect 56594 55836 56600 55888
rect 56652 55876 56658 55888
rect 135162 55876 135168 55888
rect 56652 55848 135168 55876
rect 56652 55836 56658 55848
rect 135162 55836 135168 55848
rect 135220 55836 135226 55888
rect 277302 55836 277308 55888
rect 277360 55876 277366 55888
rect 547874 55876 547880 55888
rect 277360 55848 547880 55876
rect 277360 55836 277366 55848
rect 547874 55836 547880 55848
rect 547932 55836 547938 55888
rect 208394 54680 208400 54732
rect 208452 54720 208458 54732
rect 311894 54720 311900 54732
rect 208452 54692 311900 54720
rect 208452 54680 208458 54692
rect 311894 54680 311900 54692
rect 311952 54680 311958 54732
rect 418798 54680 418804 54732
rect 418856 54720 418862 54732
rect 488626 54720 488632 54732
rect 418856 54692 488632 54720
rect 418856 54680 418862 54692
rect 488626 54680 488632 54692
rect 488684 54680 488690 54732
rect 244182 54612 244188 54664
rect 244240 54652 244246 54664
rect 430574 54652 430580 54664
rect 244240 54624 430580 54652
rect 244240 54612 244246 54624
rect 430574 54612 430580 54624
rect 430632 54612 430638 54664
rect 26234 54544 26240 54596
rect 26292 54584 26298 54596
rect 64782 54584 64788 54596
rect 26292 54556 64788 54584
rect 26292 54544 26298 54556
rect 64782 54544 64788 54556
rect 64840 54544 64846 54596
rect 251174 54544 251180 54596
rect 251232 54584 251238 54596
rect 448514 54584 448520 54596
rect 251232 54556 448520 54584
rect 251232 54544 251238 54556
rect 448514 54544 448520 54556
rect 448572 54544 448578 54596
rect 60734 54476 60740 54528
rect 60792 54516 60798 54528
rect 135898 54516 135904 54528
rect 60792 54488 135904 54516
rect 60792 54476 60798 54488
rect 135898 54476 135904 54488
rect 135956 54476 135962 54528
rect 279878 54476 279884 54528
rect 279936 54516 279942 54528
rect 557534 54516 557540 54528
rect 279936 54488 557540 54516
rect 279936 54476 279942 54488
rect 557534 54476 557540 54488
rect 557592 54476 557598 54528
rect 193214 53252 193220 53304
rect 193272 53292 193278 53304
rect 307938 53292 307944 53304
rect 193272 53264 307944 53292
rect 193272 53252 193278 53264
rect 307938 53252 307944 53264
rect 307996 53252 308002 53304
rect 257982 53184 257988 53236
rect 258040 53224 258046 53236
rect 476114 53224 476120 53236
rect 258040 53196 476120 53224
rect 258040 53184 258046 53196
rect 476114 53184 476120 53196
rect 476172 53184 476178 53236
rect 142154 53116 142160 53168
rect 142212 53156 142218 53168
rect 418154 53156 418160 53168
rect 142212 53128 418160 53156
rect 142212 53116 142218 53128
rect 418154 53116 418160 53128
rect 418212 53116 418218 53168
rect 28994 53048 29000 53100
rect 29052 53088 29058 53100
rect 65978 53088 65984 53100
rect 29052 53060 65984 53088
rect 29052 53048 29058 53060
rect 65978 53048 65984 53060
rect 66036 53048 66042 53100
rect 280062 53048 280068 53100
rect 280120 53088 280126 53100
rect 561674 53088 561680 53100
rect 280120 53060 561680 53088
rect 280120 53048 280126 53060
rect 561674 53048 561680 53060
rect 561732 53048 561738 53100
rect 260834 51960 260840 52012
rect 260892 52000 260898 52012
rect 327074 52000 327080 52012
rect 260892 51972 327080 52000
rect 260892 51960 260898 51972
rect 327074 51960 327080 51972
rect 327132 51960 327138 52012
rect 204162 51892 204168 51944
rect 204220 51932 204226 51944
rect 284294 51932 284300 51944
rect 204220 51904 284300 51932
rect 204220 51892 204226 51904
rect 284294 51892 284300 51904
rect 284352 51892 284358 51944
rect 201494 51824 201500 51876
rect 201552 51864 201558 51876
rect 310514 51864 310520 51876
rect 201552 51836 310520 51864
rect 201552 51824 201558 51836
rect 310514 51824 310520 51836
rect 310572 51824 310578 51876
rect 311158 51824 311164 51876
rect 311216 51864 311222 51876
rect 463694 51864 463700 51876
rect 311216 51836 463700 51864
rect 311216 51824 311222 51836
rect 463694 51824 463700 51836
rect 463752 51824 463758 51876
rect 187694 51756 187700 51808
rect 187752 51796 187758 51808
rect 430666 51796 430672 51808
rect 187752 51768 430672 51796
rect 187752 51756 187758 51768
rect 430666 51756 430672 51768
rect 430724 51756 430730 51808
rect 4798 51688 4804 51740
rect 4856 51728 4862 51740
rect 92198 51728 92204 51740
rect 4856 51700 92204 51728
rect 4856 51688 4862 51700
rect 92198 51688 92204 51700
rect 92256 51688 92262 51740
rect 284110 51688 284116 51740
rect 284168 51728 284174 51740
rect 572714 51728 572720 51740
rect 284168 51700 572720 51728
rect 284168 51688 284174 51700
rect 572714 51688 572720 51700
rect 572772 51688 572778 51740
rect 218054 50532 218060 50584
rect 218112 50572 218118 50584
rect 314838 50572 314844 50584
rect 218112 50544 314844 50572
rect 218112 50532 218118 50544
rect 314838 50532 314844 50544
rect 314896 50532 314902 50584
rect 227530 50464 227536 50516
rect 227588 50504 227594 50516
rect 369854 50504 369860 50516
rect 227588 50476 369860 50504
rect 227588 50464 227594 50476
rect 369854 50464 369860 50476
rect 369912 50464 369918 50516
rect 383930 50464 383936 50516
rect 383988 50504 383994 50516
rect 466454 50504 466460 50516
rect 383988 50476 466460 50504
rect 383988 50464 383994 50476
rect 466454 50464 466460 50476
rect 466512 50464 466518 50516
rect 311894 50396 311900 50448
rect 311952 50436 311958 50448
rect 465074 50436 465080 50448
rect 311952 50408 465080 50436
rect 311952 50396 311958 50408
rect 465074 50396 465080 50408
rect 465132 50396 465138 50448
rect 14458 50328 14464 50380
rect 14516 50368 14522 50380
rect 91738 50368 91744 50380
rect 14516 50340 91744 50368
rect 14516 50328 14522 50340
rect 91738 50328 91744 50340
rect 91796 50328 91802 50380
rect 110414 50328 110420 50380
rect 110472 50368 110478 50380
rect 149698 50368 149704 50380
rect 110472 50340 149704 50368
rect 110472 50328 110478 50340
rect 149698 50328 149704 50340
rect 149756 50328 149762 50380
rect 283926 50328 283932 50380
rect 283984 50368 283990 50380
rect 575474 50368 575480 50380
rect 283984 50340 575480 50368
rect 283984 50328 283990 50340
rect 575474 50328 575480 50340
rect 575532 50328 575538 50380
rect 208210 49172 208216 49224
rect 208268 49212 208274 49224
rect 295334 49212 295340 49224
rect 208268 49184 295340 49212
rect 208268 49172 208274 49184
rect 295334 49172 295340 49184
rect 295392 49172 295398 49224
rect 371878 49172 371884 49224
rect 371936 49212 371942 49224
rect 480346 49212 480352 49224
rect 371936 49184 480352 49212
rect 371936 49172 371942 49184
rect 480346 49172 480352 49184
rect 480404 49172 480410 49224
rect 224770 49104 224776 49156
rect 224828 49144 224834 49156
rect 356054 49144 356060 49156
rect 224828 49116 356060 49144
rect 224828 49104 224834 49116
rect 356054 49104 356060 49116
rect 356112 49104 356118 49156
rect 402238 49104 402244 49156
rect 402296 49144 402302 49156
rect 534074 49144 534080 49156
rect 402296 49116 534080 49144
rect 402296 49104 402302 49116
rect 534074 49104 534080 49116
rect 534132 49104 534138 49156
rect 252462 49036 252468 49088
rect 252520 49076 252526 49088
rect 458174 49076 458180 49088
rect 252520 49048 458180 49076
rect 252520 49036 252526 49048
rect 458174 49036 458180 49048
rect 458232 49036 458238 49088
rect 52454 48968 52460 49020
rect 52512 49008 52518 49020
rect 102778 49008 102784 49020
rect 52512 48980 102784 49008
rect 52512 48968 52518 48980
rect 102778 48968 102784 48980
rect 102836 48968 102842 49020
rect 135254 48968 135260 49020
rect 135312 49008 135318 49020
rect 416866 49008 416872 49020
rect 135312 48980 416872 49008
rect 135312 48968 135318 48980
rect 416866 48968 416872 48980
rect 416924 48968 416930 49020
rect 208026 47744 208032 47796
rect 208084 47784 208090 47796
rect 299474 47784 299480 47796
rect 208084 47756 299480 47784
rect 208084 47744 208090 47756
rect 299474 47744 299480 47756
rect 299532 47744 299538 47796
rect 226242 47676 226248 47728
rect 226300 47716 226306 47728
rect 362954 47716 362960 47728
rect 226300 47688 362960 47716
rect 226300 47676 226306 47688
rect 362954 47676 362960 47688
rect 363012 47676 363018 47728
rect 405182 47676 405188 47728
rect 405240 47716 405246 47728
rect 540974 47716 540980 47728
rect 405240 47688 540980 47716
rect 405240 47676 405246 47688
rect 540974 47676 540980 47688
rect 541032 47676 541038 47728
rect 244274 47608 244280 47660
rect 244332 47648 244338 47660
rect 447134 47648 447140 47660
rect 244332 47620 447140 47648
rect 244332 47608 244338 47620
rect 447134 47608 447140 47620
rect 447192 47608 447198 47660
rect 17954 47540 17960 47592
rect 18012 47580 18018 47592
rect 95142 47580 95148 47592
rect 18012 47552 95148 47580
rect 18012 47540 18018 47552
rect 95142 47540 95148 47552
rect 95200 47540 95206 47592
rect 102134 47540 102140 47592
rect 102192 47580 102198 47592
rect 148502 47580 148508 47592
rect 102192 47552 148508 47580
rect 102192 47540 102198 47552
rect 148502 47540 148508 47552
rect 148560 47540 148566 47592
rect 253750 47540 253756 47592
rect 253808 47580 253814 47592
rect 465074 47580 465080 47592
rect 253808 47552 465080 47580
rect 253808 47540 253814 47552
rect 465074 47540 465080 47552
rect 465132 47540 465138 47592
rect 222102 46384 222108 46436
rect 222160 46424 222166 46436
rect 349246 46424 349252 46436
rect 222160 46396 349252 46424
rect 222160 46384 222166 46396
rect 349246 46384 349252 46396
rect 349304 46384 349310 46436
rect 370590 46384 370596 46436
rect 370648 46424 370654 46436
rect 480438 46424 480444 46436
rect 370648 46396 480444 46424
rect 370648 46384 370654 46396
rect 480438 46384 480444 46396
rect 480496 46384 480502 46436
rect 143534 46316 143540 46368
rect 143592 46356 143598 46368
rect 290642 46356 290648 46368
rect 143592 46328 290648 46356
rect 143592 46316 143598 46328
rect 290642 46316 290648 46328
rect 290700 46316 290706 46368
rect 401042 46316 401048 46368
rect 401100 46356 401106 46368
rect 525150 46356 525156 46368
rect 401100 46328 525156 46356
rect 401100 46316 401106 46328
rect 525150 46316 525156 46328
rect 525208 46316 525214 46368
rect 242802 46248 242808 46300
rect 242860 46288 242866 46300
rect 423674 46288 423680 46300
rect 242860 46260 423680 46288
rect 242860 46248 242866 46260
rect 423674 46248 423680 46260
rect 423732 46248 423738 46300
rect 44174 46180 44180 46232
rect 44232 46220 44238 46232
rect 101582 46220 101588 46232
rect 44232 46192 101588 46220
rect 44232 46180 44238 46192
rect 101582 46180 101588 46192
rect 101640 46180 101646 46232
rect 241514 46180 241520 46232
rect 241572 46220 241578 46232
rect 445754 46220 445760 46232
rect 241572 46192 445760 46220
rect 241572 46180 241578 46192
rect 445754 46180 445760 46192
rect 445812 46180 445818 46232
rect 220538 45024 220544 45076
rect 220596 45064 220602 45076
rect 345014 45064 345020 45076
rect 220596 45036 345020 45064
rect 220596 45024 220602 45036
rect 345014 45024 345020 45036
rect 345072 45024 345078 45076
rect 399478 45024 399484 45076
rect 399536 45064 399542 45076
rect 522298 45064 522304 45076
rect 399536 45036 522304 45064
rect 399536 45024 399542 45036
rect 522298 45024 522304 45036
rect 522356 45024 522362 45076
rect 147674 44956 147680 45008
rect 147732 44996 147738 45008
rect 290458 44996 290464 45008
rect 147732 44968 290464 44996
rect 147732 44956 147738 44968
rect 290458 44956 290464 44968
rect 290516 44956 290522 45008
rect 342898 44956 342904 45008
rect 342956 44996 342962 45008
rect 473446 44996 473452 45008
rect 342956 44968 473452 44996
rect 342956 44956 342962 44968
rect 473446 44956 473452 44968
rect 473504 44956 473510 45008
rect 240042 44888 240048 44940
rect 240100 44928 240106 44940
rect 412634 44928 412640 44940
rect 240100 44900 412640 44928
rect 240100 44888 240106 44900
rect 412634 44888 412640 44900
rect 412692 44888 412698 44940
rect 80054 44820 80060 44872
rect 80112 44860 80118 44872
rect 111242 44860 111248 44872
rect 80112 44832 111248 44860
rect 80112 44820 80118 44832
rect 111242 44820 111248 44832
rect 111300 44820 111306 44872
rect 198734 44820 198740 44872
rect 198792 44860 198798 44872
rect 433518 44860 433524 44872
rect 198792 44832 433524 44860
rect 198792 44820 198798 44832
rect 433518 44820 433524 44832
rect 433576 44820 433582 44872
rect 282914 43596 282920 43648
rect 282972 43636 282978 43648
rect 332594 43636 332600 43648
rect 282972 43608 332600 43636
rect 282972 43596 282978 43608
rect 332594 43596 332600 43608
rect 332652 43596 332658 43648
rect 380158 43596 380164 43648
rect 380216 43636 380222 43648
rect 452654 43636 452660 43648
rect 380216 43608 452660 43636
rect 380216 43596 380222 43608
rect 452654 43596 452660 43608
rect 452712 43596 452718 43648
rect 213730 43528 213736 43580
rect 213788 43568 213794 43580
rect 320174 43568 320180 43580
rect 213788 43540 320180 43568
rect 213788 43528 213794 43540
rect 320174 43528 320180 43540
rect 320232 43528 320238 43580
rect 391382 43528 391388 43580
rect 391440 43568 391446 43580
rect 491294 43568 491300 43580
rect 391440 43540 491300 43568
rect 391440 43528 391446 43540
rect 491294 43528 491300 43540
rect 491352 43528 491358 43580
rect 230290 43460 230296 43512
rect 230348 43500 230354 43512
rect 376754 43500 376760 43512
rect 230348 43472 376760 43500
rect 230348 43460 230354 43472
rect 376754 43460 376760 43472
rect 376812 43460 376818 43512
rect 382918 43460 382924 43512
rect 382976 43500 382982 43512
rect 483106 43500 483112 43512
rect 382976 43472 483112 43500
rect 382976 43460 382982 43472
rect 483106 43460 483112 43472
rect 483164 43460 483170 43512
rect 180794 43392 180800 43444
rect 180852 43432 180858 43444
rect 429194 43432 429200 43444
rect 180852 43404 429200 43432
rect 180852 43392 180858 43404
rect 429194 43392 429200 43404
rect 429252 43392 429258 43444
rect 220722 42236 220728 42288
rect 220780 42276 220786 42288
rect 340874 42276 340880 42288
rect 220780 42248 340880 42276
rect 220780 42236 220786 42248
rect 340874 42236 340880 42248
rect 340932 42236 340938 42288
rect 398282 42236 398288 42288
rect 398340 42276 398346 42288
rect 520274 42276 520280 42288
rect 398340 42248 520280 42276
rect 398340 42236 398346 42248
rect 520274 42236 520280 42248
rect 520332 42236 520338 42288
rect 340138 42168 340144 42220
rect 340196 42208 340202 42220
rect 471974 42208 471980 42220
rect 340196 42180 471980 42208
rect 340196 42168 340202 42180
rect 471974 42168 471980 42180
rect 472032 42168 472038 42220
rect 237190 42100 237196 42152
rect 237248 42140 237254 42152
rect 405734 42140 405740 42152
rect 237248 42112 405740 42140
rect 237248 42100 237254 42112
rect 405734 42100 405740 42112
rect 405792 42100 405798 42152
rect 173894 42032 173900 42084
rect 173952 42072 173958 42084
rect 426526 42072 426532 42084
rect 173952 42044 426532 42072
rect 173952 42032 173958 42044
rect 426526 42032 426532 42044
rect 426584 42032 426590 42084
rect 219342 40876 219348 40928
rect 219400 40916 219406 40928
rect 338114 40916 338120 40928
rect 219400 40888 338120 40916
rect 219400 40876 219406 40888
rect 338114 40876 338120 40888
rect 338172 40876 338178 40928
rect 398098 40876 398104 40928
rect 398156 40916 398162 40928
rect 516134 40916 516140 40928
rect 398156 40888 516140 40916
rect 398156 40876 398162 40888
rect 516134 40876 516140 40888
rect 516192 40876 516198 40928
rect 329834 40808 329840 40860
rect 329892 40848 329898 40860
rect 469306 40848 469312 40860
rect 329892 40820 469312 40848
rect 329892 40808 329898 40820
rect 469306 40808 469312 40820
rect 469364 40808 469370 40860
rect 237006 40740 237012 40792
rect 237064 40780 237070 40792
rect 401594 40780 401600 40792
rect 237064 40752 401600 40780
rect 237064 40740 237070 40752
rect 401594 40740 401600 40752
rect 401652 40740 401658 40792
rect 169754 40672 169760 40724
rect 169812 40712 169818 40724
rect 426710 40712 426716 40724
rect 169812 40684 426716 40712
rect 169812 40672 169818 40684
rect 426710 40672 426716 40684
rect 426768 40672 426774 40724
rect 217870 39516 217876 39568
rect 217928 39556 217934 39568
rect 333974 39556 333980 39568
rect 217928 39528 333980 39556
rect 217928 39516 217934 39528
rect 333974 39516 333980 39528
rect 334032 39516 334038 39568
rect 392670 39516 392676 39568
rect 392728 39556 392734 39568
rect 498194 39556 498200 39568
rect 392728 39528 498200 39556
rect 392728 39516 392734 39528
rect 498194 39516 498200 39528
rect 498252 39516 498258 39568
rect 329098 39448 329104 39500
rect 329156 39488 329162 39500
rect 469490 39488 469496 39500
rect 329156 39460 469496 39488
rect 329156 39448 329162 39460
rect 469490 39448 469496 39460
rect 469548 39448 469554 39500
rect 235902 39380 235908 39432
rect 235960 39420 235966 39432
rect 398834 39420 398840 39432
rect 235960 39392 398840 39420
rect 235960 39380 235966 39392
rect 398834 39380 398840 39392
rect 398892 39380 398898 39432
rect 166994 39312 167000 39364
rect 167052 39352 167058 39364
rect 425054 39352 425060 39364
rect 167052 39324 425060 39352
rect 167052 39312 167058 39324
rect 425054 39312 425060 39324
rect 425112 39312 425118 39364
rect 314654 38088 314660 38140
rect 314712 38128 314718 38140
rect 341150 38128 341156 38140
rect 314712 38100 341156 38128
rect 314712 38088 314718 38100
rect 341150 38088 341156 38100
rect 341208 38088 341214 38140
rect 387058 38088 387064 38140
rect 387116 38128 387122 38140
rect 477494 38128 477500 38140
rect 387116 38100 477500 38128
rect 387116 38088 387122 38100
rect 477494 38088 477500 38100
rect 477552 38088 477558 38140
rect 217686 38020 217692 38072
rect 217744 38060 217750 38072
rect 331214 38060 331220 38072
rect 217744 38032 331220 38060
rect 217744 38020 217750 38032
rect 331214 38020 331220 38032
rect 331272 38020 331278 38072
rect 391198 38020 391204 38072
rect 391256 38060 391262 38072
rect 495434 38060 495440 38072
rect 391256 38032 495440 38060
rect 391256 38020 391262 38032
rect 495434 38020 495440 38032
rect 495492 38020 495498 38072
rect 234430 37952 234436 38004
rect 234488 37992 234494 38004
rect 394694 37992 394700 38004
rect 234488 37964 394700 37992
rect 234488 37952 234494 37964
rect 394694 37952 394700 37964
rect 394752 37952 394758 38004
rect 178678 37884 178684 37936
rect 178736 37924 178742 37936
rect 427906 37924 427912 37936
rect 178736 37896 427912 37924
rect 178736 37884 178742 37896
rect 427906 37884 427912 37896
rect 427964 37884 427970 37936
rect 216582 36660 216588 36712
rect 216640 36700 216646 36712
rect 327074 36700 327080 36712
rect 216640 36672 327080 36700
rect 216640 36660 216646 36672
rect 327074 36660 327080 36672
rect 327132 36660 327138 36712
rect 354030 36660 354036 36712
rect 354088 36700 354094 36712
rect 476390 36700 476396 36712
rect 354088 36672 476396 36700
rect 354088 36660 354094 36672
rect 476390 36660 476396 36672
rect 476448 36660 476454 36712
rect 233142 36592 233148 36644
rect 233200 36632 233206 36644
rect 387794 36632 387800 36644
rect 233200 36604 387800 36632
rect 233200 36592 233206 36604
rect 387794 36592 387800 36604
rect 387852 36592 387858 36644
rect 404998 36592 405004 36644
rect 405056 36632 405062 36644
rect 545114 36632 545120 36644
rect 405056 36604 545120 36632
rect 405056 36592 405062 36604
rect 545114 36592 545120 36604
rect 545172 36592 545178 36644
rect 88334 36524 88340 36576
rect 88392 36564 88398 36576
rect 144362 36564 144368 36576
rect 88392 36536 144368 36564
rect 88392 36524 88398 36536
rect 144362 36524 144368 36536
rect 144420 36524 144426 36576
rect 256602 36524 256608 36576
rect 256660 36564 256666 36576
rect 473354 36564 473360 36576
rect 256660 36536 473360 36564
rect 256660 36524 256666 36536
rect 473354 36524 473360 36536
rect 473412 36524 473418 36576
rect 215202 35300 215208 35352
rect 215260 35340 215266 35352
rect 324314 35340 324320 35352
rect 215260 35312 324320 35340
rect 215260 35300 215266 35312
rect 324314 35300 324320 35312
rect 324372 35300 324378 35352
rect 345658 35300 345664 35352
rect 345716 35340 345722 35352
rect 473630 35340 473636 35352
rect 345716 35312 473636 35340
rect 345716 35300 345722 35312
rect 473630 35300 473636 35312
rect 473688 35300 473694 35352
rect 230106 35232 230112 35284
rect 230164 35272 230170 35284
rect 380894 35272 380900 35284
rect 230164 35244 380900 35272
rect 230164 35232 230170 35244
rect 380894 35232 380900 35244
rect 380952 35232 380958 35284
rect 403618 35232 403624 35284
rect 403676 35272 403682 35284
rect 538214 35272 538220 35284
rect 403676 35244 538220 35272
rect 403676 35232 403682 35244
rect 538214 35232 538220 35244
rect 538272 35232 538278 35284
rect 85574 35164 85580 35216
rect 85632 35204 85638 35216
rect 142798 35204 142804 35216
rect 85632 35176 142804 35204
rect 85632 35164 85638 35176
rect 142798 35164 142804 35176
rect 142856 35164 142862 35216
rect 255222 35164 255228 35216
rect 255280 35204 255286 35216
rect 469214 35204 469220 35216
rect 255280 35176 469220 35204
rect 255280 35164 255286 35176
rect 469214 35164 469220 35176
rect 469272 35164 469278 35216
rect 197354 33940 197360 33992
rect 197412 33980 197418 33992
rect 309134 33980 309140 33992
rect 197412 33952 309140 33980
rect 197412 33940 197418 33952
rect 309134 33940 309140 33952
rect 309192 33940 309198 33992
rect 383010 33940 383016 33992
rect 383068 33980 383074 33992
rect 463694 33980 463700 33992
rect 383068 33952 463700 33980
rect 383068 33940 383074 33952
rect 463694 33940 463700 33952
rect 463752 33940 463758 33992
rect 223482 33872 223488 33924
rect 223540 33912 223546 33924
rect 351914 33912 351920 33924
rect 223540 33884 351920 33912
rect 223540 33872 223546 33884
rect 351914 33872 351920 33884
rect 351972 33872 351978 33924
rect 403618 33872 403624 33924
rect 403676 33912 403682 33924
rect 490006 33912 490012 33924
rect 403676 33884 490012 33912
rect 403676 33872 403682 33884
rect 490006 33872 490012 33884
rect 490064 33872 490070 33924
rect 131114 33804 131120 33856
rect 131172 33844 131178 33856
rect 415394 33844 415400 33856
rect 131172 33816 415400 33844
rect 131172 33804 131178 33816
rect 415394 33804 415400 33816
rect 415452 33804 415458 33856
rect 282822 33736 282828 33788
rect 282880 33776 282886 33788
rect 568574 33776 568580 33788
rect 282880 33748 568580 33776
rect 282880 33736 282886 33748
rect 568574 33736 568580 33748
rect 568632 33736 568638 33788
rect 176654 32580 176660 32632
rect 176712 32620 176718 32632
rect 303614 32620 303620 32632
rect 176712 32592 303620 32620
rect 176712 32580 176718 32592
rect 303614 32580 303620 32592
rect 303672 32580 303678 32632
rect 372154 32580 372160 32632
rect 372212 32620 372218 32632
rect 423766 32620 423772 32632
rect 372212 32592 423772 32620
rect 372212 32580 372218 32592
rect 423766 32580 423772 32592
rect 423824 32580 423830 32632
rect 224586 32512 224592 32564
rect 224644 32552 224650 32564
rect 358814 32552 358820 32564
rect 224644 32524 358820 32552
rect 224644 32512 224650 32524
rect 358814 32512 358820 32524
rect 358872 32512 358878 32564
rect 378870 32512 378876 32564
rect 378928 32552 378934 32564
rect 483290 32552 483296 32564
rect 378928 32524 483296 32552
rect 378928 32512 378934 32524
rect 483290 32512 483296 32524
rect 483348 32512 483354 32564
rect 201586 32444 201592 32496
rect 201644 32484 201650 32496
rect 434714 32484 434720 32496
rect 201644 32456 434720 32484
rect 201644 32444 201650 32456
rect 434714 32444 434720 32456
rect 434772 32444 434778 32496
rect 77294 32376 77300 32428
rect 77352 32416 77358 32428
rect 141602 32416 141608 32428
rect 77352 32388 141608 32416
rect 77352 32376 77358 32388
rect 141602 32376 141608 32388
rect 141660 32376 141666 32428
rect 281442 32376 281448 32428
rect 281500 32416 281506 32428
rect 564526 32416 564532 32428
rect 281500 32388 564532 32416
rect 281500 32376 281506 32388
rect 564526 32376 564532 32388
rect 564584 32376 564590 32428
rect 278774 31220 278780 31272
rect 278832 31260 278838 31272
rect 331398 31260 331404 31272
rect 278832 31232 331404 31260
rect 278832 31220 278838 31232
rect 331398 31220 331404 31232
rect 331456 31220 331462 31272
rect 140774 31152 140780 31204
rect 140832 31192 140838 31204
rect 289078 31192 289084 31204
rect 140832 31164 289084 31192
rect 140832 31152 140838 31164
rect 289078 31152 289084 31164
rect 289136 31152 289142 31204
rect 356790 31152 356796 31204
rect 356848 31192 356854 31204
rect 476206 31192 476212 31204
rect 356848 31164 476212 31192
rect 356848 31152 356854 31164
rect 476206 31152 476212 31164
rect 476264 31152 476270 31204
rect 253566 31084 253572 31136
rect 253624 31124 253630 31136
rect 462314 31124 462320 31136
rect 253624 31096 462320 31124
rect 253624 31084 253630 31096
rect 462314 31084 462320 31096
rect 462372 31084 462378 31136
rect 70394 31016 70400 31068
rect 70452 31056 70458 31068
rect 138658 31056 138664 31068
rect 70452 31028 138664 31056
rect 70452 31016 70458 31028
rect 138658 31016 138664 31028
rect 138716 31016 138722 31068
rect 202782 31016 202788 31068
rect 202840 31056 202846 31068
rect 277394 31056 277400 31068
rect 202840 31028 277400 31056
rect 202840 31016 202846 31028
rect 277394 31016 277400 31028
rect 277452 31016 277458 31068
rect 278682 31016 278688 31068
rect 278740 31056 278746 31068
rect 554774 31056 554780 31068
rect 278740 31028 554780 31056
rect 278740 31016 278746 31028
rect 554774 31016 554780 31028
rect 554832 31016 554838 31068
rect 271874 29792 271880 29844
rect 271932 29832 271938 29844
rect 329926 29832 329932 29844
rect 271932 29804 329932 29832
rect 271932 29792 271938 29804
rect 329926 29792 329932 29804
rect 329984 29792 329990 29844
rect 400950 29792 400956 29844
rect 401008 29832 401014 29844
rect 488534 29832 488540 29844
rect 401008 29804 488540 29832
rect 401008 29792 401014 29804
rect 488534 29792 488540 29804
rect 488592 29792 488598 29844
rect 250990 29724 250996 29776
rect 251048 29764 251054 29776
rect 455414 29764 455420 29776
rect 251048 29736 455420 29764
rect 251048 29724 251054 29736
rect 455414 29724 455420 29736
rect 455472 29724 455478 29776
rect 201310 29656 201316 29708
rect 201368 29696 201374 29708
rect 274634 29696 274640 29708
rect 201368 29668 274640 29696
rect 201368 29656 201374 29668
rect 274634 29656 274640 29668
rect 274692 29656 274698 29708
rect 277026 29656 277032 29708
rect 277084 29696 277090 29708
rect 550634 29696 550640 29708
rect 277084 29668 550640 29696
rect 277084 29656 277090 29668
rect 550634 29656 550640 29668
rect 550692 29656 550698 29708
rect 67634 29588 67640 29640
rect 67692 29628 67698 29640
rect 137462 29628 137468 29640
rect 67692 29600 137468 29628
rect 67692 29588 67698 29600
rect 137462 29588 137468 29600
rect 137520 29588 137526 29640
rect 144914 29588 144920 29640
rect 144972 29628 144978 29640
rect 419534 29628 419540 29640
rect 144972 29600 419540 29628
rect 144972 29588 144978 29600
rect 419534 29588 419540 29600
rect 419592 29588 419598 29640
rect 227346 28432 227352 28484
rect 227404 28472 227410 28484
rect 365714 28472 365720 28484
rect 227404 28444 365720 28472
rect 227404 28432 227410 28444
rect 365714 28432 365720 28444
rect 365772 28432 365778 28484
rect 371970 28432 371976 28484
rect 372028 28472 372034 28484
rect 420914 28472 420920 28484
rect 372028 28444 420920 28472
rect 372028 28432 372034 28444
rect 420914 28432 420920 28444
rect 420972 28432 420978 28484
rect 126974 28364 126980 28416
rect 127032 28404 127038 28416
rect 284938 28404 284944 28416
rect 127032 28376 284944 28404
rect 127032 28364 127038 28376
rect 284938 28364 284944 28376
rect 284996 28364 285002 28416
rect 376110 28364 376116 28416
rect 376168 28404 376174 28416
rect 481634 28404 481640 28416
rect 376168 28376 481640 28404
rect 376168 28364 376174 28376
rect 481634 28364 481640 28376
rect 481692 28364 481698 28416
rect 191834 28296 191840 28348
rect 191892 28336 191898 28348
rect 431954 28336 431960 28348
rect 191892 28308 431960 28336
rect 191892 28296 191898 28308
rect 431954 28296 431960 28308
rect 432012 28296 432018 28348
rect 37274 28228 37280 28280
rect 37332 28268 37338 28280
rect 98822 28268 98828 28280
rect 37332 28240 98828 28268
rect 37332 28228 37338 28240
rect 98822 28228 98828 28240
rect 98880 28228 98886 28280
rect 273162 28228 273168 28280
rect 273220 28268 273226 28280
rect 532694 28268 532700 28280
rect 273220 28240 532700 28268
rect 273220 28228 273226 28240
rect 532694 28228 532700 28240
rect 532752 28228 532758 28280
rect 264974 27004 264980 27056
rect 265032 27044 265038 27056
rect 327258 27044 327264 27056
rect 265032 27016 327264 27044
rect 265032 27004 265038 27016
rect 327258 27004 327264 27016
rect 327316 27004 327322 27056
rect 332594 27004 332600 27056
rect 332652 27044 332658 27056
rect 470686 27044 470692 27056
rect 332652 27016 470692 27044
rect 332652 27004 332658 27016
rect 470686 27004 470692 27016
rect 470744 27004 470750 27056
rect 248322 26936 248328 26988
rect 248380 26976 248386 26988
rect 444374 26976 444380 26988
rect 248380 26948 444380 26976
rect 248380 26936 248386 26948
rect 444374 26936 444380 26948
rect 444432 26936 444438 26988
rect 22094 26868 22100 26920
rect 22152 26908 22158 26920
rect 94498 26908 94504 26920
rect 22152 26880 94504 26908
rect 22152 26868 22158 26880
rect 94498 26868 94504 26880
rect 94556 26868 94562 26920
rect 200022 26868 200028 26920
rect 200080 26908 200086 26920
rect 267826 26908 267832 26920
rect 200080 26880 267832 26908
rect 200080 26868 200086 26880
rect 267826 26868 267832 26880
rect 267884 26868 267890 26920
rect 270310 26868 270316 26920
rect 270368 26908 270374 26920
rect 523218 26908 523224 26920
rect 270368 26880 523224 26908
rect 270368 26868 270374 26880
rect 523218 26868 523224 26880
rect 523276 26868 523282 26920
rect 136634 25712 136640 25764
rect 136692 25752 136698 25764
rect 287698 25752 287704 25764
rect 136692 25724 287704 25752
rect 136692 25712 136698 25724
rect 287698 25712 287704 25724
rect 287756 25712 287762 25764
rect 246850 25644 246856 25696
rect 246908 25684 246914 25696
rect 437474 25684 437480 25696
rect 246908 25656 437480 25684
rect 246908 25644 246914 25656
rect 437474 25644 437480 25656
rect 437532 25644 437538 25696
rect 248414 25576 248420 25628
rect 248472 25616 248478 25628
rect 447410 25616 447416 25628
rect 248472 25588 447416 25616
rect 248472 25576 248478 25588
rect 447410 25576 447416 25588
rect 447468 25576 447474 25628
rect 91094 25508 91100 25560
rect 91152 25548 91158 25560
rect 113818 25548 113824 25560
rect 91152 25520 113824 25548
rect 91152 25508 91158 25520
rect 113818 25508 113824 25520
rect 113876 25508 113882 25560
rect 198550 25508 198556 25560
rect 198608 25548 198614 25560
rect 259454 25548 259460 25560
rect 198608 25520 259460 25548
rect 198608 25508 198614 25520
rect 259454 25508 259460 25520
rect 259512 25508 259518 25560
rect 264882 25508 264888 25560
rect 264940 25548 264946 25560
rect 505094 25548 505100 25560
rect 264940 25520 505100 25548
rect 264940 25508 264946 25520
rect 505094 25508 505100 25520
rect 505152 25508 505158 25560
rect 247034 24284 247040 24336
rect 247092 24324 247098 24336
rect 322934 24324 322940 24336
rect 247092 24296 322940 24324
rect 247092 24284 247098 24296
rect 322934 24284 322940 24296
rect 322992 24284 322998 24336
rect 320818 24216 320824 24268
rect 320876 24256 320882 24268
rect 466638 24256 466644 24268
rect 320876 24228 466644 24256
rect 320876 24216 320882 24228
rect 466638 24216 466644 24228
rect 466696 24216 466702 24268
rect 245562 24148 245568 24200
rect 245620 24188 245626 24200
rect 433334 24188 433340 24200
rect 245620 24160 433340 24188
rect 245620 24148 245626 24160
rect 433334 24148 433340 24160
rect 433392 24148 433398 24200
rect 86954 24080 86960 24132
rect 87012 24120 87018 24132
rect 112438 24120 112444 24132
rect 87012 24092 112444 24120
rect 87012 24080 87018 24092
rect 112438 24080 112444 24092
rect 112496 24080 112502 24132
rect 194410 24080 194416 24132
rect 194468 24120 194474 24132
rect 249794 24120 249800 24132
rect 194468 24092 249800 24120
rect 194468 24080 194474 24092
rect 249794 24080 249800 24092
rect 249852 24080 249858 24132
rect 263318 24080 263324 24132
rect 263376 24120 263382 24132
rect 500954 24120 500960 24132
rect 263376 24092 500960 24120
rect 263376 24080 263382 24092
rect 500954 24080 500960 24092
rect 501012 24080 501018 24132
rect 235994 22924 236000 22976
rect 236052 22964 236058 22976
rect 320266 22964 320272 22976
rect 236052 22936 320272 22964
rect 236052 22924 236058 22936
rect 320266 22924 320272 22936
rect 320324 22924 320330 22976
rect 307018 22856 307024 22908
rect 307076 22896 307082 22908
rect 463878 22896 463884 22908
rect 307076 22868 463884 22896
rect 307076 22856 307082 22868
rect 463878 22856 463884 22868
rect 463936 22856 463942 22908
rect 81434 22788 81440 22840
rect 81492 22828 81498 22840
rect 141418 22828 141424 22840
rect 81492 22800 141424 22828
rect 81492 22788 81498 22800
rect 141418 22788 141424 22800
rect 141476 22788 141482 22840
rect 243906 22788 243912 22840
rect 243964 22828 243970 22840
rect 426434 22828 426440 22840
rect 243964 22800 426440 22828
rect 243964 22788 243970 22800
rect 426434 22788 426440 22800
rect 426492 22788 426498 22840
rect 15838 22720 15844 22772
rect 15896 22760 15902 22772
rect 93118 22760 93124 22772
rect 15896 22732 93124 22760
rect 15896 22720 15902 22732
rect 93118 22720 93124 22732
rect 93176 22720 93182 22772
rect 194226 22720 194232 22772
rect 194284 22760 194290 22772
rect 245654 22760 245660 22772
rect 194284 22732 245660 22760
rect 194284 22720 194290 22732
rect 245654 22720 245660 22732
rect 245712 22720 245718 22772
rect 263502 22720 263508 22772
rect 263560 22760 263566 22772
rect 498286 22760 498292 22772
rect 263560 22732 498292 22760
rect 263560 22720 263566 22732
rect 498286 22720 498292 22732
rect 498344 22720 498350 22772
rect 226334 21564 226340 21616
rect 226392 21604 226398 21616
rect 317598 21604 317604 21616
rect 226392 21576 317604 21604
rect 226392 21564 226398 21576
rect 317598 21564 317604 21576
rect 317656 21564 317662 21616
rect 385770 21564 385776 21616
rect 385828 21604 385834 21616
rect 484394 21604 484400 21616
rect 385828 21576 484400 21604
rect 385828 21564 385834 21576
rect 484394 21564 484400 21576
rect 484452 21564 484458 21616
rect 287054 21496 287060 21548
rect 287112 21536 287118 21548
rect 458266 21536 458272 21548
rect 287112 21508 458272 21536
rect 287112 21496 287118 21508
rect 458266 21496 458272 21508
rect 458324 21496 458330 21548
rect 241238 21428 241244 21480
rect 241296 21468 241302 21480
rect 419534 21468 419540 21480
rect 241296 21440 419540 21468
rect 241296 21428 241302 21440
rect 419534 21428 419540 21440
rect 419592 21428 419598 21480
rect 77386 21360 77392 21412
rect 77444 21400 77450 21412
rect 109678 21400 109684 21412
rect 77444 21372 109684 21400
rect 77444 21360 77450 21372
rect 109678 21360 109684 21372
rect 109736 21360 109742 21412
rect 188982 21360 188988 21412
rect 189040 21400 189046 21412
rect 227714 21400 227720 21412
rect 189040 21372 227720 21400
rect 189040 21360 189046 21372
rect 227714 21360 227720 21372
rect 227772 21360 227778 21412
rect 260558 21360 260564 21412
rect 260616 21400 260622 21412
rect 489914 21400 489920 21412
rect 260616 21372 489920 21400
rect 260616 21360 260622 21372
rect 489914 21360 489920 21372
rect 489972 21360 489978 21412
rect 404354 20136 404360 20188
rect 404412 20176 404418 20188
rect 490190 20176 490196 20188
rect 404412 20148 490196 20176
rect 404412 20136 404418 20148
rect 490190 20136 490196 20148
rect 490248 20136 490254 20188
rect 222194 20068 222200 20120
rect 222252 20108 222258 20120
rect 316126 20108 316132 20120
rect 222252 20080 316132 20108
rect 222252 20068 222258 20080
rect 316126 20068 316132 20080
rect 316184 20068 316190 20120
rect 385678 20068 385684 20120
rect 385736 20108 385742 20120
rect 473446 20108 473452 20120
rect 385736 20080 473452 20108
rect 385736 20068 385742 20080
rect 473446 20068 473452 20080
rect 473504 20068 473510 20120
rect 241422 20000 241428 20052
rect 241480 20040 241486 20052
rect 415394 20040 415400 20052
rect 241480 20012 415400 20040
rect 241480 20000 241486 20012
rect 415394 20000 415400 20012
rect 415452 20000 415458 20052
rect 55214 19932 55220 19984
rect 55272 19972 55278 19984
rect 104342 19972 104348 19984
rect 55272 19944 104348 19972
rect 55272 19932 55278 19944
rect 104342 19932 104348 19944
rect 104400 19932 104406 19984
rect 113174 19932 113180 19984
rect 113232 19972 113238 19984
rect 151262 19972 151268 19984
rect 113232 19944 151268 19972
rect 113232 19932 113238 19944
rect 151262 19932 151268 19944
rect 151320 19932 151326 19984
rect 187510 19932 187516 19984
rect 187568 19972 187574 19984
rect 224954 19972 224960 19984
rect 187568 19944 224960 19972
rect 187568 19932 187574 19944
rect 224954 19932 224960 19944
rect 225012 19932 225018 19984
rect 260742 19932 260748 19984
rect 260800 19972 260806 19984
rect 487154 19972 487160 19984
rect 260800 19944 487160 19972
rect 260800 19932 260806 19944
rect 487154 19932 487160 19944
rect 487212 19932 487218 19984
rect 363690 18776 363696 18828
rect 363748 18816 363754 18828
rect 478874 18816 478880 18828
rect 363748 18788 478880 18816
rect 363748 18776 363754 18788
rect 478874 18776 478880 18788
rect 478932 18776 478938 18828
rect 229094 18708 229100 18760
rect 229152 18748 229158 18760
rect 317414 18748 317420 18760
rect 229152 18720 317420 18748
rect 229152 18708 229158 18720
rect 317414 18708 317420 18720
rect 317472 18708 317478 18760
rect 400858 18708 400864 18760
rect 400916 18748 400922 18760
rect 531406 18748 531412 18760
rect 400916 18720 531412 18748
rect 400916 18708 400922 18720
rect 531406 18708 531412 18720
rect 531464 18708 531470 18760
rect 238662 18640 238668 18692
rect 238720 18680 238726 18692
rect 408494 18680 408500 18692
rect 238720 18652 408500 18680
rect 238720 18640 238726 18652
rect 408494 18640 408500 18652
rect 408552 18640 408558 18692
rect 48314 18572 48320 18624
rect 48372 18612 48378 18624
rect 101398 18612 101404 18624
rect 48372 18584 101404 18612
rect 48372 18572 48378 18584
rect 101398 18572 101404 18584
rect 101456 18572 101462 18624
rect 106274 18572 106280 18624
rect 106332 18612 106338 18624
rect 148318 18612 148324 18624
rect 106332 18584 148324 18612
rect 106332 18572 106338 18584
rect 148318 18572 148324 18584
rect 148376 18572 148382 18624
rect 186222 18572 186228 18624
rect 186280 18612 186286 18624
rect 218146 18612 218152 18624
rect 186280 18584 218152 18612
rect 186280 18572 186286 18584
rect 218146 18572 218152 18584
rect 218204 18572 218210 18624
rect 259362 18572 259368 18624
rect 259420 18612 259426 18624
rect 483014 18612 483020 18624
rect 259420 18584 483020 18612
rect 259420 18572 259426 18584
rect 483014 18572 483020 18584
rect 483072 18572 483078 18624
rect 211154 17348 211160 17400
rect 211212 17388 211218 17400
rect 313274 17388 313280 17400
rect 211212 17360 313280 17388
rect 211212 17348 211218 17360
rect 313274 17348 313280 17360
rect 313332 17348 313338 17400
rect 347774 17348 347780 17400
rect 347832 17388 347838 17400
rect 474734 17388 474740 17400
rect 347832 17360 474740 17388
rect 347832 17348 347838 17360
rect 474734 17348 474740 17360
rect 474792 17348 474798 17400
rect 91002 17280 91008 17332
rect 91060 17320 91066 17332
rect 121454 17320 121460 17332
rect 91060 17292 121460 17320
rect 91060 17280 91066 17292
rect 121454 17280 121460 17292
rect 121512 17280 121518 17332
rect 234246 17280 234252 17332
rect 234304 17320 234310 17332
rect 390554 17320 390560 17332
rect 234304 17292 390560 17320
rect 234304 17280 234310 17292
rect 390554 17280 390560 17292
rect 390612 17280 390618 17332
rect 395338 17280 395344 17332
rect 395396 17320 395402 17332
rect 509234 17320 509240 17332
rect 395396 17292 509240 17320
rect 395396 17280 395402 17292
rect 509234 17280 509240 17292
rect 509292 17280 509298 17332
rect 30374 17212 30380 17264
rect 30432 17252 30438 17264
rect 97258 17252 97264 17264
rect 30432 17224 97264 17252
rect 30432 17212 30438 17224
rect 97258 17212 97264 17224
rect 97316 17212 97322 17264
rect 184750 17212 184756 17264
rect 184808 17252 184814 17264
rect 213914 17252 213920 17264
rect 184808 17224 213920 17252
rect 184808 17212 184814 17224
rect 213914 17212 213920 17224
rect 213972 17212 213978 17264
rect 257706 17212 257712 17264
rect 257764 17252 257770 17264
rect 480254 17252 480260 17264
rect 257764 17224 480260 17252
rect 257764 17212 257770 17224
rect 480254 17212 480260 17224
rect 480312 17212 480318 17264
rect 284386 16464 284392 16516
rect 284444 16504 284450 16516
rect 456886 16504 456892 16516
rect 284444 16476 456892 16504
rect 284444 16464 284450 16476
rect 456886 16464 456892 16476
rect 456944 16464 456950 16516
rect 280706 16396 280712 16448
rect 280764 16436 280770 16448
rect 457070 16436 457076 16448
rect 280764 16408 457076 16436
rect 280764 16396 280770 16408
rect 457070 16396 457076 16408
rect 457128 16396 457134 16448
rect 276658 16328 276664 16380
rect 276716 16368 276722 16380
rect 455506 16368 455512 16380
rect 276716 16340 455512 16368
rect 276716 16328 276722 16340
rect 455506 16328 455512 16340
rect 455564 16328 455570 16380
rect 273254 16260 273260 16312
rect 273312 16300 273318 16312
rect 454034 16300 454040 16312
rect 273312 16272 454040 16300
rect 273312 16260 273318 16272
rect 454034 16260 454040 16272
rect 454092 16260 454098 16312
rect 270034 16192 270040 16244
rect 270092 16232 270098 16244
rect 453022 16232 453028 16244
rect 270092 16204 453028 16232
rect 270092 16192 270098 16204
rect 453022 16192 453028 16204
rect 453080 16192 453086 16244
rect 266538 16124 266544 16176
rect 266596 16164 266602 16176
rect 452838 16164 452844 16176
rect 266596 16136 452844 16164
rect 266596 16124 266602 16136
rect 452838 16124 452844 16136
rect 452896 16124 452902 16176
rect 262490 16056 262496 16108
rect 262548 16096 262554 16108
rect 451274 16096 451280 16108
rect 262548 16068 451280 16096
rect 262548 16056 262554 16068
rect 451274 16056 451280 16068
rect 451332 16056 451338 16108
rect 259546 15988 259552 16040
rect 259604 16028 259610 16040
rect 449986 16028 449992 16040
rect 259604 16000 449992 16028
rect 259604 15988 259610 16000
rect 449986 15988 449992 16000
rect 450044 15988 450050 16040
rect 255866 15920 255872 15972
rect 255924 15960 255930 15972
rect 450170 15960 450176 15972
rect 255924 15932 450176 15960
rect 255924 15920 255930 15932
rect 450170 15920 450176 15932
rect 450228 15920 450234 15972
rect 85298 15852 85304 15904
rect 85356 15892 85362 15904
rect 104066 15892 104072 15904
rect 85356 15864 104072 15892
rect 85356 15852 85362 15864
rect 104066 15852 104072 15864
rect 104124 15852 104130 15904
rect 109034 15852 109040 15904
rect 109092 15892 109098 15904
rect 117958 15892 117964 15904
rect 109092 15864 117964 15892
rect 109092 15852 109098 15864
rect 117958 15852 117964 15864
rect 118016 15852 118022 15904
rect 138842 15852 138848 15904
rect 138900 15892 138906 15904
rect 417050 15892 417056 15904
rect 138900 15864 417056 15892
rect 138900 15852 138906 15864
rect 417050 15852 417056 15864
rect 417108 15852 417114 15904
rect 234614 14968 234620 15020
rect 234672 15008 234678 15020
rect 443086 15008 443092 15020
rect 234672 14980 443092 15008
rect 234672 14968 234678 14980
rect 443086 14968 443092 14980
rect 443144 14968 443150 15020
rect 231026 14900 231032 14952
rect 231084 14940 231090 14952
rect 443270 14940 443276 14952
rect 231084 14912 443276 14940
rect 231084 14900 231090 14912
rect 443270 14900 443276 14912
rect 443328 14900 443334 14952
rect 227530 14832 227536 14884
rect 227588 14872 227594 14884
rect 441614 14872 441620 14884
rect 227588 14844 441620 14872
rect 227588 14832 227594 14844
rect 441614 14832 441620 14844
rect 441672 14832 441678 14884
rect 223574 14764 223580 14816
rect 223632 14804 223638 14816
rect 440510 14804 440516 14816
rect 223632 14776 440516 14804
rect 223632 14764 223638 14776
rect 440510 14764 440516 14776
rect 440568 14764 440574 14816
rect 219986 14696 219992 14748
rect 220044 14736 220050 14748
rect 440326 14736 440332 14748
rect 220044 14708 440332 14736
rect 220044 14696 220050 14708
rect 440326 14696 440332 14708
rect 440384 14696 440390 14748
rect 216858 14628 216864 14680
rect 216916 14668 216922 14680
rect 438854 14668 438860 14680
rect 216916 14640 438860 14668
rect 216916 14628 216922 14640
rect 438854 14628 438860 14640
rect 438912 14628 438918 14680
rect 213362 14560 213368 14612
rect 213420 14600 213426 14612
rect 437566 14600 437572 14612
rect 213420 14572 437572 14600
rect 213420 14560 213426 14572
rect 437566 14560 437572 14572
rect 437624 14560 437630 14612
rect 493042 14560 493048 14612
rect 493100 14600 493106 14612
rect 514754 14600 514760 14612
rect 493100 14572 514760 14600
rect 493100 14560 493106 14572
rect 514754 14560 514760 14572
rect 514812 14560 514818 14612
rect 73338 14492 73344 14544
rect 73396 14532 73402 14544
rect 108482 14532 108488 14544
rect 73396 14504 108488 14532
rect 73396 14492 73402 14504
rect 108482 14492 108488 14504
rect 108540 14492 108546 14544
rect 147122 14492 147128 14544
rect 147180 14532 147186 14544
rect 166258 14532 166264 14544
rect 147180 14504 166264 14532
rect 147180 14492 147186 14504
rect 166258 14492 166264 14504
rect 166316 14492 166322 14544
rect 209774 14492 209780 14544
rect 209832 14532 209838 14544
rect 436186 14532 436192 14544
rect 209832 14504 436192 14532
rect 209832 14492 209838 14504
rect 436186 14492 436192 14504
rect 436244 14492 436250 14544
rect 33594 14424 33600 14476
rect 33652 14464 33658 14476
rect 65518 14464 65524 14476
rect 33652 14436 65524 14464
rect 33652 14424 33658 14436
rect 65518 14424 65524 14436
rect 65576 14424 65582 14476
rect 99834 14424 99840 14476
rect 99892 14464 99898 14476
rect 146938 14464 146944 14476
rect 99892 14436 146944 14464
rect 99892 14424 99898 14436
rect 146938 14424 146944 14436
rect 146996 14424 147002 14476
rect 206186 14424 206192 14476
rect 206244 14464 206250 14476
rect 436370 14464 436376 14476
rect 206244 14436 436376 14464
rect 206244 14424 206250 14436
rect 436370 14424 436376 14436
rect 436428 14424 436434 14476
rect 440878 14424 440884 14476
rect 440936 14464 440942 14476
rect 492950 14464 492956 14476
rect 440936 14436 492956 14464
rect 440936 14424 440942 14436
rect 492950 14424 492956 14436
rect 493008 14424 493014 14476
rect 158898 13404 158904 13456
rect 158956 13444 158962 13456
rect 293402 13444 293408 13456
rect 158956 13416 293408 13444
rect 158956 13404 158962 13416
rect 293402 13404 293408 13416
rect 293460 13404 293466 13456
rect 301498 13404 301504 13456
rect 301556 13444 301562 13456
rect 462406 13444 462412 13456
rect 301556 13416 462412 13444
rect 301556 13404 301562 13416
rect 462406 13404 462412 13416
rect 462464 13404 462470 13456
rect 155126 13336 155132 13388
rect 155184 13376 155190 13388
rect 293218 13376 293224 13388
rect 155184 13348 293224 13376
rect 155184 13336 155190 13348
rect 293218 13336 293224 13348
rect 293276 13336 293282 13388
rect 298094 13336 298100 13388
rect 298152 13376 298158 13388
rect 460934 13376 460940 13388
rect 298152 13348 460940 13376
rect 298152 13336 298158 13348
rect 460934 13336 460940 13348
rect 460992 13336 460998 13388
rect 151814 13268 151820 13320
rect 151872 13308 151878 13320
rect 291838 13308 291844 13320
rect 151872 13280 291844 13308
rect 151872 13268 151878 13280
rect 291838 13268 291844 13280
rect 291896 13268 291902 13320
rect 294874 13268 294880 13320
rect 294932 13308 294938 13320
rect 459830 13308 459836 13320
rect 294932 13280 459836 13308
rect 294932 13268 294938 13280
rect 459830 13268 459836 13280
rect 459888 13268 459894 13320
rect 291378 13200 291384 13252
rect 291436 13240 291442 13252
rect 459646 13240 459652 13252
rect 291436 13212 459652 13240
rect 291436 13200 291442 13212
rect 459646 13200 459652 13212
rect 459704 13200 459710 13252
rect 163682 13132 163688 13184
rect 163740 13172 163746 13184
rect 423950 13172 423956 13184
rect 163740 13144 423956 13172
rect 163740 13132 163746 13144
rect 423950 13132 423956 13144
rect 424008 13132 424014 13184
rect 21818 13064 21824 13116
rect 21876 13104 21882 13116
rect 62758 13104 62764 13116
rect 21876 13076 62764 13104
rect 21876 13064 21882 13076
rect 62758 13064 62764 13076
rect 62816 13064 62822 13116
rect 65058 13064 65064 13116
rect 65116 13104 65122 13116
rect 75362 13104 75368 13116
rect 65116 13076 75368 13104
rect 65116 13064 65122 13076
rect 75362 13064 75368 13076
rect 75420 13064 75426 13116
rect 89438 13064 89444 13116
rect 89496 13104 89502 13116
rect 118786 13104 118792 13116
rect 89496 13076 118792 13104
rect 89496 13064 89502 13076
rect 118786 13064 118792 13076
rect 118844 13064 118850 13116
rect 127526 13064 127532 13116
rect 127584 13104 127590 13116
rect 414014 13104 414020 13116
rect 127584 13076 414020 13104
rect 127584 13064 127590 13076
rect 414014 13064 414020 13076
rect 414072 13064 414078 13116
rect 486418 13064 486424 13116
rect 486476 13104 486482 13116
rect 513466 13104 513472 13116
rect 486476 13076 513472 13104
rect 486476 13064 486482 13076
rect 513466 13064 513472 13076
rect 513524 13064 513530 13116
rect 258258 12044 258264 12096
rect 258316 12084 258322 12096
rect 325694 12084 325700 12096
rect 258316 12056 325700 12084
rect 258316 12044 258322 12056
rect 325694 12044 325700 12056
rect 325752 12044 325758 12096
rect 254210 11976 254216 12028
rect 254268 12016 254274 12028
rect 324498 12016 324504 12028
rect 254268 11988 324504 12016
rect 254268 11976 254274 11988
rect 324498 11976 324504 11988
rect 324556 11976 324562 12028
rect 251266 11908 251272 11960
rect 251324 11948 251330 11960
rect 324682 11948 324688 11960
rect 251324 11920 324688 11948
rect 251324 11908 251330 11920
rect 324682 11908 324688 11920
rect 324740 11908 324746 11960
rect 240134 11840 240140 11892
rect 240192 11880 240198 11892
rect 321738 11880 321744 11892
rect 240192 11852 321744 11880
rect 240192 11840 240198 11852
rect 321738 11840 321744 11852
rect 321796 11840 321802 11892
rect 386690 11840 386696 11892
rect 386748 11880 386754 11892
rect 485958 11880 485964 11892
rect 386748 11852 485964 11880
rect 386748 11840 386754 11852
rect 485958 11840 485964 11852
rect 486016 11840 486022 11892
rect 61562 11772 61568 11824
rect 61620 11812 61626 11824
rect 73798 11812 73804 11824
rect 61620 11784 73804 11812
rect 61620 11772 61626 11784
rect 73798 11772 73804 11784
rect 73856 11772 73862 11824
rect 218054 11772 218060 11824
rect 218112 11812 218118 11824
rect 219250 11812 219256 11824
rect 218112 11784 219256 11812
rect 218112 11772 218118 11784
rect 219250 11772 219256 11784
rect 219308 11772 219314 11824
rect 233418 11772 233424 11824
rect 233476 11812 233482 11824
rect 318794 11812 318800 11824
rect 233476 11784 318800 11812
rect 233476 11772 233482 11784
rect 318794 11772 318800 11784
rect 318852 11772 318858 11824
rect 324406 11772 324412 11824
rect 324464 11812 324470 11824
rect 343818 11812 343824 11824
rect 324464 11784 343824 11812
rect 324464 11772 324470 11784
rect 343818 11772 343824 11784
rect 343876 11772 343882 11824
rect 357434 11772 357440 11824
rect 357492 11812 357498 11824
rect 477586 11812 477592 11824
rect 357492 11784 477592 11812
rect 357492 11772 357498 11784
rect 477586 11772 477592 11784
rect 477644 11772 477650 11824
rect 11606 11704 11612 11756
rect 11664 11744 11670 11756
rect 61378 11744 61384 11756
rect 11664 11716 61384 11744
rect 11664 11704 11670 11716
rect 61378 11704 61384 11716
rect 61436 11704 61442 11756
rect 89622 11704 89628 11756
rect 89680 11744 89686 11756
rect 114738 11744 114744 11756
rect 89680 11716 114744 11744
rect 89680 11704 89686 11716
rect 114738 11704 114744 11716
rect 114796 11704 114802 11756
rect 133874 11704 133880 11756
rect 133932 11744 133938 11756
rect 286502 11744 286508 11756
rect 133932 11716 286508 11744
rect 133932 11704 133938 11716
rect 286502 11704 286508 11716
rect 286560 11704 286566 11756
rect 322934 11704 322940 11756
rect 322992 11744 322998 11756
rect 467834 11744 467840 11756
rect 322992 11716 467840 11744
rect 322992 11704 322998 11716
rect 467834 11704 467840 11716
rect 467892 11704 467898 11756
rect 490006 11704 490012 11756
rect 490064 11744 490070 11756
rect 513650 11744 513656 11756
rect 490064 11716 513656 11744
rect 490064 11704 490070 11716
rect 513650 11704 513656 11716
rect 513708 11704 513714 11756
rect 259454 11636 259460 11688
rect 259512 11676 259518 11688
rect 260650 11676 260656 11688
rect 259512 11648 260656 11676
rect 259512 11636 259518 11648
rect 260650 11636 260656 11648
rect 260708 11636 260714 11688
rect 374638 10752 374644 10804
rect 374696 10792 374702 10804
rect 432046 10792 432052 10804
rect 374696 10764 432052 10792
rect 374696 10752 374702 10764
rect 432046 10752 432052 10764
rect 432104 10752 432110 10804
rect 186866 10684 186872 10736
rect 186924 10724 186930 10736
rect 306374 10724 306380 10736
rect 186924 10696 306380 10724
rect 186924 10684 186930 10696
rect 306374 10684 306380 10696
rect 306432 10684 306438 10736
rect 374822 10684 374828 10736
rect 374880 10724 374886 10736
rect 435082 10724 435088 10736
rect 374880 10696 435088 10724
rect 374880 10684 374886 10696
rect 435082 10684 435088 10696
rect 435140 10684 435146 10736
rect 183738 10616 183744 10668
rect 183796 10656 183802 10668
rect 305270 10656 305276 10668
rect 183796 10628 305276 10656
rect 183796 10616 183802 10628
rect 305270 10616 305276 10628
rect 305328 10616 305334 10668
rect 376018 10616 376024 10668
rect 376076 10656 376082 10668
rect 439130 10656 439136 10668
rect 376076 10628 439136 10656
rect 376076 10616 376082 10628
rect 439130 10616 439136 10628
rect 439188 10616 439194 10668
rect 180242 10548 180248 10600
rect 180300 10588 180306 10600
rect 305086 10588 305092 10600
rect 180300 10560 305092 10588
rect 180300 10548 180306 10560
rect 305086 10548 305092 10560
rect 305144 10548 305150 10600
rect 377398 10548 377404 10600
rect 377456 10588 377462 10600
rect 442626 10588 442632 10600
rect 377456 10560 442632 10588
rect 377456 10548 377462 10560
rect 442626 10548 442632 10560
rect 442684 10548 442690 10600
rect 169570 10480 169576 10532
rect 169628 10520 169634 10532
rect 296162 10520 296168 10532
rect 169628 10492 296168 10520
rect 169628 10480 169634 10492
rect 296162 10480 296168 10492
rect 296220 10480 296226 10532
rect 339586 10480 339592 10532
rect 339644 10520 339650 10532
rect 347958 10520 347964 10532
rect 339644 10492 347964 10520
rect 339644 10480 339650 10492
rect 347958 10480 347964 10492
rect 348016 10480 348022 10532
rect 377582 10480 377588 10532
rect 377640 10520 377646 10532
rect 445754 10520 445760 10532
rect 377640 10492 445760 10520
rect 377640 10480 377646 10492
rect 445754 10480 445760 10492
rect 445812 10480 445818 10532
rect 172698 10412 172704 10464
rect 172756 10452 172762 10464
rect 302234 10452 302240 10464
rect 172756 10424 302240 10452
rect 172756 10412 172762 10424
rect 302234 10412 302240 10424
rect 302292 10412 302298 10464
rect 332686 10412 332692 10464
rect 332744 10452 332750 10464
rect 346486 10452 346492 10464
rect 332744 10424 346492 10452
rect 332744 10412 332750 10424
rect 346486 10412 346492 10424
rect 346544 10412 346550 10464
rect 378778 10412 378784 10464
rect 378836 10452 378842 10464
rect 448514 10452 448520 10464
rect 378836 10424 448520 10452
rect 378836 10412 378842 10424
rect 448514 10412 448520 10424
rect 448572 10412 448578 10464
rect 84102 10344 84108 10396
rect 84160 10384 84166 10396
rect 97442 10384 97448 10396
rect 84160 10356 97448 10384
rect 84160 10344 84166 10356
rect 97442 10344 97448 10356
rect 97500 10344 97506 10396
rect 166074 10344 166080 10396
rect 166132 10384 166138 10396
rect 295978 10384 295984 10396
rect 166132 10356 295984 10384
rect 166132 10344 166138 10356
rect 295978 10344 295984 10356
rect 296036 10344 296042 10396
rect 307938 10344 307944 10396
rect 307996 10384 308002 10396
rect 339494 10384 339500 10396
rect 307996 10356 339500 10384
rect 307996 10344 308002 10356
rect 339494 10344 339500 10356
rect 339552 10344 339558 10396
rect 381722 10344 381728 10396
rect 381780 10384 381786 10396
rect 456886 10384 456892 10396
rect 381780 10356 456892 10384
rect 381780 10344 381786 10356
rect 456886 10344 456892 10356
rect 456944 10344 456950 10396
rect 51074 10276 51080 10328
rect 51132 10316 51138 10328
rect 71038 10316 71044 10328
rect 51132 10288 71044 10316
rect 51132 10276 51138 10288
rect 71038 10276 71044 10288
rect 71096 10276 71102 10328
rect 84194 10276 84200 10328
rect 84252 10316 84258 10328
rect 111058 10316 111064 10328
rect 84252 10288 111064 10316
rect 84252 10276 84258 10288
rect 111058 10276 111064 10288
rect 111116 10276 111122 10328
rect 130286 10276 130292 10328
rect 130344 10316 130350 10328
rect 286318 10316 286324 10328
rect 130344 10288 286324 10316
rect 130344 10276 130350 10288
rect 286318 10276 286324 10288
rect 286376 10276 286382 10328
rect 297266 10276 297272 10328
rect 297324 10316 297330 10328
rect 336734 10316 336740 10328
rect 297324 10288 336740 10316
rect 297324 10276 297330 10288
rect 336734 10276 336740 10288
rect 336792 10276 336798 10328
rect 355318 10276 355324 10328
rect 355376 10316 355382 10328
rect 364610 10316 364616 10328
rect 355376 10288 364616 10316
rect 355376 10276 355382 10288
rect 364610 10276 364616 10288
rect 364668 10276 364674 10328
rect 381538 10276 381544 10328
rect 381596 10316 381602 10328
rect 459922 10316 459928 10328
rect 381596 10288 459928 10316
rect 381596 10276 381602 10288
rect 459922 10276 459928 10288
rect 459980 10276 459986 10328
rect 482370 10276 482376 10328
rect 482428 10316 482434 10328
rect 511994 10316 512000 10328
rect 482428 10288 512000 10316
rect 482428 10276 482434 10288
rect 511994 10276 512000 10288
rect 512052 10276 512058 10328
rect 429654 9256 429660 9308
rect 429712 9296 429718 9308
rect 496906 9296 496912 9308
rect 429712 9268 496912 9296
rect 429712 9256 429718 9268
rect 496906 9256 496912 9268
rect 496964 9256 496970 9308
rect 412266 9188 412272 9240
rect 412324 9228 412330 9240
rect 492766 9228 492772 9240
rect 412324 9200 492772 9228
rect 412324 9188 412330 9200
rect 492766 9188 492772 9200
rect 492824 9188 492830 9240
rect 394234 9120 394240 9172
rect 394292 9160 394298 9172
rect 487246 9160 487252 9172
rect 394292 9132 487252 9160
rect 394292 9120 394298 9132
rect 487246 9120 487252 9132
rect 487304 9120 487310 9172
rect 180702 9052 180708 9104
rect 180760 9092 180766 9104
rect 196802 9092 196808 9104
rect 180760 9064 196808 9092
rect 180760 9052 180766 9064
rect 196802 9052 196808 9064
rect 196860 9052 196866 9104
rect 246666 9052 246672 9104
rect 246724 9092 246730 9104
rect 441522 9092 441528 9104
rect 246724 9064 441528 9092
rect 246724 9052 246730 9064
rect 441522 9052 441528 9064
rect 441580 9052 441586 9104
rect 86862 8984 86868 9036
rect 86920 9024 86926 9036
rect 108114 9024 108120 9036
rect 86920 8996 108120 9024
rect 86920 8984 86926 8996
rect 108114 8984 108120 8996
rect 108172 8984 108178 9036
rect 143626 8984 143632 9036
rect 143684 9024 143690 9036
rect 165062 9024 165068 9036
rect 143684 8996 165068 9024
rect 143684 8984 143690 8996
rect 165062 8984 165068 8996
rect 165120 8984 165126 9036
rect 184566 8984 184572 9036
rect 184624 9024 184630 9036
rect 211062 9024 211068 9036
rect 184624 8996 211068 9024
rect 184624 8984 184630 8996
rect 211062 8984 211068 8996
rect 211120 8984 211126 9036
rect 249702 8984 249708 9036
rect 249760 9024 249766 9036
rect 448606 9024 448612 9036
rect 249760 8996 448612 9024
rect 249760 8984 249766 8996
rect 448606 8984 448612 8996
rect 448664 8984 448670 9036
rect 47854 8916 47860 8968
rect 47912 8956 47918 8968
rect 69658 8956 69664 8968
rect 47912 8928 69664 8956
rect 47912 8916 47918 8928
rect 69658 8916 69664 8928
rect 69716 8916 69722 8968
rect 96246 8916 96252 8968
rect 96304 8956 96310 8968
rect 145558 8956 145564 8968
rect 96304 8928 145564 8956
rect 96304 8916 96310 8928
rect 145558 8916 145564 8928
rect 145616 8916 145622 8968
rect 193122 8916 193128 8968
rect 193180 8956 193186 8968
rect 242894 8956 242900 8968
rect 193180 8928 242900 8956
rect 193180 8916 193186 8928
rect 242894 8916 242900 8928
rect 242952 8916 242958 8968
rect 250806 8916 250812 8968
rect 250864 8956 250870 8968
rect 452102 8956 452108 8968
rect 250864 8928 452108 8956
rect 250864 8916 250870 8928
rect 452102 8916 452108 8928
rect 452160 8916 452166 8968
rect 461578 8916 461584 8968
rect 461636 8956 461642 8968
rect 506566 8956 506572 8968
rect 461636 8928 506572 8956
rect 461636 8916 461642 8928
rect 506566 8916 506572 8928
rect 506624 8916 506630 8968
rect 69106 8304 69112 8356
rect 69164 8344 69170 8356
rect 75178 8344 75184 8356
rect 69164 8316 75184 8344
rect 69164 8304 69170 8316
rect 75178 8304 75184 8316
rect 75236 8304 75242 8356
rect 81342 8304 81348 8356
rect 81400 8344 81406 8356
rect 86862 8344 86868 8356
rect 81400 8316 86868 8344
rect 81400 8304 81406 8316
rect 86862 8304 86868 8316
rect 86920 8304 86926 8356
rect 79962 8236 79968 8288
rect 80020 8276 80026 8288
rect 83274 8276 83280 8288
rect 80020 8248 83280 8276
rect 80020 8236 80026 8248
rect 83274 8236 83280 8248
rect 83332 8236 83338 8288
rect 369118 8236 369124 8288
rect 369176 8276 369182 8288
rect 414290 8276 414296 8288
rect 369176 8248 414296 8276
rect 369176 8236 369182 8248
rect 414290 8236 414296 8248
rect 414348 8236 414354 8288
rect 370498 8168 370504 8220
rect 370556 8208 370562 8220
rect 417878 8208 417884 8220
rect 370556 8180 417884 8208
rect 370556 8168 370562 8180
rect 417878 8168 417884 8180
rect 417936 8168 417942 8220
rect 422570 8168 422576 8220
rect 422628 8208 422634 8220
rect 495526 8208 495532 8220
rect 422628 8180 495532 8208
rect 422628 8168 422634 8180
rect 495526 8168 495532 8180
rect 495584 8168 495590 8220
rect 406378 8100 406384 8152
rect 406436 8140 406442 8152
rect 549070 8140 549076 8152
rect 406436 8112 549076 8140
rect 406436 8100 406442 8112
rect 549070 8100 549076 8112
rect 549128 8100 549134 8152
rect 407942 8032 407948 8084
rect 408000 8072 408006 8084
rect 552658 8072 552664 8084
rect 408000 8044 552664 8072
rect 408000 8032 408006 8044
rect 552658 8032 552664 8044
rect 552716 8032 552722 8084
rect 407758 7964 407764 8016
rect 407816 8004 407822 8016
rect 556154 8004 556160 8016
rect 407816 7976 556160 8004
rect 407816 7964 407822 7976
rect 556154 7964 556160 7976
rect 556212 7964 556218 8016
rect 365162 7896 365168 7948
rect 365220 7936 365226 7948
rect 400122 7936 400128 7948
rect 365220 7908 400128 7936
rect 365220 7896 365226 7908
rect 400122 7896 400128 7908
rect 400180 7896 400186 7948
rect 409138 7896 409144 7948
rect 409196 7936 409202 7948
rect 559742 7936 559748 7948
rect 409196 7908 559748 7936
rect 409196 7896 409202 7908
rect 559742 7896 559748 7908
rect 559800 7896 559806 7948
rect 366358 7828 366364 7880
rect 366416 7868 366422 7880
rect 403710 7868 403716 7880
rect 366416 7840 403716 7868
rect 366416 7828 366422 7840
rect 403710 7828 403716 7840
rect 403768 7828 403774 7880
rect 410702 7828 410708 7880
rect 410760 7868 410766 7880
rect 563238 7868 563244 7880
rect 410760 7840 563244 7868
rect 410760 7828 410766 7840
rect 563238 7828 563244 7840
rect 563296 7828 563302 7880
rect 367738 7760 367744 7812
rect 367796 7800 367802 7812
rect 407206 7800 407212 7812
rect 367796 7772 407212 7800
rect 367796 7760 367802 7772
rect 407206 7760 407212 7772
rect 407264 7760 407270 7812
rect 410518 7760 410524 7812
rect 410576 7800 410582 7812
rect 566826 7800 566832 7812
rect 410576 7772 566832 7800
rect 410576 7760 410582 7772
rect 566826 7760 566832 7772
rect 566884 7760 566890 7812
rect 179322 7692 179328 7744
rect 179380 7732 179386 7744
rect 193306 7732 193312 7744
rect 179380 7704 193312 7732
rect 179380 7692 179386 7704
rect 193306 7692 193312 7704
rect 193364 7692 193370 7744
rect 244090 7692 244096 7744
rect 244148 7732 244154 7744
rect 321922 7732 321928 7744
rect 244148 7704 321928 7732
rect 244148 7692 244154 7704
rect 321922 7692 321928 7704
rect 321980 7692 321986 7744
rect 329190 7692 329196 7744
rect 329248 7732 329254 7744
rect 345106 7732 345112 7744
rect 329248 7704 345112 7732
rect 329248 7692 329254 7704
rect 345106 7692 345112 7704
rect 345164 7692 345170 7744
rect 367922 7692 367928 7744
rect 367980 7732 367986 7744
rect 410794 7732 410800 7744
rect 367980 7704 410800 7732
rect 367980 7692 367986 7704
rect 410794 7692 410800 7704
rect 410852 7692 410858 7744
rect 411898 7692 411904 7744
rect 411956 7732 411962 7744
rect 570322 7732 570328 7744
rect 411956 7704 570328 7732
rect 411956 7692 411962 7704
rect 570322 7692 570328 7704
rect 570380 7692 570386 7744
rect 58434 7624 58440 7676
rect 58492 7664 58498 7676
rect 72418 7664 72424 7676
rect 58492 7636 72424 7664
rect 58492 7624 58498 7636
rect 72418 7624 72424 7636
rect 72476 7624 72482 7676
rect 82538 7624 82544 7676
rect 82596 7664 82602 7676
rect 93946 7664 93952 7676
rect 82596 7636 93952 7664
rect 82596 7624 82602 7636
rect 93946 7624 93952 7636
rect 94004 7624 94010 7676
rect 136450 7624 136456 7676
rect 136508 7664 136514 7676
rect 163498 7664 163504 7676
rect 136508 7636 163504 7664
rect 136508 7624 136514 7636
rect 163498 7624 163504 7636
rect 163556 7624 163562 7676
rect 181990 7624 181996 7676
rect 182048 7664 182054 7676
rect 203886 7664 203892 7676
rect 182048 7636 203892 7664
rect 182048 7624 182054 7636
rect 203886 7624 203892 7636
rect 203944 7624 203950 7676
rect 229002 7624 229008 7676
rect 229060 7664 229066 7676
rect 374086 7664 374092 7676
rect 229060 7636 374092 7664
rect 229060 7624 229066 7636
rect 374086 7624 374092 7636
rect 374144 7624 374150 7676
rect 413278 7624 413284 7676
rect 413336 7664 413342 7676
rect 573910 7664 573916 7676
rect 413336 7636 573916 7664
rect 413336 7624 413342 7636
rect 573910 7624 573916 7636
rect 573968 7624 573974 7676
rect 2866 7556 2872 7608
rect 2924 7596 2930 7608
rect 58618 7596 58624 7608
rect 2924 7568 58624 7596
rect 2924 7556 2930 7568
rect 58618 7556 58624 7568
rect 58676 7556 58682 7608
rect 88242 7556 88248 7608
rect 88300 7596 88306 7608
rect 111610 7596 111616 7608
rect 88300 7568 111616 7596
rect 88300 7556 88306 7568
rect 111610 7556 111616 7568
rect 111668 7556 111674 7608
rect 117590 7556 117596 7608
rect 117648 7596 117654 7608
rect 151078 7596 151084 7608
rect 117648 7568 151084 7596
rect 117648 7556 117654 7568
rect 151078 7556 151084 7568
rect 151136 7556 151142 7608
rect 157794 7556 157800 7608
rect 157852 7596 157858 7608
rect 169018 7596 169024 7608
rect 157852 7568 169024 7596
rect 157852 7556 157858 7568
rect 169018 7556 169024 7568
rect 169076 7556 169082 7608
rect 187326 7556 187332 7608
rect 187384 7596 187390 7608
rect 221550 7596 221556 7608
rect 187384 7568 221556 7596
rect 187384 7556 187390 7568
rect 221550 7556 221556 7568
rect 221608 7556 221614 7608
rect 231762 7556 231768 7608
rect 231820 7596 231826 7608
rect 384758 7596 384764 7608
rect 231820 7568 384764 7596
rect 231820 7556 231826 7568
rect 384758 7556 384764 7568
rect 384816 7556 384822 7608
rect 414658 7556 414664 7608
rect 414716 7596 414722 7608
rect 577406 7596 577412 7608
rect 414716 7568 577412 7596
rect 414716 7556 414722 7568
rect 577406 7556 577412 7568
rect 577464 7556 577470 7608
rect 72602 6876 72608 6928
rect 72660 6916 72666 6928
rect 76558 6916 76564 6928
rect 72660 6888 76564 6916
rect 72660 6876 72666 6888
rect 76558 6876 76564 6888
rect 76616 6876 76622 6928
rect 41874 6672 41880 6724
rect 41932 6712 41938 6724
rect 100018 6712 100024 6724
rect 41932 6684 100024 6712
rect 41932 6672 41938 6684
rect 100018 6672 100024 6684
rect 100076 6672 100082 6724
rect 300762 6672 300768 6724
rect 300820 6712 300826 6724
rect 338482 6712 338488 6724
rect 300820 6684 338488 6712
rect 300820 6672 300826 6684
rect 338482 6672 338488 6684
rect 338540 6672 338546 6724
rect 356698 6672 356704 6724
rect 356756 6712 356762 6724
rect 368198 6712 368204 6724
rect 356756 6684 368204 6712
rect 356756 6672 356762 6684
rect 368198 6672 368204 6684
rect 368256 6672 368262 6724
rect 34790 6604 34796 6656
rect 34848 6644 34854 6656
rect 98638 6644 98644 6656
rect 34848 6616 98644 6644
rect 34848 6604 34854 6616
rect 98638 6604 98644 6616
rect 98696 6604 98702 6656
rect 286594 6604 286600 6656
rect 286652 6644 286658 6656
rect 334342 6644 334348 6656
rect 286652 6616 334348 6644
rect 286652 6604 286658 6616
rect 334342 6604 334348 6616
rect 334400 6604 334406 6656
rect 358262 6604 358268 6656
rect 358320 6644 358326 6656
rect 371694 6644 371700 6656
rect 358320 6616 371700 6644
rect 358320 6604 358326 6616
rect 371694 6604 371700 6616
rect 371752 6604 371758 6656
rect 74994 6536 75000 6588
rect 75052 6576 75058 6588
rect 140038 6576 140044 6588
rect 75052 6548 140044 6576
rect 75052 6536 75058 6548
rect 140038 6536 140044 6548
rect 140096 6536 140102 6588
rect 205542 6536 205548 6588
rect 205600 6576 205606 6588
rect 288986 6576 288992 6588
rect 205600 6548 288992 6576
rect 205600 6536 205606 6548
rect 288986 6536 288992 6548
rect 289044 6536 289050 6588
rect 290182 6536 290188 6588
rect 290240 6576 290246 6588
rect 334158 6576 334164 6588
rect 290240 6548 334164 6576
rect 290240 6536 290246 6548
rect 334158 6536 334164 6548
rect 334216 6536 334222 6588
rect 358078 6536 358084 6588
rect 358136 6576 358142 6588
rect 375282 6576 375288 6588
rect 358136 6548 375288 6576
rect 358136 6536 358142 6548
rect 375282 6536 375288 6548
rect 375340 6536 375346 6588
rect 27706 6468 27712 6520
rect 27764 6508 27770 6520
rect 95878 6508 95884 6520
rect 27764 6480 95884 6508
rect 27764 6468 27770 6480
rect 95878 6468 95884 6480
rect 95936 6468 95942 6520
rect 206922 6468 206928 6520
rect 206980 6508 206986 6520
rect 292574 6508 292580 6520
rect 206980 6480 292580 6508
rect 206980 6468 206986 6480
rect 292574 6468 292580 6480
rect 292632 6468 292638 6520
rect 293678 6468 293684 6520
rect 293736 6508 293742 6520
rect 335446 6508 335452 6520
rect 293736 6480 335452 6508
rect 293736 6468 293742 6480
rect 335446 6468 335452 6480
rect 335504 6468 335510 6520
rect 359550 6468 359556 6520
rect 359608 6508 359614 6520
rect 378870 6508 378876 6520
rect 359608 6480 378876 6508
rect 359608 6468 359614 6480
rect 378870 6468 378876 6480
rect 378928 6468 378934 6520
rect 388622 6468 388628 6520
rect 388680 6508 388686 6520
rect 481726 6508 481732 6520
rect 388680 6480 481732 6508
rect 388680 6468 388686 6480
rect 481726 6468 481732 6480
rect 481784 6468 481790 6520
rect 64322 6400 64328 6452
rect 64380 6440 64386 6452
rect 137278 6440 137284 6452
rect 64380 6412 137284 6440
rect 64380 6400 64386 6412
rect 137278 6400 137284 6412
rect 137336 6400 137342 6452
rect 209682 6400 209688 6452
rect 209740 6440 209746 6452
rect 303154 6440 303160 6452
rect 209740 6412 303160 6440
rect 209740 6400 209746 6412
rect 303154 6400 303160 6412
rect 303212 6400 303218 6452
rect 304350 6400 304356 6452
rect 304408 6440 304414 6452
rect 338298 6440 338304 6452
rect 304408 6412 338304 6440
rect 304408 6400 304414 6412
rect 338298 6400 338304 6412
rect 338356 6400 338362 6452
rect 360838 6400 360844 6452
rect 360896 6440 360902 6452
rect 382366 6440 382372 6452
rect 360896 6412 382372 6440
rect 360896 6400 360902 6412
rect 382366 6400 382372 6412
rect 382424 6400 382430 6452
rect 388438 6400 388444 6452
rect 388496 6440 388502 6452
rect 485222 6440 485228 6452
rect 388496 6412 485228 6440
rect 388496 6400 388502 6412
rect 485222 6400 485228 6412
rect 485280 6400 485286 6452
rect 53742 6332 53748 6384
rect 53800 6372 53806 6384
rect 134518 6372 134524 6384
rect 53800 6344 134524 6372
rect 53800 6332 53806 6344
rect 134518 6332 134524 6344
rect 134576 6332 134582 6384
rect 210786 6332 210792 6384
rect 210844 6372 210850 6384
rect 306742 6372 306748 6384
rect 210844 6344 306748 6372
rect 210844 6332 210850 6344
rect 306742 6332 306748 6344
rect 306800 6332 306806 6384
rect 361022 6332 361028 6384
rect 361080 6372 361086 6384
rect 385954 6372 385960 6384
rect 361080 6344 385960 6372
rect 361080 6332 361086 6344
rect 385954 6332 385960 6344
rect 386012 6332 386018 6384
rect 389818 6332 389824 6384
rect 389876 6372 389882 6384
rect 488810 6372 488816 6384
rect 389876 6344 488816 6372
rect 389876 6332 389882 6344
rect 488810 6332 488816 6344
rect 488868 6332 488874 6384
rect 50154 6264 50160 6316
rect 50212 6304 50218 6316
rect 133138 6304 133144 6316
rect 50212 6276 133144 6304
rect 50212 6264 50218 6276
rect 133138 6264 133144 6276
rect 133196 6264 133202 6316
rect 177758 6264 177764 6316
rect 177816 6304 177822 6316
rect 186130 6304 186136 6316
rect 177816 6276 186136 6304
rect 177816 6264 177822 6276
rect 186130 6264 186136 6276
rect 186188 6264 186194 6316
rect 210970 6264 210976 6316
rect 211028 6304 211034 6316
rect 310238 6304 310244 6316
rect 211028 6276 310244 6304
rect 211028 6264 211034 6276
rect 310238 6264 310244 6276
rect 310296 6264 310302 6316
rect 311434 6264 311440 6316
rect 311492 6304 311498 6316
rect 340966 6304 340972 6316
rect 311492 6276 340972 6304
rect 311492 6264 311498 6276
rect 340966 6264 340972 6276
rect 341024 6264 341030 6316
rect 343358 6264 343364 6316
rect 343416 6304 343422 6316
rect 349338 6304 349344 6316
rect 343416 6276 349344 6304
rect 343416 6264 343422 6276
rect 349338 6264 349344 6276
rect 349396 6264 349402 6316
rect 362218 6264 362224 6316
rect 362276 6304 362282 6316
rect 389450 6304 389456 6316
rect 362276 6276 389456 6304
rect 362276 6264 362282 6276
rect 389450 6264 389456 6276
rect 389508 6264 389514 6316
rect 394142 6264 394148 6316
rect 394200 6304 394206 6316
rect 502978 6304 502984 6316
rect 394200 6276 502984 6304
rect 394200 6264 394206 6276
rect 502978 6264 502984 6276
rect 503036 6264 503042 6316
rect 14734 6196 14740 6248
rect 14792 6236 14798 6248
rect 125042 6236 125048 6248
rect 14792 6208 125048 6236
rect 14792 6196 14798 6208
rect 125042 6196 125048 6208
rect 125100 6196 125106 6248
rect 161290 6196 161296 6248
rect 161348 6236 161354 6248
rect 170582 6236 170588 6248
rect 161348 6208 170588 6236
rect 161348 6196 161354 6208
rect 170582 6196 170588 6208
rect 170640 6196 170646 6248
rect 181806 6196 181812 6248
rect 181864 6236 181870 6248
rect 200298 6236 200304 6248
rect 181864 6208 200304 6236
rect 181864 6196 181870 6208
rect 200298 6196 200304 6208
rect 200356 6196 200362 6248
rect 212442 6196 212448 6248
rect 212500 6236 212506 6248
rect 313826 6236 313832 6248
rect 212500 6208 313832 6236
rect 212500 6196 212506 6208
rect 313826 6196 313832 6208
rect 313884 6196 313890 6248
rect 363598 6196 363604 6248
rect 363656 6236 363662 6248
rect 393038 6236 393044 6248
rect 363656 6208 393044 6236
rect 363656 6196 363662 6208
rect 393038 6196 393044 6208
rect 393096 6196 393102 6248
rect 393958 6196 393964 6248
rect 394016 6236 394022 6248
rect 506474 6236 506480 6248
rect 394016 6208 506480 6236
rect 394016 6196 394022 6208
rect 506474 6196 506480 6208
rect 506532 6196 506538 6248
rect 9950 6128 9956 6180
rect 10008 6168 10014 6180
rect 123478 6168 123484 6180
rect 10008 6140 123484 6168
rect 10008 6128 10014 6140
rect 123478 6128 123484 6140
rect 123536 6128 123542 6180
rect 154206 6128 154212 6180
rect 154264 6168 154270 6180
rect 167638 6168 167644 6180
rect 154264 6140 167644 6168
rect 154264 6128 154270 6140
rect 167638 6128 167644 6140
rect 167696 6128 167702 6180
rect 183462 6128 183468 6180
rect 183520 6168 183526 6180
rect 207382 6168 207388 6180
rect 183520 6140 207388 6168
rect 183520 6128 183526 6140
rect 207382 6128 207388 6140
rect 207440 6128 207446 6180
rect 213546 6128 213552 6180
rect 213604 6168 213610 6180
rect 317322 6168 317328 6180
rect 213604 6140 317328 6168
rect 213604 6128 213610 6140
rect 317322 6128 317328 6140
rect 317380 6128 317386 6180
rect 318518 6128 318524 6180
rect 318576 6168 318582 6180
rect 342254 6168 342260 6180
rect 318576 6140 342260 6168
rect 318576 6128 318582 6140
rect 342254 6128 342260 6140
rect 342312 6128 342318 6180
rect 353846 6128 353852 6180
rect 353904 6168 353910 6180
rect 357526 6168 357532 6180
rect 353904 6140 357532 6168
rect 353904 6128 353910 6140
rect 357526 6128 357532 6140
rect 357584 6128 357590 6180
rect 364978 6128 364984 6180
rect 365036 6168 365042 6180
rect 396534 6168 396540 6180
rect 365036 6140 396540 6168
rect 365036 6128 365042 6140
rect 396534 6128 396540 6140
rect 396592 6128 396598 6180
rect 396718 6128 396724 6180
rect 396776 6168 396782 6180
rect 513558 6168 513564 6180
rect 396776 6140 513564 6168
rect 396776 6128 396782 6140
rect 513558 6128 513564 6140
rect 513616 6128 513622 6180
rect 174906 5516 174912 5568
rect 174964 5556 174970 5568
rect 179046 5556 179052 5568
rect 174964 5528 179052 5556
rect 174964 5516 174970 5528
rect 179046 5516 179052 5528
rect 179104 5516 179110 5568
rect 352558 5516 352564 5568
rect 352616 5556 352622 5568
rect 354030 5556 354036 5568
rect 352616 5528 354036 5556
rect 352616 5516 352622 5528
rect 354030 5516 354036 5528
rect 354088 5516 354094 5568
rect 98638 5312 98644 5364
rect 98696 5352 98702 5364
rect 105538 5352 105544 5364
rect 98696 5324 105544 5352
rect 98696 5312 98702 5324
rect 105538 5312 105544 5324
rect 105596 5312 105602 5364
rect 102226 5244 102232 5296
rect 102284 5284 102290 5296
rect 116578 5284 116584 5296
rect 102284 5256 116584 5284
rect 102284 5244 102290 5256
rect 116578 5244 116584 5256
rect 116636 5244 116642 5296
rect 267366 5244 267372 5296
rect 267424 5284 267430 5296
rect 512454 5284 512460 5296
rect 267424 5256 512460 5284
rect 267424 5244 267430 5256
rect 512454 5244 512460 5256
rect 512512 5244 512518 5296
rect 98730 5176 98736 5228
rect 98788 5216 98794 5228
rect 115382 5216 115388 5228
rect 98788 5188 115388 5216
rect 98788 5176 98794 5188
rect 115382 5176 115388 5188
rect 115440 5176 115446 5228
rect 267550 5176 267556 5228
rect 267608 5216 267614 5228
rect 515950 5216 515956 5228
rect 267608 5188 515956 5216
rect 267608 5176 267614 5188
rect 515950 5176 515956 5188
rect 516008 5176 516014 5228
rect 44266 5108 44272 5160
rect 44324 5148 44330 5160
rect 68462 5148 68468 5160
rect 44324 5120 68468 5148
rect 44324 5108 44330 5120
rect 68462 5108 68468 5120
rect 68520 5108 68526 5160
rect 95142 5108 95148 5160
rect 95200 5148 95206 5160
rect 115198 5148 115204 5160
rect 95200 5120 115204 5148
rect 95200 5108 95206 5120
rect 115198 5108 115204 5120
rect 115256 5108 115262 5160
rect 191466 5108 191472 5160
rect 191524 5148 191530 5160
rect 235810 5148 235816 5160
rect 191524 5120 235816 5148
rect 191524 5108 191530 5120
rect 235810 5108 235816 5120
rect 235868 5108 235874 5160
rect 269022 5108 269028 5160
rect 269080 5148 269086 5160
rect 519538 5148 519544 5160
rect 269080 5120 519544 5148
rect 269080 5108 269086 5120
rect 519538 5108 519544 5120
rect 519596 5108 519602 5160
rect 40678 5040 40684 5092
rect 40736 5080 40742 5092
rect 68278 5080 68284 5092
rect 40736 5052 68284 5080
rect 40736 5040 40742 5052
rect 68278 5040 68284 5052
rect 68336 5040 68342 5092
rect 70302 5040 70308 5092
rect 70360 5080 70366 5092
rect 108298 5080 108304 5092
rect 70360 5052 108304 5080
rect 70360 5040 70366 5052
rect 108298 5040 108304 5052
rect 108356 5040 108362 5092
rect 140038 5040 140044 5092
rect 140096 5080 140102 5092
rect 164878 5080 164884 5092
rect 140096 5052 164884 5080
rect 140096 5040 140102 5052
rect 164878 5040 164884 5052
rect 164936 5040 164942 5092
rect 191650 5040 191656 5092
rect 191708 5080 191714 5092
rect 239306 5080 239312 5092
rect 191708 5052 239312 5080
rect 191708 5040 191714 5052
rect 239306 5040 239312 5052
rect 239364 5040 239370 5092
rect 270126 5040 270132 5092
rect 270184 5080 270190 5092
rect 526622 5080 526628 5092
rect 270184 5052 526628 5080
rect 270184 5040 270190 5052
rect 526622 5040 526628 5052
rect 526680 5040 526686 5092
rect 66714 4972 66720 5024
rect 66772 5012 66778 5024
rect 106918 5012 106924 5024
rect 66772 4984 106924 5012
rect 66772 4972 66778 4984
rect 106918 4972 106924 4984
rect 106976 4972 106982 5024
rect 132954 4972 132960 5024
rect 133012 5012 133018 5024
rect 162118 5012 162124 5024
rect 133012 4984 162124 5012
rect 133012 4972 133018 4984
rect 162118 4972 162124 4984
rect 162176 4972 162182 5024
rect 195882 4972 195888 5024
rect 195940 5012 195946 5024
rect 253474 5012 253480 5024
rect 195940 4984 253480 5012
rect 195940 4972 195946 4984
rect 253474 4972 253480 4984
rect 253532 4972 253538 5024
rect 271782 4972 271788 5024
rect 271840 5012 271846 5024
rect 530118 5012 530124 5024
rect 271840 4984 530124 5012
rect 271840 4972 271846 4984
rect 530118 4972 530124 4984
rect 530176 4972 530182 5024
rect 63218 4904 63224 4956
rect 63276 4944 63282 4956
rect 98638 4944 98644 4956
rect 63276 4916 98644 4944
rect 63276 4904 63282 4916
rect 98638 4904 98644 4916
rect 98696 4904 98702 4956
rect 129366 4904 129372 4956
rect 129424 4944 129430 4956
rect 160738 4944 160744 4956
rect 129424 4916 160744 4944
rect 129424 4904 129430 4916
rect 160738 4904 160744 4916
rect 160796 4904 160802 4956
rect 197262 4904 197268 4956
rect 197320 4944 197326 4956
rect 257062 4944 257068 4956
rect 197320 4916 257068 4944
rect 197320 4904 197326 4916
rect 257062 4904 257068 4916
rect 257120 4904 257126 4956
rect 274450 4904 274456 4956
rect 274508 4944 274514 4956
rect 537202 4944 537208 4956
rect 274508 4916 537208 4944
rect 274508 4904 274514 4916
rect 537202 4904 537208 4916
rect 537260 4904 537266 4956
rect 59630 4836 59636 4888
rect 59688 4876 59694 4888
rect 104158 4876 104164 4888
rect 59688 4848 104164 4876
rect 59688 4836 59694 4848
rect 104158 4836 104164 4848
rect 104216 4836 104222 4888
rect 112806 4836 112812 4888
rect 112864 4876 112870 4888
rect 119338 4876 119344 4888
rect 112864 4848 119344 4876
rect 112864 4836 112870 4848
rect 119338 4836 119344 4848
rect 119396 4836 119402 4888
rect 125870 4836 125876 4888
rect 125928 4876 125934 4888
rect 160922 4876 160928 4888
rect 125928 4848 160928 4876
rect 125928 4836 125934 4848
rect 160922 4836 160928 4848
rect 160980 4836 160986 4888
rect 176562 4836 176568 4888
rect 176620 4876 176626 4888
rect 182542 4876 182548 4888
rect 176620 4848 182548 4876
rect 176620 4836 176626 4848
rect 182542 4836 182548 4848
rect 182600 4836 182606 4888
rect 198366 4836 198372 4888
rect 198424 4876 198430 4888
rect 264146 4876 264152 4888
rect 198424 4848 264152 4876
rect 198424 4836 198430 4848
rect 264146 4836 264152 4848
rect 264204 4836 264210 4888
rect 274266 4836 274272 4888
rect 274324 4876 274330 4888
rect 540790 4876 540796 4888
rect 274324 4848 540796 4876
rect 274324 4836 274330 4848
rect 540790 4836 540796 4848
rect 540848 4836 540854 4888
rect 37182 4768 37188 4820
rect 37240 4808 37246 4820
rect 66898 4808 66904 4820
rect 37240 4780 66904 4808
rect 37240 4768 37246 4780
rect 66898 4768 66904 4780
rect 66956 4768 66962 4820
rect 92750 4768 92756 4820
rect 92808 4808 92814 4820
rect 92808 4780 122834 4808
rect 92808 4768 92814 4780
rect 122806 4740 122834 4780
rect 177942 4768 177948 4820
rect 178000 4808 178006 4820
rect 189718 4808 189724 4820
rect 178000 4780 189724 4808
rect 178000 4768 178006 4780
rect 189718 4768 189724 4780
rect 189776 4768 189782 4820
rect 201126 4768 201132 4820
rect 201184 4808 201190 4820
rect 271230 4808 271236 4820
rect 201184 4780 271236 4808
rect 201184 4768 201190 4780
rect 271230 4768 271236 4780
rect 271288 4768 271294 4820
rect 275922 4768 275928 4820
rect 275980 4808 275986 4820
rect 544378 4808 544384 4820
rect 275980 4780 544384 4808
rect 275980 4768 275986 4780
rect 544378 4768 544384 4780
rect 544436 4768 544442 4820
rect 144178 4740 144184 4752
rect 122806 4712 144184 4740
rect 144178 4700 144184 4712
rect 144236 4700 144242 4752
rect 116394 4224 116400 4276
rect 116452 4264 116458 4276
rect 120902 4264 120908 4276
rect 116452 4236 120908 4264
rect 116452 4224 116458 4236
rect 120902 4224 120908 4236
rect 120960 4224 120966 4276
rect 7650 4156 7656 4208
rect 7708 4196 7714 4208
rect 11698 4196 11704 4208
rect 7708 4168 11704 4196
rect 7708 4156 7714 4168
rect 11698 4156 11704 4168
rect 11756 4156 11762 4208
rect 119890 4156 119896 4208
rect 119948 4196 119954 4208
rect 120718 4196 120724 4208
rect 119948 4168 120724 4196
rect 119948 4156 119954 4168
rect 120718 4156 120724 4168
rect 120776 4156 120782 4208
rect 164878 4156 164884 4208
rect 164936 4196 164942 4208
rect 170398 4196 170404 4208
rect 164936 4168 170404 4196
rect 164936 4156 164942 4168
rect 170398 4156 170404 4168
rect 170456 4156 170462 4208
rect 171962 4156 171968 4208
rect 172020 4196 172026 4208
rect 173158 4196 173164 4208
rect 172020 4168 173164 4196
rect 172020 4156 172026 4168
rect 173158 4156 173164 4168
rect 173216 4156 173222 4208
rect 39574 4088 39580 4140
rect 39632 4128 39638 4140
rect 130378 4128 130384 4140
rect 39632 4100 130384 4128
rect 39632 4088 39638 4100
rect 130378 4088 130384 4100
rect 130436 4088 130442 4140
rect 344554 4088 344560 4140
rect 344612 4128 344618 4140
rect 345658 4128 345664 4140
rect 344612 4100 345664 4128
rect 344612 4088 344618 4100
rect 345658 4088 345664 4100
rect 345716 4088 345722 4140
rect 468662 4088 468668 4140
rect 468720 4128 468726 4140
rect 507946 4128 507952 4140
rect 468720 4100 507952 4128
rect 468720 4088 468726 4100
rect 507946 4088 507952 4100
rect 508004 4088 508010 4140
rect 525058 4088 525064 4140
rect 525116 4128 525122 4140
rect 529014 4128 529020 4140
rect 525116 4100 529020 4128
rect 525116 4088 525122 4100
rect 529014 4088 529020 4100
rect 529072 4088 529078 4140
rect 530762 4088 530768 4140
rect 530820 4128 530826 4140
rect 550266 4128 550272 4140
rect 530820 4100 550272 4128
rect 530820 4088 530826 4100
rect 550266 4088 550272 4100
rect 550324 4088 550330 4140
rect 35986 4020 35992 4072
rect 36044 4060 36050 4072
rect 128998 4060 129004 4072
rect 36044 4032 129004 4060
rect 36044 4020 36050 4032
rect 128998 4020 129004 4032
rect 129056 4020 129062 4072
rect 465166 4020 465172 4072
rect 465224 4060 465230 4072
rect 506750 4060 506756 4072
rect 465224 4032 506756 4060
rect 465224 4020 465230 4032
rect 506750 4020 506756 4032
rect 506808 4020 506814 4072
rect 531958 4020 531964 4072
rect 532016 4060 532022 4072
rect 553762 4060 553768 4072
rect 532016 4032 553768 4060
rect 532016 4020 532022 4032
rect 553762 4020 553768 4032
rect 553820 4020 553826 4072
rect 32398 3952 32404 4004
rect 32456 3992 32462 4004
rect 127618 3992 127624 4004
rect 32456 3964 127624 3992
rect 32456 3952 32462 3964
rect 127618 3952 127624 3964
rect 127676 3952 127682 4004
rect 372890 3952 372896 4004
rect 372948 3992 372954 4004
rect 376110 3992 376116 4004
rect 372948 3964 376116 3992
rect 372948 3952 372954 3964
rect 376110 3952 376116 3964
rect 376168 3952 376174 4004
rect 458082 3952 458088 4004
rect 458140 3992 458146 4004
rect 505186 3992 505192 4004
rect 458140 3964 505192 3992
rect 458140 3952 458146 3964
rect 505186 3952 505192 3964
rect 505244 3952 505250 4004
rect 533522 3952 533528 4004
rect 533580 3992 533586 4004
rect 557350 3992 557356 4004
rect 533580 3964 557356 3992
rect 533580 3952 533586 3964
rect 557350 3952 557356 3964
rect 557408 3952 557414 4004
rect 28902 3884 28908 3936
rect 28960 3924 28966 3936
rect 127802 3924 127808 3936
rect 28960 3896 127808 3924
rect 28960 3884 28966 3896
rect 127802 3884 127808 3896
rect 127860 3884 127866 3936
rect 143534 3884 143540 3936
rect 143592 3924 143598 3936
rect 144730 3924 144736 3936
rect 143592 3896 144736 3924
rect 143592 3884 143598 3896
rect 144730 3884 144736 3896
rect 144788 3884 144794 3936
rect 454494 3884 454500 3936
rect 454552 3924 454558 3936
rect 503714 3924 503720 3936
rect 454552 3896 503720 3924
rect 454552 3884 454558 3896
rect 503714 3884 503720 3896
rect 503772 3884 503778 3936
rect 533338 3884 533344 3936
rect 533396 3924 533402 3936
rect 560846 3924 560852 3936
rect 533396 3896 560852 3924
rect 533396 3884 533402 3896
rect 560846 3884 560852 3896
rect 560904 3884 560910 3936
rect 25314 3816 25320 3868
rect 25372 3856 25378 3868
rect 157978 3856 157984 3868
rect 25372 3828 157984 3856
rect 25372 3816 25378 3828
rect 157978 3816 157984 3828
rect 158036 3816 158042 3868
rect 450906 3816 450912 3868
rect 450964 3856 450970 3868
rect 502426 3856 502432 3868
rect 450964 3828 502432 3856
rect 450964 3816 450970 3828
rect 502426 3816 502432 3828
rect 502484 3816 502490 3868
rect 534718 3816 534724 3868
rect 534776 3856 534782 3868
rect 564434 3856 564440 3868
rect 534776 3828 564440 3856
rect 534776 3816 534782 3828
rect 564434 3816 564440 3828
rect 564492 3816 564498 3868
rect 20622 3748 20628 3800
rect 20680 3788 20686 3800
rect 156598 3788 156604 3800
rect 20680 3760 156604 3788
rect 20680 3748 20686 3760
rect 156598 3748 156604 3760
rect 156656 3748 156662 3800
rect 383562 3748 383568 3800
rect 383620 3788 383626 3800
rect 385770 3788 385776 3800
rect 383620 3760 385776 3788
rect 383620 3748 383626 3760
rect 385770 3748 385776 3760
rect 385828 3748 385834 3800
rect 401318 3748 401324 3800
rect 401376 3788 401382 3800
rect 403618 3788 403624 3800
rect 401376 3760 403624 3788
rect 401376 3748 401382 3760
rect 403618 3748 403624 3760
rect 403676 3748 403682 3800
rect 408402 3748 408408 3800
rect 408460 3788 408466 3800
rect 418798 3788 418804 3800
rect 408460 3760 418804 3788
rect 408460 3748 408466 3760
rect 418798 3748 418804 3760
rect 418856 3748 418862 3800
rect 447410 3748 447416 3800
rect 447468 3788 447474 3800
rect 502610 3788 502616 3800
rect 447468 3760 502616 3788
rect 447468 3748 447474 3760
rect 502610 3748 502616 3760
rect 502668 3748 502674 3800
rect 518342 3748 518348 3800
rect 518400 3788 518406 3800
rect 521654 3788 521660 3800
rect 518400 3760 521660 3788
rect 518400 3748 518406 3760
rect 521654 3748 521660 3760
rect 521712 3748 521718 3800
rect 536282 3748 536288 3800
rect 536340 3788 536346 3800
rect 568022 3788 568028 3800
rect 536340 3760 568028 3788
rect 536340 3748 536346 3760
rect 568022 3748 568028 3760
rect 568080 3748 568086 3800
rect 15930 3680 15936 3732
rect 15988 3720 15994 3732
rect 155218 3720 155224 3732
rect 15988 3692 155224 3720
rect 15988 3680 15994 3692
rect 155218 3680 155224 3692
rect 155276 3680 155282 3732
rect 193214 3680 193220 3732
rect 193272 3720 193278 3732
rect 194410 3720 194416 3732
rect 193272 3692 194416 3720
rect 193272 3680 193278 3692
rect 194410 3680 194416 3692
rect 194468 3680 194474 3732
rect 251174 3680 251180 3732
rect 251232 3720 251238 3732
rect 252370 3720 252376 3732
rect 251232 3692 252376 3720
rect 251232 3680 251238 3692
rect 252370 3680 252376 3692
rect 252428 3680 252434 3732
rect 267734 3680 267740 3732
rect 267792 3720 267798 3732
rect 268470 3720 268476 3732
rect 267792 3692 268476 3720
rect 267792 3680 267798 3692
rect 268470 3680 268476 3692
rect 268528 3680 268534 3732
rect 284294 3680 284300 3732
rect 284352 3720 284358 3732
rect 285030 3720 285036 3732
rect 284352 3692 285036 3720
rect 284352 3680 284358 3692
rect 285030 3680 285036 3692
rect 285088 3680 285094 3732
rect 365806 3680 365812 3732
rect 365864 3720 365870 3732
rect 371878 3720 371884 3732
rect 365864 3692 371884 3720
rect 365864 3680 365870 3692
rect 371878 3680 371884 3692
rect 371936 3680 371942 3732
rect 415486 3680 415492 3732
rect 415544 3720 415550 3732
rect 440878 3720 440884 3732
rect 415544 3692 440884 3720
rect 415544 3680 415550 3692
rect 440878 3680 440884 3692
rect 440936 3680 440942 3732
rect 443822 3680 443828 3732
rect 443880 3720 443886 3732
rect 501046 3720 501052 3732
rect 443880 3692 501052 3720
rect 443880 3680 443886 3692
rect 501046 3680 501052 3692
rect 501104 3680 501110 3732
rect 516134 3680 516140 3732
rect 516192 3720 516198 3732
rect 516318 3720 516324 3732
rect 516192 3692 516324 3720
rect 516192 3680 516198 3692
rect 516318 3680 516324 3692
rect 516376 3680 516382 3732
rect 536098 3680 536104 3732
rect 536156 3720 536162 3732
rect 571518 3720 571524 3732
rect 536156 3692 571524 3720
rect 536156 3680 536162 3692
rect 571518 3680 571524 3692
rect 571576 3680 571582 3732
rect 5258 3612 5264 3664
rect 5316 3652 5322 3664
rect 158162 3652 158168 3664
rect 5316 3624 158168 3652
rect 5316 3612 5322 3624
rect 158162 3612 158168 3624
rect 158220 3612 158226 3664
rect 160094 3612 160100 3664
rect 160152 3652 160158 3664
rect 424134 3652 424140 3664
rect 160152 3624 424140 3652
rect 160152 3612 160158 3624
rect 424134 3612 424140 3624
rect 424192 3612 424198 3664
rect 440326 3612 440332 3664
rect 440384 3652 440390 3664
rect 499850 3652 499856 3664
rect 440384 3624 499856 3652
rect 440384 3612 440390 3624
rect 499850 3612 499856 3624
rect 499908 3612 499914 3664
rect 511258 3612 511264 3664
rect 511316 3652 511322 3664
rect 518986 3652 518992 3664
rect 511316 3624 518992 3652
rect 511316 3612 511322 3624
rect 518986 3612 518992 3624
rect 519044 3612 519050 3664
rect 537478 3612 537484 3664
rect 537536 3652 537542 3664
rect 575106 3652 575112 3664
rect 537536 3624 575112 3652
rect 537536 3612 537542 3624
rect 575106 3612 575112 3624
rect 575164 3612 575170 3664
rect 11146 3544 11152 3596
rect 11204 3584 11210 3596
rect 154022 3584 154028 3596
rect 11204 3556 154028 3584
rect 11204 3544 11210 3556
rect 154022 3544 154028 3556
rect 154080 3544 154086 3596
rect 156598 3544 156604 3596
rect 156656 3584 156662 3596
rect 422386 3584 422392 3596
rect 156656 3556 422392 3584
rect 156656 3544 156662 3556
rect 422386 3544 422392 3556
rect 422444 3544 422450 3596
rect 436738 3544 436744 3596
rect 436796 3584 436802 3596
rect 499666 3584 499672 3596
rect 436796 3556 499672 3584
rect 436796 3544 436802 3556
rect 499666 3544 499672 3556
rect 499724 3544 499730 3596
rect 507670 3544 507676 3596
rect 507728 3584 507734 3596
rect 519170 3584 519176 3596
rect 507728 3556 519176 3584
rect 507728 3544 507734 3556
rect 519170 3544 519176 3556
rect 519228 3544 519234 3596
rect 526438 3544 526444 3596
rect 526496 3584 526502 3596
rect 532510 3584 532516 3596
rect 526496 3556 532516 3584
rect 526496 3544 526502 3556
rect 532510 3544 532516 3556
rect 532568 3544 532574 3596
rect 541618 3544 541624 3596
rect 541676 3584 541682 3596
rect 582190 3584 582196 3596
rect 541676 3556 582196 3584
rect 541676 3544 541682 3556
rect 582190 3544 582196 3556
rect 582248 3544 582254 3596
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 3418 3516 3424 3528
rect 624 3488 3424 3516
rect 624 3476 630 3488
rect 3418 3476 3424 3488
rect 3476 3476 3482 3528
rect 24210 3476 24216 3528
rect 24268 3516 24274 3528
rect 126238 3516 126244 3528
rect 24268 3488 126244 3516
rect 24268 3476 24274 3488
rect 126238 3476 126244 3488
rect 126296 3476 126302 3528
rect 153010 3476 153016 3528
rect 153068 3516 153074 3528
rect 153068 3488 415348 3516
rect 153068 3476 153074 3488
rect 1670 3408 1676 3460
rect 1728 3448 1734 3460
rect 10318 3448 10324 3460
rect 1728 3420 10324 3448
rect 1728 3408 1734 3420
rect 10318 3408 10324 3420
rect 10376 3408 10382 3460
rect 19426 3408 19432 3460
rect 19484 3448 19490 3460
rect 124858 3448 124864 3460
rect 19484 3420 124864 3448
rect 19484 3408 19490 3420
rect 124858 3408 124864 3420
rect 124916 3408 124922 3460
rect 149514 3408 149520 3460
rect 149572 3448 149578 3460
rect 415320 3448 415348 3488
rect 415394 3476 415400 3528
rect 415452 3516 415458 3528
rect 416682 3516 416688 3528
rect 415452 3488 416688 3516
rect 415452 3476 415458 3488
rect 416682 3476 416688 3488
rect 416740 3476 416746 3528
rect 423766 3476 423772 3528
rect 423824 3516 423830 3528
rect 424962 3516 424968 3528
rect 423824 3488 424968 3516
rect 423824 3476 423830 3488
rect 424962 3476 424968 3488
rect 425020 3476 425026 3528
rect 433242 3476 433248 3528
rect 433300 3516 433306 3528
rect 433300 3488 497228 3516
rect 433300 3476 433306 3488
rect 421282 3448 421288 3460
rect 149572 3420 412772 3448
rect 415320 3420 421288 3448
rect 149572 3408 149578 3420
rect 43070 3340 43076 3392
rect 43128 3380 43134 3392
rect 131942 3380 131948 3392
rect 43128 3352 131948 3380
rect 43128 3340 43134 3352
rect 131942 3340 131948 3352
rect 132000 3340 132006 3392
rect 177850 3340 177856 3392
rect 177908 3380 177914 3392
rect 178678 3380 178684 3392
rect 177908 3352 178684 3380
rect 177908 3340 177914 3352
rect 178678 3340 178684 3352
rect 178736 3340 178742 3392
rect 184934 3340 184940 3392
rect 184992 3380 184998 3392
rect 186958 3380 186964 3392
rect 184992 3352 186964 3380
rect 184992 3340 184998 3352
rect 186958 3340 186964 3352
rect 187016 3340 187022 3392
rect 324406 3340 324412 3392
rect 324464 3380 324470 3392
rect 325602 3380 325608 3392
rect 324464 3352 325608 3380
rect 324464 3340 324470 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 332594 3340 332600 3392
rect 332652 3380 332658 3392
rect 333882 3380 333888 3392
rect 332652 3352 333888 3380
rect 332652 3340 332658 3352
rect 333882 3340 333888 3352
rect 333940 3340 333946 3392
rect 337470 3340 337476 3392
rect 337528 3380 337534 3392
rect 340138 3380 340144 3392
rect 337528 3352 340144 3380
rect 337528 3340 337534 3352
rect 340138 3340 340144 3352
rect 340196 3340 340202 3392
rect 340874 3340 340880 3392
rect 340932 3380 340938 3392
rect 342162 3380 342168 3392
rect 340932 3352 342168 3380
rect 340932 3340 340938 3352
rect 342162 3340 342168 3352
rect 342220 3340 342226 3392
rect 349154 3340 349160 3392
rect 349212 3380 349218 3392
rect 350442 3380 350448 3392
rect 349212 3352 350448 3380
rect 349212 3340 349218 3352
rect 350442 3340 350448 3352
rect 350500 3340 350506 3392
rect 351638 3340 351644 3392
rect 351696 3380 351702 3392
rect 353938 3380 353944 3392
rect 351696 3352 353944 3380
rect 351696 3340 351702 3352
rect 353938 3340 353944 3352
rect 353996 3340 354002 3392
rect 355226 3340 355232 3392
rect 355284 3380 355290 3392
rect 356790 3380 356796 3392
rect 355284 3352 356796 3380
rect 355284 3340 355290 3352
rect 356790 3340 356796 3352
rect 356848 3340 356854 3392
rect 357434 3340 357440 3392
rect 357492 3380 357498 3392
rect 358722 3380 358728 3392
rect 357492 3352 358728 3380
rect 357492 3340 357498 3352
rect 358722 3340 358728 3352
rect 358780 3340 358786 3392
rect 362310 3340 362316 3392
rect 362368 3380 362374 3392
rect 363690 3380 363696 3392
rect 362368 3352 363696 3380
rect 362368 3340 362374 3352
rect 363690 3340 363696 3352
rect 363748 3340 363754 3392
rect 365714 3340 365720 3392
rect 365772 3380 365778 3392
rect 367002 3380 367008 3392
rect 365772 3352 367008 3380
rect 365772 3340 365778 3352
rect 367002 3340 367008 3352
rect 367060 3340 367066 3392
rect 369394 3340 369400 3392
rect 369452 3380 369458 3392
rect 370590 3380 370596 3392
rect 369452 3352 370596 3380
rect 369452 3340 369458 3352
rect 370590 3340 370596 3352
rect 370648 3340 370654 3392
rect 376478 3340 376484 3392
rect 376536 3380 376542 3392
rect 378778 3380 378784 3392
rect 376536 3352 378784 3380
rect 376536 3340 376542 3352
rect 378778 3340 378784 3352
rect 378836 3340 378842 3392
rect 379974 3340 379980 3392
rect 380032 3380 380038 3392
rect 382918 3380 382924 3392
rect 380032 3352 382924 3380
rect 380032 3340 380038 3352
rect 382918 3340 382924 3352
rect 382976 3340 382982 3392
rect 412744 3380 412772 3420
rect 421282 3408 421288 3420
rect 421340 3408 421346 3460
rect 426158 3408 426164 3460
rect 426216 3448 426222 3460
rect 497090 3448 497096 3460
rect 426216 3420 497096 3448
rect 426216 3408 426222 3420
rect 497090 3408 497096 3420
rect 497148 3408 497154 3460
rect 497200 3448 497228 3488
rect 498194 3476 498200 3528
rect 498252 3516 498258 3528
rect 499022 3516 499028 3528
rect 498252 3488 499028 3516
rect 498252 3476 498258 3488
rect 499022 3476 499028 3488
rect 499080 3476 499086 3528
rect 504174 3476 504180 3528
rect 504232 3516 504238 3528
rect 517514 3516 517520 3528
rect 504232 3488 517520 3516
rect 504232 3476 504238 3488
rect 517514 3476 517520 3488
rect 517572 3476 517578 3528
rect 521838 3476 521844 3528
rect 521896 3516 521902 3528
rect 523126 3516 523132 3528
rect 521896 3488 523132 3516
rect 521896 3476 521902 3488
rect 523126 3476 523132 3488
rect 523184 3476 523190 3528
rect 526714 3476 526720 3528
rect 526772 3516 526778 3528
rect 536098 3516 536104 3528
rect 526772 3488 536104 3516
rect 526772 3476 526778 3488
rect 536098 3476 536104 3488
rect 536156 3476 536162 3528
rect 538858 3476 538864 3528
rect 538916 3516 538922 3528
rect 578602 3516 578608 3528
rect 538916 3488 578608 3516
rect 538916 3476 538922 3488
rect 578602 3476 578608 3488
rect 578660 3476 578666 3528
rect 498378 3448 498384 3460
rect 497200 3420 498384 3448
rect 498378 3408 498384 3420
rect 498436 3408 498442 3460
rect 500586 3408 500592 3460
rect 500644 3448 500650 3460
rect 516134 3448 516140 3460
rect 500644 3420 516140 3448
rect 500644 3408 500650 3420
rect 516134 3408 516140 3420
rect 516192 3408 516198 3460
rect 527910 3408 527916 3460
rect 527968 3448 527974 3460
rect 539594 3448 539600 3460
rect 527968 3420 539600 3448
rect 527968 3408 527974 3420
rect 539594 3408 539600 3420
rect 539652 3408 539658 3460
rect 540238 3408 540244 3460
rect 540296 3448 540302 3460
rect 580994 3448 581000 3460
rect 540296 3420 581000 3448
rect 540296 3408 540302 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 421098 3380 421104 3392
rect 412744 3352 421104 3380
rect 421098 3340 421104 3352
rect 421156 3340 421162 3392
rect 448514 3340 448520 3392
rect 448572 3380 448578 3392
rect 449802 3380 449808 3392
rect 448572 3352 449808 3380
rect 448572 3340 448578 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 472250 3340 472256 3392
rect 472308 3380 472314 3392
rect 509418 3380 509424 3392
rect 472308 3352 509424 3380
rect 472308 3340 472314 3352
rect 509418 3340 509424 3352
rect 509476 3340 509482 3392
rect 530578 3340 530584 3392
rect 530636 3380 530642 3392
rect 546678 3380 546684 3392
rect 530636 3352 546684 3380
rect 530636 3340 530642 3352
rect 546678 3340 546684 3352
rect 546736 3340 546742 3392
rect 4062 3272 4068 3324
rect 4120 3312 4126 3324
rect 4798 3312 4804 3324
rect 4120 3284 4804 3312
rect 4120 3272 4126 3284
rect 4798 3272 4804 3284
rect 4856 3272 4862 3324
rect 46658 3272 46664 3324
rect 46716 3312 46722 3324
rect 131758 3312 131764 3324
rect 46716 3284 131764 3312
rect 46716 3272 46722 3284
rect 131758 3272 131764 3284
rect 131816 3272 131822 3324
rect 319714 3272 319720 3324
rect 319772 3312 319778 3324
rect 320818 3312 320824 3324
rect 319772 3284 320824 3312
rect 319772 3272 319778 3284
rect 320818 3272 320824 3284
rect 320876 3272 320882 3324
rect 340966 3272 340972 3324
rect 341024 3312 341030 3324
rect 342898 3312 342904 3324
rect 341024 3284 342904 3312
rect 341024 3272 341030 3284
rect 342898 3272 342904 3284
rect 342956 3272 342962 3324
rect 475746 3272 475752 3324
rect 475804 3312 475810 3324
rect 509694 3312 509700 3324
rect 475804 3284 509700 3312
rect 475804 3272 475810 3284
rect 509694 3272 509700 3284
rect 509752 3272 509758 3324
rect 529198 3272 529204 3324
rect 529256 3312 529262 3324
rect 543182 3312 543188 3324
rect 529256 3284 543188 3312
rect 529256 3272 529262 3284
rect 543182 3272 543188 3284
rect 543240 3272 543246 3324
rect 77294 3204 77300 3256
rect 77352 3244 77358 3256
rect 78214 3244 78220 3256
rect 77352 3216 78220 3244
rect 77352 3204 77358 3216
rect 78214 3204 78220 3216
rect 78272 3204 78278 3256
rect 102134 3204 102140 3256
rect 102192 3244 102198 3256
rect 103330 3244 103336 3256
rect 102192 3216 103336 3244
rect 102192 3204 102198 3216
rect 103330 3204 103336 3216
rect 103388 3204 103394 3256
rect 121086 3204 121092 3256
rect 121144 3244 121150 3256
rect 152458 3244 152464 3256
rect 121144 3216 152464 3244
rect 121144 3204 121150 3216
rect 152458 3204 152464 3216
rect 152516 3204 152522 3256
rect 305546 3204 305552 3256
rect 305604 3244 305610 3256
rect 307018 3244 307024 3256
rect 305604 3216 307024 3244
rect 305604 3204 305610 3216
rect 307018 3204 307024 3216
rect 307076 3204 307082 3256
rect 479334 3204 479340 3256
rect 479392 3244 479398 3256
rect 510614 3244 510620 3256
rect 479392 3216 510620 3244
rect 479392 3204 479398 3216
rect 510614 3204 510620 3216
rect 510672 3204 510678 3256
rect 516502 3244 516508 3256
rect 512840 3216 516508 3244
rect 13538 3136 13544 3188
rect 13596 3176 13602 3188
rect 15838 3176 15844 3188
rect 13596 3148 15844 3176
rect 13596 3136 13602 3148
rect 15838 3136 15844 3148
rect 15896 3136 15902 3188
rect 124674 3136 124680 3188
rect 124732 3176 124738 3188
rect 153838 3176 153844 3188
rect 124732 3148 153844 3176
rect 124732 3136 124738 3148
rect 153838 3136 153844 3148
rect 153896 3136 153902 3188
rect 390554 3136 390560 3188
rect 390612 3176 390618 3188
rect 391842 3176 391848 3188
rect 390612 3148 391848 3176
rect 390612 3136 390618 3148
rect 391842 3136 391848 3148
rect 391900 3136 391906 3188
rect 397730 3136 397736 3188
rect 397788 3176 397794 3188
rect 400950 3176 400956 3188
rect 397788 3148 400956 3176
rect 397788 3136 397794 3148
rect 400950 3136 400956 3148
rect 401008 3136 401014 3188
rect 489914 3136 489920 3188
rect 489972 3176 489978 3188
rect 490742 3176 490748 3188
rect 489972 3148 490748 3176
rect 489972 3136 489978 3148
rect 490742 3136 490748 3148
rect 490800 3136 490806 3188
rect 497090 3136 497096 3188
rect 497148 3176 497154 3188
rect 512840 3176 512868 3216
rect 516502 3204 516508 3216
rect 516560 3204 516566 3256
rect 497148 3148 512868 3176
rect 497148 3136 497154 3148
rect 514754 3136 514760 3188
rect 514812 3176 514818 3188
rect 520366 3176 520372 3188
rect 514812 3148 520372 3176
rect 514812 3136 514818 3148
rect 520366 3136 520372 3148
rect 520424 3136 520430 3188
rect 525150 3136 525156 3188
rect 525208 3176 525214 3188
rect 527818 3176 527824 3188
rect 525208 3148 527824 3176
rect 525208 3136 525214 3148
rect 527818 3136 527824 3148
rect 527876 3136 527882 3188
rect 309042 3000 309048 3052
rect 309100 3040 309106 3052
rect 311158 3040 311164 3052
rect 309100 3012 311164 3040
rect 309100 3000 309106 3012
rect 311158 3000 311164 3012
rect 311216 3000 311222 3052
rect 522298 3000 522304 3052
rect 522356 3040 522362 3052
rect 524230 3040 524236 3052
rect 522356 3012 524236 3040
rect 522356 3000 522362 3012
rect 524230 3000 524236 3012
rect 524288 3000 524294 3052
rect 8754 2932 8760 2984
rect 8812 2972 8818 2984
rect 14458 2972 14464 2984
rect 8812 2944 14464 2972
rect 8812 2932 8818 2944
rect 14458 2932 14464 2944
rect 14516 2932 14522 2984
rect 523678 2932 523684 2984
rect 523736 2972 523742 2984
rect 525426 2972 525432 2984
rect 523736 2944 525432 2972
rect 523736 2932 523742 2944
rect 525426 2932 525432 2944
rect 525484 2932 525490 2984
rect 326798 2864 326804 2916
rect 326856 2904 326862 2916
rect 329098 2904 329104 2916
rect 326856 2876 329104 2904
rect 326856 2864 326862 2876
rect 329098 2864 329104 2876
rect 329156 2864 329162 2916
rect 390646 2864 390652 2916
rect 390704 2904 390710 2916
rect 392578 2904 392584 2916
rect 390704 2876 392584 2904
rect 390704 2864 390710 2876
rect 392578 2864 392584 2876
rect 392636 2864 392642 2916
<< via1 >>
rect 10324 558900 10376 558952
rect 57428 558900 57480 558952
rect 381912 59780 381964 59832
rect 383292 59780 383344 59832
rect 64788 59712 64840 59764
rect 65892 59712 65944 59764
rect 94504 59712 94556 59764
rect 97080 59712 97132 59764
rect 98828 59712 98880 59764
rect 100944 59712 100996 59764
rect 105544 59712 105596 59764
rect 107752 59712 107804 59764
rect 108488 59712 108540 59764
rect 110696 59712 110748 59764
rect 113824 59712 113876 59764
rect 115572 59712 115624 59764
rect 124864 59712 124916 59764
rect 127256 59712 127308 59764
rect 129004 59712 129056 59764
rect 131120 59712 131172 59764
rect 131764 59712 131816 59764
rect 134064 59712 134116 59764
rect 135168 59712 135220 59764
rect 137008 59712 137060 59764
rect 141424 59712 141476 59764
rect 143816 59712 143868 59764
rect 145564 59712 145616 59764
rect 147680 59712 147732 59764
rect 148324 59712 148376 59764
rect 150624 59712 150676 59764
rect 155224 59712 155276 59764
rect 157432 59712 157484 59764
rect 160744 59712 160796 59764
rect 163320 59712 163372 59764
rect 179328 59712 179380 59764
rect 180800 59712 180852 59764
rect 184756 59712 184808 59764
rect 186596 59712 186648 59764
rect 193220 59712 193272 59764
rect 193772 59712 193824 59764
rect 202788 59712 202840 59764
rect 204168 59712 204220 59764
rect 208032 59712 208084 59764
rect 209688 59712 209740 59764
rect 210976 59712 211028 59764
rect 212908 59712 212960 59764
rect 220544 59712 220596 59764
rect 222660 59712 222712 59764
rect 227536 59712 227588 59764
rect 229468 59712 229520 59764
rect 230112 59712 230164 59764
rect 232412 59712 232464 59764
rect 238668 59712 238720 59764
rect 240140 59712 240192 59764
rect 246672 59712 246724 59764
rect 248972 59712 249024 59764
rect 250996 59712 251048 59764
rect 252836 59712 252888 59764
rect 271788 59712 271840 59764
rect 273260 59712 273312 59764
rect 278688 59712 278740 59764
rect 280068 59712 280120 59764
rect 287704 59712 287756 59764
rect 289820 59712 289872 59764
rect 290464 59712 290516 59764
rect 292764 59712 292816 59764
rect 315764 59712 315816 59764
rect 317604 59712 317656 59764
rect 322572 59712 322624 59764
rect 324688 59712 324740 59764
rect 334348 59712 334400 59764
rect 335268 59712 335320 59764
rect 339132 59712 339184 59764
rect 340972 59712 341024 59764
rect 355600 59712 355652 59764
rect 358268 59712 358320 59764
rect 365352 59712 365404 59764
rect 367744 59712 367796 59764
rect 369308 59712 369360 59764
rect 371976 59712 372028 59764
rect 385960 59712 386012 59764
rect 388628 59712 388680 59764
rect 388720 59712 388772 59764
rect 391388 59712 391440 59764
rect 391664 59712 391716 59764
rect 394148 59712 394200 59764
rect 395712 59712 395764 59764
rect 398104 59712 398156 59764
rect 398472 59712 398524 59764
rect 401048 59712 401100 59764
rect 402428 59712 402480 59764
rect 405188 59712 405240 59764
rect 405280 59712 405332 59764
rect 407948 59712 408000 59764
rect 410156 59712 410208 59764
rect 411904 59712 411956 59764
rect 413100 59712 413152 59764
rect 414664 59712 414716 59764
rect 438032 59712 438084 59764
rect 438860 59712 438912 59764
rect 456616 59712 456668 59764
rect 457076 59712 457128 59764
rect 461584 59712 461636 59764
rect 462412 59712 462464 59764
rect 470600 59712 470652 59764
rect 471980 59712 472032 59764
rect 474372 59712 474424 59764
rect 476396 59712 476448 59764
rect 480260 59712 480312 59764
rect 481640 59712 481692 59764
rect 495900 59712 495952 59764
rect 496912 59712 496964 59764
rect 500684 59712 500736 59764
rect 502616 59712 502668 59764
rect 503628 59712 503680 59764
rect 505192 59712 505244 59764
rect 517244 59712 517296 59764
rect 519176 59712 519228 59764
rect 522120 59712 522172 59764
rect 523684 59712 523736 59764
rect 524052 59712 524104 59764
rect 526444 59712 526496 59764
rect 526996 59712 527048 59764
rect 529204 59712 529256 59764
rect 530860 59712 530912 59764
rect 533528 59712 533580 59764
rect 533804 59712 533856 59764
rect 536288 59712 536340 59764
rect 123484 59576 123536 59628
rect 125324 59576 125376 59628
rect 159364 59576 159416 59628
rect 161296 59576 161348 59628
rect 198372 59576 198424 59628
rect 200028 59576 200080 59628
rect 242808 59576 242860 59628
rect 244096 59576 244148 59628
rect 269028 59576 269080 59628
rect 270316 59576 270368 59628
rect 275928 59576 275980 59628
rect 277124 59576 277176 59628
rect 284944 59576 284996 59628
rect 286876 59576 286928 59628
rect 295248 59576 295300 59628
rect 296628 59576 296680 59628
rect 324504 59576 324556 59628
rect 325700 59576 325752 59628
rect 374092 59576 374144 59628
rect 376024 59576 376076 59628
rect 419816 59576 419868 59628
rect 421104 59576 421156 59628
rect 456892 59576 456944 59628
rect 458272 59576 458324 59628
rect 492864 59576 492916 59628
rect 494152 59576 494204 59628
rect 61936 59440 61988 59492
rect 63960 59440 64012 59492
rect 113272 59440 113324 59492
rect 114652 59440 114704 59492
rect 152464 59440 152516 59492
rect 154488 59440 154540 59492
rect 165068 59440 165120 59492
rect 167184 59440 167236 59492
rect 235908 59440 235960 59492
rect 237380 59440 237432 59492
rect 244188 59440 244240 59492
rect 246028 59440 246080 59492
rect 352748 59440 352800 59492
rect 354680 59440 354732 59492
rect 497740 59440 497792 59492
rect 499672 59440 499724 59492
rect 507492 59440 507544 59492
rect 509424 59440 509476 59492
rect 11704 59372 11756 59424
rect 59360 59372 59412 59424
rect 103520 59372 103572 59424
rect 104900 59372 104952 59424
rect 542268 59372 542320 59424
rect 582380 59372 582432 59424
rect 85028 59304 85080 59356
rect 89720 59304 89772 59356
rect 168380 59304 168432 59356
rect 173992 59304 174044 59356
rect 346400 59304 346452 59356
rect 347780 59304 347832 59356
rect 447140 58896 447192 58948
rect 448520 58896 448572 58948
rect 267740 58828 267792 58880
rect 326160 58828 326212 58880
rect 371148 58828 371200 58880
rect 427820 58828 427872 58880
rect 91008 58760 91060 58812
rect 92296 58760 92348 58812
rect 190460 58760 190512 58812
rect 305000 58760 305052 58812
rect 319628 58760 319680 58812
rect 321744 58760 321796 58812
rect 335360 58760 335412 58812
rect 345388 58760 345440 58812
rect 392584 58760 392636 58812
rect 483480 58760 483532 58812
rect 237380 58692 237432 58744
rect 441988 58692 442040 58744
rect 3424 58624 3476 58676
rect 57980 58624 58032 58676
rect 104900 58624 104952 58676
rect 118608 58624 118660 58676
rect 150440 58624 150492 58676
rect 168288 58624 168340 58676
rect 193036 58624 193088 58676
rect 231860 58624 231912 58676
rect 264796 58624 264848 58676
rect 494060 58624 494112 58676
rect 91744 58488 91796 58540
rect 94136 58488 94188 58540
rect 253572 58488 253624 58540
rect 254308 58488 254360 58540
rect 320456 58488 320508 58540
rect 321928 58488 321980 58540
rect 448152 58352 448204 58404
rect 450176 58352 450228 58404
rect 446404 58080 446456 58132
rect 447416 58080 447468 58132
rect 75920 57944 75972 57996
rect 78496 57944 78548 57996
rect 354680 57944 354732 57996
rect 360200 57944 360252 57996
rect 215300 57400 215352 57452
rect 311992 57400 312044 57452
rect 161480 57332 161532 57384
rect 295248 57332 295300 57384
rect 321560 57332 321612 57384
rect 340880 57332 340932 57384
rect 383844 57332 383896 57384
rect 470600 57332 470652 57384
rect 194600 57264 194652 57316
rect 430580 57264 430632 57316
rect 53840 57196 53892 57248
rect 71780 57196 71832 57248
rect 87972 57196 88024 57248
rect 100760 57196 100812 57248
rect 267648 57196 267700 57248
rect 507860 57196 507912 57248
rect 276020 56108 276072 56160
rect 328552 56108 328604 56160
rect 206744 56040 206796 56092
rect 281540 56040 281592 56092
rect 204260 55972 204312 56024
rect 308956 55972 309008 56024
rect 316040 55972 316092 56024
rect 463608 55972 463660 56024
rect 16580 55904 16632 55956
rect 61936 55904 61988 55956
rect 186964 55904 187016 55956
rect 427636 55904 427688 55956
rect 56600 55836 56652 55888
rect 135168 55836 135220 55888
rect 277308 55836 277360 55888
rect 547880 55836 547932 55888
rect 208400 54680 208452 54732
rect 311900 54680 311952 54732
rect 418804 54680 418856 54732
rect 488632 54680 488684 54732
rect 244188 54612 244240 54664
rect 430580 54612 430632 54664
rect 26240 54544 26292 54596
rect 64788 54544 64840 54596
rect 251180 54544 251232 54596
rect 448520 54544 448572 54596
rect 60740 54476 60792 54528
rect 135904 54476 135956 54528
rect 279884 54476 279936 54528
rect 557540 54476 557592 54528
rect 193220 53252 193272 53304
rect 307944 53252 307996 53304
rect 257988 53184 258040 53236
rect 476120 53184 476172 53236
rect 142160 53116 142212 53168
rect 418160 53116 418212 53168
rect 29000 53048 29052 53100
rect 65984 53048 66036 53100
rect 280068 53048 280120 53100
rect 561680 53048 561732 53100
rect 260840 51960 260892 52012
rect 327080 51960 327132 52012
rect 204168 51892 204220 51944
rect 284300 51892 284352 51944
rect 201500 51824 201552 51876
rect 310520 51824 310572 51876
rect 311164 51824 311216 51876
rect 463700 51824 463752 51876
rect 187700 51756 187752 51808
rect 430672 51756 430724 51808
rect 4804 51688 4856 51740
rect 92204 51688 92256 51740
rect 284116 51688 284168 51740
rect 572720 51688 572772 51740
rect 218060 50532 218112 50584
rect 314844 50532 314896 50584
rect 227536 50464 227588 50516
rect 369860 50464 369912 50516
rect 383936 50464 383988 50516
rect 466460 50464 466512 50516
rect 311900 50396 311952 50448
rect 465080 50396 465132 50448
rect 14464 50328 14516 50380
rect 91744 50328 91796 50380
rect 110420 50328 110472 50380
rect 149704 50328 149756 50380
rect 283932 50328 283984 50380
rect 575480 50328 575532 50380
rect 208216 49172 208268 49224
rect 295340 49172 295392 49224
rect 371884 49172 371936 49224
rect 480352 49172 480404 49224
rect 224776 49104 224828 49156
rect 356060 49104 356112 49156
rect 402244 49104 402296 49156
rect 534080 49104 534132 49156
rect 252468 49036 252520 49088
rect 458180 49036 458232 49088
rect 52460 48968 52512 49020
rect 102784 48968 102836 49020
rect 135260 48968 135312 49020
rect 416872 48968 416924 49020
rect 208032 47744 208084 47796
rect 299480 47744 299532 47796
rect 226248 47676 226300 47728
rect 362960 47676 363012 47728
rect 405188 47676 405240 47728
rect 540980 47676 541032 47728
rect 244280 47608 244332 47660
rect 447140 47608 447192 47660
rect 17960 47540 18012 47592
rect 95148 47540 95200 47592
rect 102140 47540 102192 47592
rect 148508 47540 148560 47592
rect 253756 47540 253808 47592
rect 465080 47540 465132 47592
rect 222108 46384 222160 46436
rect 349252 46384 349304 46436
rect 370596 46384 370648 46436
rect 480444 46384 480496 46436
rect 143540 46316 143592 46368
rect 290648 46316 290700 46368
rect 401048 46316 401100 46368
rect 525156 46316 525208 46368
rect 242808 46248 242860 46300
rect 423680 46248 423732 46300
rect 44180 46180 44232 46232
rect 101588 46180 101640 46232
rect 241520 46180 241572 46232
rect 445760 46180 445812 46232
rect 220544 45024 220596 45076
rect 345020 45024 345072 45076
rect 399484 45024 399536 45076
rect 522304 45024 522356 45076
rect 147680 44956 147732 45008
rect 290464 44956 290516 45008
rect 342904 44956 342956 45008
rect 473452 44956 473504 45008
rect 240048 44888 240100 44940
rect 412640 44888 412692 44940
rect 80060 44820 80112 44872
rect 111248 44820 111300 44872
rect 198740 44820 198792 44872
rect 433524 44820 433576 44872
rect 282920 43596 282972 43648
rect 332600 43596 332652 43648
rect 380164 43596 380216 43648
rect 452660 43596 452712 43648
rect 213736 43528 213788 43580
rect 320180 43528 320232 43580
rect 391388 43528 391440 43580
rect 491300 43528 491352 43580
rect 230296 43460 230348 43512
rect 376760 43460 376812 43512
rect 382924 43460 382976 43512
rect 483112 43460 483164 43512
rect 180800 43392 180852 43444
rect 429200 43392 429252 43444
rect 220728 42236 220780 42288
rect 340880 42236 340932 42288
rect 398288 42236 398340 42288
rect 520280 42236 520332 42288
rect 340144 42168 340196 42220
rect 471980 42168 472032 42220
rect 237196 42100 237248 42152
rect 405740 42100 405792 42152
rect 173900 42032 173952 42084
rect 426532 42032 426584 42084
rect 219348 40876 219400 40928
rect 338120 40876 338172 40928
rect 398104 40876 398156 40928
rect 516140 40876 516192 40928
rect 329840 40808 329892 40860
rect 469312 40808 469364 40860
rect 237012 40740 237064 40792
rect 401600 40740 401652 40792
rect 169760 40672 169812 40724
rect 426716 40672 426768 40724
rect 217876 39516 217928 39568
rect 333980 39516 334032 39568
rect 392676 39516 392728 39568
rect 498200 39516 498252 39568
rect 329104 39448 329156 39500
rect 469496 39448 469548 39500
rect 235908 39380 235960 39432
rect 398840 39380 398892 39432
rect 167000 39312 167052 39364
rect 425060 39312 425112 39364
rect 314660 38088 314712 38140
rect 341156 38088 341208 38140
rect 387064 38088 387116 38140
rect 477500 38088 477552 38140
rect 217692 38020 217744 38072
rect 331220 38020 331272 38072
rect 391204 38020 391256 38072
rect 495440 38020 495492 38072
rect 234436 37952 234488 38004
rect 394700 37952 394752 38004
rect 178684 37884 178736 37936
rect 427912 37884 427964 37936
rect 216588 36660 216640 36712
rect 327080 36660 327132 36712
rect 354036 36660 354088 36712
rect 476396 36660 476448 36712
rect 233148 36592 233200 36644
rect 387800 36592 387852 36644
rect 405004 36592 405056 36644
rect 545120 36592 545172 36644
rect 88340 36524 88392 36576
rect 144368 36524 144420 36576
rect 256608 36524 256660 36576
rect 473360 36524 473412 36576
rect 215208 35300 215260 35352
rect 324320 35300 324372 35352
rect 345664 35300 345716 35352
rect 473636 35300 473688 35352
rect 230112 35232 230164 35284
rect 380900 35232 380952 35284
rect 403624 35232 403676 35284
rect 538220 35232 538272 35284
rect 85580 35164 85632 35216
rect 142804 35164 142856 35216
rect 255228 35164 255280 35216
rect 469220 35164 469272 35216
rect 197360 33940 197412 33992
rect 309140 33940 309192 33992
rect 383016 33940 383068 33992
rect 463700 33940 463752 33992
rect 223488 33872 223540 33924
rect 351920 33872 351972 33924
rect 403624 33872 403676 33924
rect 490012 33872 490064 33924
rect 131120 33804 131172 33856
rect 415400 33804 415452 33856
rect 282828 33736 282880 33788
rect 568580 33736 568632 33788
rect 176660 32580 176712 32632
rect 303620 32580 303672 32632
rect 372160 32580 372212 32632
rect 423772 32580 423824 32632
rect 224592 32512 224644 32564
rect 358820 32512 358872 32564
rect 378876 32512 378928 32564
rect 483296 32512 483348 32564
rect 201592 32444 201644 32496
rect 434720 32444 434772 32496
rect 77300 32376 77352 32428
rect 141608 32376 141660 32428
rect 281448 32376 281500 32428
rect 564532 32376 564584 32428
rect 278780 31220 278832 31272
rect 331404 31220 331456 31272
rect 140780 31152 140832 31204
rect 289084 31152 289136 31204
rect 356796 31152 356848 31204
rect 476212 31152 476264 31204
rect 253572 31084 253624 31136
rect 462320 31084 462372 31136
rect 70400 31016 70452 31068
rect 138664 31016 138716 31068
rect 202788 31016 202840 31068
rect 277400 31016 277452 31068
rect 278688 31016 278740 31068
rect 554780 31016 554832 31068
rect 271880 29792 271932 29844
rect 329932 29792 329984 29844
rect 400956 29792 401008 29844
rect 488540 29792 488592 29844
rect 250996 29724 251048 29776
rect 455420 29724 455472 29776
rect 201316 29656 201368 29708
rect 274640 29656 274692 29708
rect 277032 29656 277084 29708
rect 550640 29656 550692 29708
rect 67640 29588 67692 29640
rect 137468 29588 137520 29640
rect 144920 29588 144972 29640
rect 419540 29588 419592 29640
rect 227352 28432 227404 28484
rect 365720 28432 365772 28484
rect 371976 28432 372028 28484
rect 420920 28432 420972 28484
rect 126980 28364 127032 28416
rect 284944 28364 284996 28416
rect 376116 28364 376168 28416
rect 481640 28364 481692 28416
rect 191840 28296 191892 28348
rect 431960 28296 432012 28348
rect 37280 28228 37332 28280
rect 98828 28228 98880 28280
rect 273168 28228 273220 28280
rect 532700 28228 532752 28280
rect 264980 27004 265032 27056
rect 327264 27004 327316 27056
rect 332600 27004 332652 27056
rect 470692 27004 470744 27056
rect 248328 26936 248380 26988
rect 444380 26936 444432 26988
rect 22100 26868 22152 26920
rect 94504 26868 94556 26920
rect 200028 26868 200080 26920
rect 267832 26868 267884 26920
rect 270316 26868 270368 26920
rect 523224 26868 523276 26920
rect 136640 25712 136692 25764
rect 287704 25712 287756 25764
rect 246856 25644 246908 25696
rect 437480 25644 437532 25696
rect 248420 25576 248472 25628
rect 447416 25576 447468 25628
rect 91100 25508 91152 25560
rect 113824 25508 113876 25560
rect 198556 25508 198608 25560
rect 259460 25508 259512 25560
rect 264888 25508 264940 25560
rect 505100 25508 505152 25560
rect 247040 24284 247092 24336
rect 322940 24284 322992 24336
rect 320824 24216 320876 24268
rect 466644 24216 466696 24268
rect 245568 24148 245620 24200
rect 433340 24148 433392 24200
rect 86960 24080 87012 24132
rect 112444 24080 112496 24132
rect 194416 24080 194468 24132
rect 249800 24080 249852 24132
rect 263324 24080 263376 24132
rect 500960 24080 501012 24132
rect 236000 22924 236052 22976
rect 320272 22924 320324 22976
rect 307024 22856 307076 22908
rect 463884 22856 463936 22908
rect 81440 22788 81492 22840
rect 141424 22788 141476 22840
rect 243912 22788 243964 22840
rect 426440 22788 426492 22840
rect 15844 22720 15896 22772
rect 93124 22720 93176 22772
rect 194232 22720 194284 22772
rect 245660 22720 245712 22772
rect 263508 22720 263560 22772
rect 498292 22720 498344 22772
rect 226340 21564 226392 21616
rect 317604 21564 317656 21616
rect 385776 21564 385828 21616
rect 484400 21564 484452 21616
rect 287060 21496 287112 21548
rect 458272 21496 458324 21548
rect 241244 21428 241296 21480
rect 419540 21428 419592 21480
rect 77392 21360 77444 21412
rect 109684 21360 109736 21412
rect 188988 21360 189040 21412
rect 227720 21360 227772 21412
rect 260564 21360 260616 21412
rect 489920 21360 489972 21412
rect 404360 20136 404412 20188
rect 490196 20136 490248 20188
rect 222200 20068 222252 20120
rect 316132 20068 316184 20120
rect 385684 20068 385736 20120
rect 473452 20068 473504 20120
rect 241428 20000 241480 20052
rect 415400 20000 415452 20052
rect 55220 19932 55272 19984
rect 104348 19932 104400 19984
rect 113180 19932 113232 19984
rect 151268 19932 151320 19984
rect 187516 19932 187568 19984
rect 224960 19932 225012 19984
rect 260748 19932 260800 19984
rect 487160 19932 487212 19984
rect 363696 18776 363748 18828
rect 478880 18776 478932 18828
rect 229100 18708 229152 18760
rect 317420 18708 317472 18760
rect 400864 18708 400916 18760
rect 531412 18708 531464 18760
rect 238668 18640 238720 18692
rect 408500 18640 408552 18692
rect 48320 18572 48372 18624
rect 101404 18572 101456 18624
rect 106280 18572 106332 18624
rect 148324 18572 148376 18624
rect 186228 18572 186280 18624
rect 218152 18572 218204 18624
rect 259368 18572 259420 18624
rect 483020 18572 483072 18624
rect 211160 17348 211212 17400
rect 313280 17348 313332 17400
rect 347780 17348 347832 17400
rect 474740 17348 474792 17400
rect 91008 17280 91060 17332
rect 121460 17280 121512 17332
rect 234252 17280 234304 17332
rect 390560 17280 390612 17332
rect 395344 17280 395396 17332
rect 509240 17280 509292 17332
rect 30380 17212 30432 17264
rect 97264 17212 97316 17264
rect 184756 17212 184808 17264
rect 213920 17212 213972 17264
rect 257712 17212 257764 17264
rect 480260 17212 480312 17264
rect 284392 16464 284444 16516
rect 456892 16464 456944 16516
rect 280712 16396 280764 16448
rect 457076 16396 457128 16448
rect 276664 16328 276716 16380
rect 455512 16328 455564 16380
rect 273260 16260 273312 16312
rect 454040 16260 454092 16312
rect 270040 16192 270092 16244
rect 453028 16192 453080 16244
rect 266544 16124 266596 16176
rect 452844 16124 452896 16176
rect 262496 16056 262548 16108
rect 451280 16056 451332 16108
rect 259552 15988 259604 16040
rect 449992 15988 450044 16040
rect 255872 15920 255924 15972
rect 450176 15920 450228 15972
rect 85304 15852 85356 15904
rect 104072 15852 104124 15904
rect 109040 15852 109092 15904
rect 117964 15852 118016 15904
rect 138848 15852 138900 15904
rect 417056 15852 417108 15904
rect 234620 14968 234672 15020
rect 443092 14968 443144 15020
rect 231032 14900 231084 14952
rect 443276 14900 443328 14952
rect 227536 14832 227588 14884
rect 441620 14832 441672 14884
rect 223580 14764 223632 14816
rect 440516 14764 440568 14816
rect 219992 14696 220044 14748
rect 440332 14696 440384 14748
rect 216864 14628 216916 14680
rect 438860 14628 438912 14680
rect 213368 14560 213420 14612
rect 437572 14560 437624 14612
rect 493048 14560 493100 14612
rect 514760 14560 514812 14612
rect 73344 14492 73396 14544
rect 108488 14492 108540 14544
rect 147128 14492 147180 14544
rect 166264 14492 166316 14544
rect 209780 14492 209832 14544
rect 436192 14492 436244 14544
rect 33600 14424 33652 14476
rect 65524 14424 65576 14476
rect 99840 14424 99892 14476
rect 146944 14424 146996 14476
rect 206192 14424 206244 14476
rect 436376 14424 436428 14476
rect 440884 14424 440936 14476
rect 492956 14424 493008 14476
rect 158904 13404 158956 13456
rect 293408 13404 293460 13456
rect 301504 13404 301556 13456
rect 462412 13404 462464 13456
rect 155132 13336 155184 13388
rect 293224 13336 293276 13388
rect 298100 13336 298152 13388
rect 460940 13336 460992 13388
rect 151820 13268 151872 13320
rect 291844 13268 291896 13320
rect 294880 13268 294932 13320
rect 459836 13268 459888 13320
rect 291384 13200 291436 13252
rect 459652 13200 459704 13252
rect 163688 13132 163740 13184
rect 423956 13132 424008 13184
rect 21824 13064 21876 13116
rect 62764 13064 62816 13116
rect 65064 13064 65116 13116
rect 75368 13064 75420 13116
rect 89444 13064 89496 13116
rect 118792 13064 118844 13116
rect 127532 13064 127584 13116
rect 414020 13064 414072 13116
rect 486424 13064 486476 13116
rect 513472 13064 513524 13116
rect 258264 12044 258316 12096
rect 325700 12044 325752 12096
rect 254216 11976 254268 12028
rect 324504 11976 324556 12028
rect 251272 11908 251324 11960
rect 324688 11908 324740 11960
rect 240140 11840 240192 11892
rect 321744 11840 321796 11892
rect 386696 11840 386748 11892
rect 485964 11840 486016 11892
rect 61568 11772 61620 11824
rect 73804 11772 73856 11824
rect 218060 11772 218112 11824
rect 219256 11772 219308 11824
rect 233424 11772 233476 11824
rect 318800 11772 318852 11824
rect 324412 11772 324464 11824
rect 343824 11772 343876 11824
rect 357440 11772 357492 11824
rect 477592 11772 477644 11824
rect 11612 11704 11664 11756
rect 61384 11704 61436 11756
rect 89628 11704 89680 11756
rect 114744 11704 114796 11756
rect 133880 11704 133932 11756
rect 286508 11704 286560 11756
rect 322940 11704 322992 11756
rect 467840 11704 467892 11756
rect 490012 11704 490064 11756
rect 513656 11704 513708 11756
rect 259460 11636 259512 11688
rect 260656 11636 260708 11688
rect 374644 10752 374696 10804
rect 432052 10752 432104 10804
rect 186872 10684 186924 10736
rect 306380 10684 306432 10736
rect 374828 10684 374880 10736
rect 435088 10684 435140 10736
rect 183744 10616 183796 10668
rect 305276 10616 305328 10668
rect 376024 10616 376076 10668
rect 439136 10616 439188 10668
rect 180248 10548 180300 10600
rect 305092 10548 305144 10600
rect 377404 10548 377456 10600
rect 442632 10548 442684 10600
rect 169576 10480 169628 10532
rect 296168 10480 296220 10532
rect 339592 10480 339644 10532
rect 347964 10480 348016 10532
rect 377588 10480 377640 10532
rect 445760 10480 445812 10532
rect 172704 10412 172756 10464
rect 302240 10412 302292 10464
rect 332692 10412 332744 10464
rect 346492 10412 346544 10464
rect 378784 10412 378836 10464
rect 448520 10412 448572 10464
rect 84108 10344 84160 10396
rect 97448 10344 97500 10396
rect 166080 10344 166132 10396
rect 295984 10344 296036 10396
rect 307944 10344 307996 10396
rect 339500 10344 339552 10396
rect 381728 10344 381780 10396
rect 456892 10344 456944 10396
rect 51080 10276 51132 10328
rect 71044 10276 71096 10328
rect 84200 10276 84252 10328
rect 111064 10276 111116 10328
rect 130292 10276 130344 10328
rect 286324 10276 286376 10328
rect 297272 10276 297324 10328
rect 336740 10276 336792 10328
rect 355324 10276 355376 10328
rect 364616 10276 364668 10328
rect 381544 10276 381596 10328
rect 459928 10276 459980 10328
rect 482376 10276 482428 10328
rect 512000 10276 512052 10328
rect 429660 9256 429712 9308
rect 496912 9256 496964 9308
rect 412272 9188 412324 9240
rect 492772 9188 492824 9240
rect 394240 9120 394292 9172
rect 487252 9120 487304 9172
rect 180708 9052 180760 9104
rect 196808 9052 196860 9104
rect 246672 9052 246724 9104
rect 441528 9052 441580 9104
rect 86868 8984 86920 9036
rect 108120 8984 108172 9036
rect 143632 8984 143684 9036
rect 165068 8984 165120 9036
rect 184572 8984 184624 9036
rect 211068 8984 211120 9036
rect 249708 8984 249760 9036
rect 448612 8984 448664 9036
rect 47860 8916 47912 8968
rect 69664 8916 69716 8968
rect 96252 8916 96304 8968
rect 145564 8916 145616 8968
rect 193128 8916 193180 8968
rect 242900 8916 242952 8968
rect 250812 8916 250864 8968
rect 452108 8916 452160 8968
rect 461584 8916 461636 8968
rect 506572 8916 506624 8968
rect 69112 8304 69164 8356
rect 75184 8304 75236 8356
rect 81348 8304 81400 8356
rect 86868 8304 86920 8356
rect 79968 8236 80020 8288
rect 83280 8236 83332 8288
rect 369124 8236 369176 8288
rect 414296 8236 414348 8288
rect 370504 8168 370556 8220
rect 417884 8168 417936 8220
rect 422576 8168 422628 8220
rect 495532 8168 495584 8220
rect 406384 8100 406436 8152
rect 549076 8100 549128 8152
rect 407948 8032 408000 8084
rect 552664 8032 552716 8084
rect 407764 7964 407816 8016
rect 556160 7964 556212 8016
rect 365168 7896 365220 7948
rect 400128 7896 400180 7948
rect 409144 7896 409196 7948
rect 559748 7896 559800 7948
rect 366364 7828 366416 7880
rect 403716 7828 403768 7880
rect 410708 7828 410760 7880
rect 563244 7828 563296 7880
rect 367744 7760 367796 7812
rect 407212 7760 407264 7812
rect 410524 7760 410576 7812
rect 566832 7760 566884 7812
rect 179328 7692 179380 7744
rect 193312 7692 193364 7744
rect 244096 7692 244148 7744
rect 321928 7692 321980 7744
rect 329196 7692 329248 7744
rect 345112 7692 345164 7744
rect 367928 7692 367980 7744
rect 410800 7692 410852 7744
rect 411904 7692 411956 7744
rect 570328 7692 570380 7744
rect 58440 7624 58492 7676
rect 72424 7624 72476 7676
rect 82544 7624 82596 7676
rect 93952 7624 94004 7676
rect 136456 7624 136508 7676
rect 163504 7624 163556 7676
rect 181996 7624 182048 7676
rect 203892 7624 203944 7676
rect 229008 7624 229060 7676
rect 374092 7624 374144 7676
rect 413284 7624 413336 7676
rect 573916 7624 573968 7676
rect 2872 7556 2924 7608
rect 58624 7556 58676 7608
rect 88248 7556 88300 7608
rect 111616 7556 111668 7608
rect 117596 7556 117648 7608
rect 151084 7556 151136 7608
rect 157800 7556 157852 7608
rect 169024 7556 169076 7608
rect 187332 7556 187384 7608
rect 221556 7556 221608 7608
rect 231768 7556 231820 7608
rect 384764 7556 384816 7608
rect 414664 7556 414716 7608
rect 577412 7556 577464 7608
rect 72608 6876 72660 6928
rect 76564 6876 76616 6928
rect 41880 6672 41932 6724
rect 100024 6672 100076 6724
rect 300768 6672 300820 6724
rect 338488 6672 338540 6724
rect 356704 6672 356756 6724
rect 368204 6672 368256 6724
rect 34796 6604 34848 6656
rect 98644 6604 98696 6656
rect 286600 6604 286652 6656
rect 334348 6604 334400 6656
rect 358268 6604 358320 6656
rect 371700 6604 371752 6656
rect 75000 6536 75052 6588
rect 140044 6536 140096 6588
rect 205548 6536 205600 6588
rect 288992 6536 289044 6588
rect 290188 6536 290240 6588
rect 334164 6536 334216 6588
rect 358084 6536 358136 6588
rect 375288 6536 375340 6588
rect 27712 6468 27764 6520
rect 95884 6468 95936 6520
rect 206928 6468 206980 6520
rect 292580 6468 292632 6520
rect 293684 6468 293736 6520
rect 335452 6468 335504 6520
rect 359556 6468 359608 6520
rect 378876 6468 378928 6520
rect 388628 6468 388680 6520
rect 481732 6468 481784 6520
rect 64328 6400 64380 6452
rect 137284 6400 137336 6452
rect 209688 6400 209740 6452
rect 303160 6400 303212 6452
rect 304356 6400 304408 6452
rect 338304 6400 338356 6452
rect 360844 6400 360896 6452
rect 382372 6400 382424 6452
rect 388444 6400 388496 6452
rect 485228 6400 485280 6452
rect 53748 6332 53800 6384
rect 134524 6332 134576 6384
rect 210792 6332 210844 6384
rect 306748 6332 306800 6384
rect 361028 6332 361080 6384
rect 385960 6332 386012 6384
rect 389824 6332 389876 6384
rect 488816 6332 488868 6384
rect 50160 6264 50212 6316
rect 133144 6264 133196 6316
rect 177764 6264 177816 6316
rect 186136 6264 186188 6316
rect 210976 6264 211028 6316
rect 310244 6264 310296 6316
rect 311440 6264 311492 6316
rect 340972 6264 341024 6316
rect 343364 6264 343416 6316
rect 349344 6264 349396 6316
rect 362224 6264 362276 6316
rect 389456 6264 389508 6316
rect 394148 6264 394200 6316
rect 502984 6264 503036 6316
rect 14740 6196 14792 6248
rect 125048 6196 125100 6248
rect 161296 6196 161348 6248
rect 170588 6196 170640 6248
rect 181812 6196 181864 6248
rect 200304 6196 200356 6248
rect 212448 6196 212500 6248
rect 313832 6196 313884 6248
rect 363604 6196 363656 6248
rect 393044 6196 393096 6248
rect 393964 6196 394016 6248
rect 506480 6196 506532 6248
rect 9956 6128 10008 6180
rect 123484 6128 123536 6180
rect 154212 6128 154264 6180
rect 167644 6128 167696 6180
rect 183468 6128 183520 6180
rect 207388 6128 207440 6180
rect 213552 6128 213604 6180
rect 317328 6128 317380 6180
rect 318524 6128 318576 6180
rect 342260 6128 342312 6180
rect 353852 6128 353904 6180
rect 357532 6128 357584 6180
rect 364984 6128 365036 6180
rect 396540 6128 396592 6180
rect 396724 6128 396776 6180
rect 513564 6128 513616 6180
rect 174912 5516 174964 5568
rect 179052 5516 179104 5568
rect 352564 5516 352616 5568
rect 354036 5516 354088 5568
rect 98644 5312 98696 5364
rect 105544 5312 105596 5364
rect 102232 5244 102284 5296
rect 116584 5244 116636 5296
rect 267372 5244 267424 5296
rect 512460 5244 512512 5296
rect 98736 5176 98788 5228
rect 115388 5176 115440 5228
rect 267556 5176 267608 5228
rect 515956 5176 516008 5228
rect 44272 5108 44324 5160
rect 68468 5108 68520 5160
rect 95148 5108 95200 5160
rect 115204 5108 115256 5160
rect 191472 5108 191524 5160
rect 235816 5108 235868 5160
rect 269028 5108 269080 5160
rect 519544 5108 519596 5160
rect 40684 5040 40736 5092
rect 68284 5040 68336 5092
rect 70308 5040 70360 5092
rect 108304 5040 108356 5092
rect 140044 5040 140096 5092
rect 164884 5040 164936 5092
rect 191656 5040 191708 5092
rect 239312 5040 239364 5092
rect 270132 5040 270184 5092
rect 526628 5040 526680 5092
rect 66720 4972 66772 5024
rect 106924 4972 106976 5024
rect 132960 4972 133012 5024
rect 162124 4972 162176 5024
rect 195888 4972 195940 5024
rect 253480 4972 253532 5024
rect 271788 4972 271840 5024
rect 530124 4972 530176 5024
rect 63224 4904 63276 4956
rect 98644 4904 98696 4956
rect 129372 4904 129424 4956
rect 160744 4904 160796 4956
rect 197268 4904 197320 4956
rect 257068 4904 257120 4956
rect 274456 4904 274508 4956
rect 537208 4904 537260 4956
rect 59636 4836 59688 4888
rect 104164 4836 104216 4888
rect 112812 4836 112864 4888
rect 119344 4836 119396 4888
rect 125876 4836 125928 4888
rect 160928 4836 160980 4888
rect 176568 4836 176620 4888
rect 182548 4836 182600 4888
rect 198372 4836 198424 4888
rect 264152 4836 264204 4888
rect 274272 4836 274324 4888
rect 540796 4836 540848 4888
rect 37188 4768 37240 4820
rect 66904 4768 66956 4820
rect 92756 4768 92808 4820
rect 177948 4768 178000 4820
rect 189724 4768 189776 4820
rect 201132 4768 201184 4820
rect 271236 4768 271288 4820
rect 275928 4768 275980 4820
rect 544384 4768 544436 4820
rect 144184 4700 144236 4752
rect 116400 4224 116452 4276
rect 120908 4224 120960 4276
rect 7656 4156 7708 4208
rect 11704 4156 11756 4208
rect 119896 4156 119948 4208
rect 120724 4156 120776 4208
rect 164884 4156 164936 4208
rect 170404 4156 170456 4208
rect 171968 4156 172020 4208
rect 173164 4156 173216 4208
rect 39580 4088 39632 4140
rect 130384 4088 130436 4140
rect 344560 4088 344612 4140
rect 345664 4088 345716 4140
rect 468668 4088 468720 4140
rect 507952 4088 508004 4140
rect 525064 4088 525116 4140
rect 529020 4088 529072 4140
rect 530768 4088 530820 4140
rect 550272 4088 550324 4140
rect 35992 4020 36044 4072
rect 129004 4020 129056 4072
rect 465172 4020 465224 4072
rect 506756 4020 506808 4072
rect 531964 4020 532016 4072
rect 553768 4020 553820 4072
rect 32404 3952 32456 4004
rect 127624 3952 127676 4004
rect 372896 3952 372948 4004
rect 376116 3952 376168 4004
rect 458088 3952 458140 4004
rect 505192 3952 505244 4004
rect 533528 3952 533580 4004
rect 557356 3952 557408 4004
rect 28908 3884 28960 3936
rect 127808 3884 127860 3936
rect 143540 3884 143592 3936
rect 144736 3884 144788 3936
rect 454500 3884 454552 3936
rect 503720 3884 503772 3936
rect 533344 3884 533396 3936
rect 560852 3884 560904 3936
rect 25320 3816 25372 3868
rect 157984 3816 158036 3868
rect 450912 3816 450964 3868
rect 502432 3816 502484 3868
rect 534724 3816 534776 3868
rect 564440 3816 564492 3868
rect 20628 3748 20680 3800
rect 156604 3748 156656 3800
rect 383568 3748 383620 3800
rect 385776 3748 385828 3800
rect 401324 3748 401376 3800
rect 403624 3748 403676 3800
rect 408408 3748 408460 3800
rect 418804 3748 418856 3800
rect 447416 3748 447468 3800
rect 502616 3748 502668 3800
rect 518348 3748 518400 3800
rect 521660 3748 521712 3800
rect 536288 3748 536340 3800
rect 568028 3748 568080 3800
rect 15936 3680 15988 3732
rect 155224 3680 155276 3732
rect 193220 3680 193272 3732
rect 194416 3680 194468 3732
rect 251180 3680 251232 3732
rect 252376 3680 252428 3732
rect 267740 3680 267792 3732
rect 268476 3680 268528 3732
rect 284300 3680 284352 3732
rect 285036 3680 285088 3732
rect 365812 3680 365864 3732
rect 371884 3680 371936 3732
rect 415492 3680 415544 3732
rect 440884 3680 440936 3732
rect 443828 3680 443880 3732
rect 501052 3680 501104 3732
rect 516140 3680 516192 3732
rect 516324 3680 516376 3732
rect 536104 3680 536156 3732
rect 571524 3680 571576 3732
rect 5264 3612 5316 3664
rect 158168 3612 158220 3664
rect 160100 3612 160152 3664
rect 424140 3612 424192 3664
rect 440332 3612 440384 3664
rect 499856 3612 499908 3664
rect 511264 3612 511316 3664
rect 518992 3612 519044 3664
rect 537484 3612 537536 3664
rect 575112 3612 575164 3664
rect 11152 3544 11204 3596
rect 154028 3544 154080 3596
rect 156604 3544 156656 3596
rect 422392 3544 422444 3596
rect 436744 3544 436796 3596
rect 499672 3544 499724 3596
rect 507676 3544 507728 3596
rect 519176 3544 519228 3596
rect 526444 3544 526496 3596
rect 532516 3544 532568 3596
rect 541624 3544 541676 3596
rect 582196 3544 582248 3596
rect 572 3476 624 3528
rect 3424 3476 3476 3528
rect 24216 3476 24268 3528
rect 126244 3476 126296 3528
rect 153016 3476 153068 3528
rect 1676 3408 1728 3460
rect 10324 3408 10376 3460
rect 19432 3408 19484 3460
rect 124864 3408 124916 3460
rect 149520 3408 149572 3460
rect 415400 3476 415452 3528
rect 416688 3476 416740 3528
rect 423772 3476 423824 3528
rect 424968 3476 425020 3528
rect 433248 3476 433300 3528
rect 43076 3340 43128 3392
rect 131948 3340 132000 3392
rect 177856 3340 177908 3392
rect 178684 3340 178736 3392
rect 184940 3340 184992 3392
rect 186964 3340 187016 3392
rect 324412 3340 324464 3392
rect 325608 3340 325660 3392
rect 332600 3340 332652 3392
rect 333888 3340 333940 3392
rect 337476 3340 337528 3392
rect 340144 3340 340196 3392
rect 340880 3340 340932 3392
rect 342168 3340 342220 3392
rect 349160 3340 349212 3392
rect 350448 3340 350500 3392
rect 351644 3340 351696 3392
rect 353944 3340 353996 3392
rect 355232 3340 355284 3392
rect 356796 3340 356848 3392
rect 357440 3340 357492 3392
rect 358728 3340 358780 3392
rect 362316 3340 362368 3392
rect 363696 3340 363748 3392
rect 365720 3340 365772 3392
rect 367008 3340 367060 3392
rect 369400 3340 369452 3392
rect 370596 3340 370648 3392
rect 376484 3340 376536 3392
rect 378784 3340 378836 3392
rect 379980 3340 380032 3392
rect 382924 3340 382976 3392
rect 421288 3408 421340 3460
rect 426164 3408 426216 3460
rect 497096 3408 497148 3460
rect 498200 3476 498252 3528
rect 499028 3476 499080 3528
rect 504180 3476 504232 3528
rect 517520 3476 517572 3528
rect 521844 3476 521896 3528
rect 523132 3476 523184 3528
rect 526720 3476 526772 3528
rect 536104 3476 536156 3528
rect 538864 3476 538916 3528
rect 578608 3476 578660 3528
rect 498384 3408 498436 3460
rect 500592 3408 500644 3460
rect 516140 3408 516192 3460
rect 527916 3408 527968 3460
rect 539600 3408 539652 3460
rect 540244 3408 540296 3460
rect 581000 3408 581052 3460
rect 421104 3340 421156 3392
rect 448520 3340 448572 3392
rect 449808 3340 449860 3392
rect 472256 3340 472308 3392
rect 509424 3340 509476 3392
rect 530584 3340 530636 3392
rect 546684 3340 546736 3392
rect 4068 3272 4120 3324
rect 4804 3272 4856 3324
rect 46664 3272 46716 3324
rect 131764 3272 131816 3324
rect 319720 3272 319772 3324
rect 320824 3272 320876 3324
rect 340972 3272 341024 3324
rect 342904 3272 342956 3324
rect 475752 3272 475804 3324
rect 509700 3272 509752 3324
rect 529204 3272 529256 3324
rect 543188 3272 543240 3324
rect 77300 3204 77352 3256
rect 78220 3204 78272 3256
rect 102140 3204 102192 3256
rect 103336 3204 103388 3256
rect 121092 3204 121144 3256
rect 152464 3204 152516 3256
rect 305552 3204 305604 3256
rect 307024 3204 307076 3256
rect 479340 3204 479392 3256
rect 510620 3204 510672 3256
rect 13544 3136 13596 3188
rect 15844 3136 15896 3188
rect 124680 3136 124732 3188
rect 153844 3136 153896 3188
rect 390560 3136 390612 3188
rect 391848 3136 391900 3188
rect 397736 3136 397788 3188
rect 400956 3136 401008 3188
rect 489920 3136 489972 3188
rect 490748 3136 490800 3188
rect 497096 3136 497148 3188
rect 516508 3204 516560 3256
rect 514760 3136 514812 3188
rect 520372 3136 520424 3188
rect 525156 3136 525208 3188
rect 527824 3136 527876 3188
rect 309048 3000 309100 3052
rect 311164 3000 311216 3052
rect 522304 3000 522356 3052
rect 524236 3000 524288 3052
rect 8760 2932 8812 2984
rect 14464 2932 14516 2984
rect 523684 2932 523736 2984
rect 525432 2932 525484 2984
rect 326804 2864 326856 2916
rect 329104 2864 329156 2916
rect 390652 2864 390704 2916
rect 392584 2864 392636 2916
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 57426 559464 57482 559473
rect 57426 559399 57482 559408
rect 57440 558958 57468 559399
rect 10324 558952 10376 558958
rect 10324 558894 10376 558900
rect 57428 558952 57480 558958
rect 57428 558894 57480 558900
rect 3424 58676 3476 58682
rect 3424 58618 3476 58624
rect 2872 7608 2924 7614
rect 2872 7550 2924 7556
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 584 480 612 3470
rect 1676 3460 1728 3466
rect 1676 3402 1728 3408
rect 1688 480 1716 3402
rect 2884 480 2912 7550
rect 3436 3534 3464 58618
rect 4804 51740 4856 51746
rect 4804 51682 4856 51688
rect 3424 3528 3476 3534
rect 3424 3470 3476 3476
rect 4816 3330 4844 51682
rect 9956 6180 10008 6186
rect 9956 6122 10008 6128
rect 7656 4208 7708 4214
rect 7656 4150 7708 4156
rect 5264 3664 5316 3670
rect 5264 3606 5316 3612
rect 4068 3324 4120 3330
rect 4068 3266 4120 3272
rect 4804 3324 4856 3330
rect 4804 3266 4856 3272
rect 4080 480 4108 3266
rect 5276 480 5304 3606
rect 6458 3360 6514 3369
rect 6458 3295 6514 3304
rect 6472 480 6500 3295
rect 7668 480 7696 4150
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 8772 480 8800 2926
rect 9968 480 9996 6122
rect 10336 3466 10364 558894
rect 381912 59832 381964 59838
rect 57978 59800 58034 59809
rect 65890 59800 65946 59809
rect 57978 59735 58034 59744
rect 64788 59764 64840 59770
rect 11704 59424 11756 59430
rect 11704 59366 11756 59372
rect 11612 11756 11664 11762
rect 11612 11698 11664 11704
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 10324 3460 10376 3466
rect 10324 3402 10376 3408
rect 11164 480 11192 3538
rect 11624 490 11652 11698
rect 11716 4214 11744 59366
rect 57992 58682 58020 59735
rect 65890 59735 65892 59744
rect 64788 59706 64840 59712
rect 65944 59735 65946 59744
rect 67914 59800 67970 59809
rect 67914 59735 67970 59744
rect 68834 59800 68890 59809
rect 68834 59735 68890 59744
rect 69846 59800 69902 59809
rect 75642 59800 75698 59809
rect 69846 59735 69902 59744
rect 75472 59758 75642 59786
rect 65892 59706 65944 59712
rect 58622 59664 58678 59673
rect 58622 59599 58678 59608
rect 62026 59664 62082 59673
rect 62026 59599 62082 59608
rect 57980 58676 58032 58682
rect 57980 58618 58032 58624
rect 53840 57248 53892 57254
rect 53840 57190 53892 57196
rect 16580 55956 16632 55962
rect 16580 55898 16632 55904
rect 14464 50380 14516 50386
rect 14464 50322 14516 50328
rect 11704 4208 11756 4214
rect 11704 4150 11756 4156
rect 13544 3188 13596 3194
rect 13544 3130 13596 3136
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 11624 462 12020 490
rect 13556 480 13584 3130
rect 14476 2990 14504 50322
rect 15844 22772 15896 22778
rect 15844 22714 15896 22720
rect 14740 6248 14792 6254
rect 14740 6190 14792 6196
rect 14464 2984 14516 2990
rect 14464 2926 14516 2932
rect 14752 480 14780 6190
rect 15856 3194 15884 22714
rect 16592 16574 16620 55898
rect 26240 54596 26292 54602
rect 26240 54538 26292 54544
rect 17960 47592 18012 47598
rect 17960 47534 18012 47540
rect 16592 16546 17080 16574
rect 15936 3732 15988 3738
rect 15936 3674 15988 3680
rect 15844 3188 15896 3194
rect 15844 3130 15896 3136
rect 15948 480 15976 3674
rect 17052 480 17080 16546
rect 11992 354 12020 462
rect 12318 354 12430 480
rect 11992 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 47534
rect 22100 26920 22152 26926
rect 22100 26862 22152 26868
rect 22112 16574 22140 26862
rect 22112 16546 22600 16574
rect 21824 13116 21876 13122
rect 21824 13058 21876 13064
rect 20628 3800 20680 3806
rect 20628 3742 20680 3748
rect 19432 3460 19484 3466
rect 19432 3402 19484 3408
rect 19444 480 19472 3402
rect 20640 480 20668 3742
rect 21836 480 21864 13058
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 25320 3868 25372 3874
rect 25320 3810 25372 3816
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 24228 480 24256 3470
rect 25332 480 25360 3810
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 54538
rect 29000 53100 29052 53106
rect 29000 53042 29052 53048
rect 29012 16574 29040 53042
rect 52460 49020 52512 49026
rect 52460 48962 52512 48968
rect 44180 46232 44232 46238
rect 44180 46174 44232 46180
rect 37280 28280 37332 28286
rect 37280 28222 37332 28228
rect 30380 17264 30432 17270
rect 30380 17206 30432 17212
rect 30392 16574 30420 17206
rect 37292 16574 37320 28222
rect 44192 16574 44220 46174
rect 48320 18624 48372 18630
rect 48320 18566 48372 18572
rect 48332 16574 48360 18566
rect 52472 16574 52500 48962
rect 53852 16574 53880 57190
rect 56600 55888 56652 55894
rect 56600 55830 56652 55836
rect 55220 19984 55272 19990
rect 55220 19926 55272 19932
rect 55232 16574 55260 19926
rect 56612 16574 56640 55830
rect 29012 16546 30144 16574
rect 30392 16546 30880 16574
rect 37292 16546 38424 16574
rect 44192 16546 45048 16574
rect 48332 16546 48544 16574
rect 52472 16546 52592 16574
rect 53852 16546 54984 16574
rect 55232 16546 56088 16574
rect 56612 16546 56824 16574
rect 27712 6520 27764 6526
rect 27712 6462 27764 6468
rect 27724 480 27752 6462
rect 28908 3936 28960 3942
rect 28908 3878 28960 3884
rect 28920 480 28948 3878
rect 30116 480 30144 16546
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 33600 14476 33652 14482
rect 33600 14418 33652 14424
rect 32404 4004 32456 4010
rect 32404 3946 32456 3952
rect 32416 480 32444 3946
rect 33612 480 33640 14418
rect 34796 6656 34848 6662
rect 34796 6598 34848 6604
rect 34808 480 34836 6598
rect 37188 4820 37240 4826
rect 37188 4762 37240 4768
rect 35992 4072 36044 4078
rect 35992 4014 36044 4020
rect 36004 480 36032 4014
rect 37200 480 37228 4762
rect 38396 480 38424 16546
rect 41880 6724 41932 6730
rect 41880 6666 41932 6672
rect 40684 5092 40736 5098
rect 40684 5034 40736 5040
rect 39580 4140 39632 4146
rect 39580 4082 39632 4088
rect 39592 480 39620 4082
rect 40696 480 40724 5034
rect 41892 480 41920 6666
rect 44272 5160 44324 5166
rect 44272 5102 44324 5108
rect 43076 3392 43128 3398
rect 43076 3334 43128 3340
rect 43088 480 43116 3334
rect 44284 480 44312 5102
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31270 -960 31382 326
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 47860 8968 47912 8974
rect 47860 8910 47912 8916
rect 46664 3324 46716 3330
rect 46664 3266 46716 3272
rect 46676 480 46704 3266
rect 47872 480 47900 8910
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48516 354 48544 16546
rect 51080 10328 51132 10334
rect 51080 10270 51132 10276
rect 50160 6316 50212 6322
rect 50160 6258 50212 6264
rect 50172 480 50200 6258
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51092 354 51120 10270
rect 52564 480 52592 16546
rect 53748 6384 53800 6390
rect 53748 6326 53800 6332
rect 53760 480 53788 6326
rect 54956 480 54984 16546
rect 56060 480 56088 16546
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58440 7676 58492 7682
rect 58440 7618 58492 7624
rect 58452 480 58480 7618
rect 58636 7614 58664 59599
rect 61382 59528 61438 59537
rect 61382 59463 61438 59472
rect 61936 59492 61988 59498
rect 59360 59424 59412 59430
rect 59358 59392 59360 59401
rect 59412 59392 59414 59401
rect 59358 59327 59414 59336
rect 60740 54528 60792 54534
rect 60740 54470 60792 54476
rect 60752 16574 60780 54470
rect 60752 16546 60872 16574
rect 58624 7608 58676 7614
rect 58624 7550 58676 7556
rect 59636 4888 59688 4894
rect 59636 4830 59688 4836
rect 59648 480 59676 4830
rect 60844 480 60872 16546
rect 61396 11762 61424 59463
rect 61936 59434 61988 59440
rect 61948 55962 61976 59434
rect 62040 59401 62068 59599
rect 63958 59528 64014 59537
rect 63958 59463 63960 59472
rect 64012 59463 64014 59472
rect 63960 59434 64012 59440
rect 62026 59392 62082 59401
rect 62026 59327 62082 59336
rect 62762 59392 62818 59401
rect 62762 59327 62818 59336
rect 61936 55956 61988 55962
rect 61936 55898 61988 55904
rect 62776 13122 62804 59327
rect 64800 54602 64828 59706
rect 65982 59664 66038 59673
rect 65982 59599 66038 59608
rect 65890 59392 65946 59401
rect 65890 59327 65946 59336
rect 64788 54596 64840 54602
rect 64788 54538 64840 54544
rect 65904 51074 65932 59327
rect 65996 53106 66024 59599
rect 66902 59528 66958 59537
rect 66902 59463 66958 59472
rect 65984 53100 66036 53106
rect 65984 53042 66036 53048
rect 65536 51046 65932 51074
rect 65536 14482 65564 51046
rect 65524 14476 65576 14482
rect 65524 14418 65576 14424
rect 62764 13116 62816 13122
rect 62764 13058 62816 13064
rect 65064 13116 65116 13122
rect 65064 13058 65116 13064
rect 61568 11824 61620 11830
rect 61568 11766 61620 11772
rect 61384 11756 61436 11762
rect 61384 11698 61436 11704
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61580 354 61608 11766
rect 64328 6452 64380 6458
rect 64328 6394 64380 6400
rect 63224 4956 63276 4962
rect 63224 4898 63276 4904
rect 63236 480 63264 4898
rect 64340 480 64368 6394
rect 61998 354 62110 480
rect 61580 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 13058
rect 66720 5024 66772 5030
rect 66720 4966 66772 4972
rect 66732 480 66760 4966
rect 66916 4826 66944 59463
rect 67928 59401 67956 59735
rect 68466 59664 68522 59673
rect 68466 59599 68522 59608
rect 67914 59392 67970 59401
rect 67914 59327 67970 59336
rect 68282 59392 68338 59401
rect 68282 59327 68338 59336
rect 67640 29640 67692 29646
rect 67640 29582 67692 29588
rect 66904 4820 66956 4826
rect 66904 4762 66956 4768
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 29582
rect 68296 5098 68324 59327
rect 68480 5166 68508 59599
rect 68848 59537 68876 59735
rect 69860 59537 69888 59735
rect 71042 59664 71098 59673
rect 71042 59599 71098 59608
rect 74998 59664 75054 59673
rect 74998 59599 75054 59608
rect 68834 59528 68890 59537
rect 68834 59463 68890 59472
rect 69846 59528 69902 59537
rect 69846 59463 69902 59472
rect 69662 59392 69718 59401
rect 69662 59327 69718 59336
rect 69676 8974 69704 59327
rect 70400 31068 70452 31074
rect 70400 31010 70452 31016
rect 69664 8968 69716 8974
rect 69664 8910 69716 8916
rect 69112 8356 69164 8362
rect 69112 8298 69164 8304
rect 68468 5160 68520 5166
rect 68468 5102 68520 5108
rect 68284 5092 68336 5098
rect 68284 5034 68336 5040
rect 69124 480 69152 8298
rect 70412 6914 70440 31010
rect 71056 10334 71084 59599
rect 71778 59528 71834 59537
rect 71778 59463 71834 59472
rect 71792 57254 71820 59463
rect 75012 59401 75040 59599
rect 75472 59537 75500 59758
rect 75642 59735 75698 59744
rect 85026 59800 85082 59809
rect 85026 59735 85082 59744
rect 85210 59800 85266 59809
rect 85210 59735 85266 59744
rect 87970 59800 88026 59809
rect 87970 59735 88026 59744
rect 92294 59800 92350 59809
rect 92294 59735 92350 59744
rect 94134 59800 94190 59809
rect 97078 59800 97134 59809
rect 94134 59735 94190 59744
rect 94504 59764 94556 59770
rect 75642 59664 75698 59673
rect 75642 59599 75698 59608
rect 77574 59664 77630 59673
rect 78770 59664 78826 59673
rect 77574 59599 77630 59608
rect 78508 59622 78770 59650
rect 75458 59528 75514 59537
rect 75458 59463 75514 59472
rect 72422 59392 72478 59401
rect 72422 59327 72478 59336
rect 73802 59392 73858 59401
rect 73802 59327 73858 59336
rect 74998 59392 75054 59401
rect 74998 59327 75054 59336
rect 71780 57248 71832 57254
rect 71780 57190 71832 57196
rect 71044 10328 71096 10334
rect 71044 10270 71096 10276
rect 72436 7682 72464 59327
rect 73344 14544 73396 14550
rect 73344 14486 73396 14492
rect 72424 7676 72476 7682
rect 72424 7618 72476 7624
rect 72608 6928 72660 6934
rect 70412 6886 71544 6914
rect 70308 5092 70360 5098
rect 70308 5034 70360 5040
rect 70320 480 70348 5034
rect 71516 480 71544 6886
rect 72608 6870 72660 6876
rect 72620 480 72648 6870
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 14486
rect 73816 11830 73844 59327
rect 75182 59256 75238 59265
rect 75182 59191 75238 59200
rect 73804 11824 73856 11830
rect 73804 11766 73856 11772
rect 75196 8362 75224 59191
rect 75656 45554 75684 59599
rect 76562 59528 76618 59537
rect 76562 59463 76618 59472
rect 75920 57996 75972 58002
rect 75920 57938 75972 57944
rect 75380 45526 75684 45554
rect 75380 13122 75408 45526
rect 75368 13116 75420 13122
rect 75368 13058 75420 13064
rect 75184 8356 75236 8362
rect 75184 8298 75236 8304
rect 75000 6588 75052 6594
rect 75000 6530 75052 6536
rect 75012 480 75040 6530
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 57938
rect 76576 6934 76604 59463
rect 77588 59401 77616 59599
rect 77574 59392 77630 59401
rect 77574 59327 77630 59336
rect 78508 58002 78536 59622
rect 78770 59599 78826 59608
rect 79966 59664 80022 59673
rect 79966 59599 80022 59608
rect 84106 59664 84162 59673
rect 84106 59599 84162 59608
rect 78586 59392 78642 59401
rect 78586 59327 78642 59336
rect 78600 58018 78628 59327
rect 78496 57996 78548 58002
rect 78600 57990 78720 58018
rect 78496 57938 78548 57944
rect 77300 32428 77352 32434
rect 77300 32370 77352 32376
rect 76564 6928 76616 6934
rect 76564 6870 76616 6876
rect 77312 3262 77340 32370
rect 77392 21412 77444 21418
rect 77392 21354 77444 21360
rect 77300 3256 77352 3262
rect 77300 3198 77352 3204
rect 77404 480 77432 21354
rect 78692 16574 78720 57990
rect 78692 16546 79272 16574
rect 78220 3256 78272 3262
rect 78220 3198 78272 3204
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78232 354 78260 3198
rect 78558 354 78670 480
rect 78232 326 78670 354
rect 79244 354 79272 16546
rect 79980 8294 80008 59599
rect 81346 59528 81402 59537
rect 81346 59463 81402 59472
rect 80060 44872 80112 44878
rect 80060 44814 80112 44820
rect 80072 16574 80100 44814
rect 80072 16546 80928 16574
rect 79968 8288 80020 8294
rect 79968 8230 80020 8236
rect 80900 480 80928 16546
rect 81360 8362 81388 59463
rect 82542 59392 82598 59401
rect 82542 59327 82598 59336
rect 81440 22840 81492 22846
rect 81440 22782 81492 22788
rect 81452 16574 81480 22782
rect 81452 16546 81664 16574
rect 81348 8356 81400 8362
rect 81348 8298 81400 8304
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 82556 7682 82584 59327
rect 84120 10402 84148 59599
rect 85040 59362 85068 59735
rect 85224 59401 85252 59735
rect 85394 59528 85450 59537
rect 85394 59463 85450 59472
rect 86866 59528 86922 59537
rect 86866 59463 86922 59472
rect 85210 59392 85266 59401
rect 85028 59356 85080 59362
rect 85210 59327 85266 59336
rect 85028 59298 85080 59304
rect 85408 45554 85436 59463
rect 85316 45526 85436 45554
rect 85316 15910 85344 45526
rect 85580 35216 85632 35222
rect 85580 35158 85632 35164
rect 85592 16574 85620 35158
rect 85592 16546 85712 16574
rect 85304 15904 85356 15910
rect 85304 15846 85356 15852
rect 84108 10396 84160 10402
rect 84108 10338 84160 10344
rect 84200 10328 84252 10334
rect 84200 10270 84252 10276
rect 83280 8288 83332 8294
rect 83280 8230 83332 8236
rect 82544 7676 82596 7682
rect 82544 7618 82596 7624
rect 83292 480 83320 8230
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 10270
rect 85684 480 85712 16546
rect 86880 9042 86908 59463
rect 87984 57254 88012 59735
rect 89626 59528 89682 59537
rect 91282 59528 91338 59537
rect 89626 59463 89682 59472
rect 90836 59486 91282 59514
rect 88246 59392 88302 59401
rect 88246 59327 88302 59336
rect 89442 59392 89498 59401
rect 89442 59327 89498 59336
rect 87972 57248 88024 57254
rect 87972 57190 88024 57196
rect 86960 24132 87012 24138
rect 86960 24074 87012 24080
rect 86972 16574 87000 24074
rect 86972 16546 87552 16574
rect 86868 9036 86920 9042
rect 86868 8978 86920 8984
rect 86868 8356 86920 8362
rect 86868 8298 86920 8304
rect 86880 480 86908 8298
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87524 354 87552 16546
rect 88260 7614 88288 59327
rect 88340 36576 88392 36582
rect 88340 36518 88392 36524
rect 88352 16574 88380 36518
rect 88352 16546 89208 16574
rect 88248 7608 88300 7614
rect 88248 7550 88300 7556
rect 89180 480 89208 16546
rect 89456 13122 89484 59327
rect 89444 13116 89496 13122
rect 89444 13058 89496 13064
rect 89640 11762 89668 59463
rect 90836 59401 90864 59486
rect 91282 59463 91338 59472
rect 90822 59392 90878 59401
rect 89720 59356 89772 59362
rect 90822 59327 90878 59336
rect 89720 59298 89772 59304
rect 89732 16574 89760 59298
rect 92308 58818 92336 59735
rect 92386 59528 92442 59537
rect 92386 59463 92442 59472
rect 91008 58812 91060 58818
rect 91008 58754 91060 58760
rect 92296 58812 92348 58818
rect 92296 58754 92348 58760
rect 91020 17338 91048 58754
rect 91744 58540 91796 58546
rect 91744 58482 91796 58488
rect 91756 50386 91784 58482
rect 92400 57974 92428 59463
rect 93214 59392 93270 59401
rect 93214 59327 93270 59336
rect 92216 57946 92428 57974
rect 92216 51746 92244 57946
rect 92204 51740 92256 51746
rect 92204 51682 92256 51688
rect 93228 51074 93256 59327
rect 94148 58546 94176 59735
rect 97078 59735 97080 59744
rect 94504 59706 94556 59712
rect 97132 59735 97134 59744
rect 98090 59800 98146 59809
rect 100942 59800 100998 59809
rect 98090 59735 98146 59744
rect 98828 59764 98880 59770
rect 97080 59706 97132 59712
rect 94136 58540 94188 58546
rect 94136 58482 94188 58488
rect 93136 51046 93256 51074
rect 91744 50380 91796 50386
rect 91744 50322 91796 50328
rect 91100 25560 91152 25566
rect 91100 25502 91152 25508
rect 91008 17332 91060 17338
rect 91008 17274 91060 17280
rect 91112 16574 91140 25502
rect 93136 22778 93164 51046
rect 94516 26926 94544 59706
rect 97262 59664 97318 59673
rect 97262 59599 97318 59608
rect 95146 59528 95202 59537
rect 95146 59463 95202 59472
rect 95160 47598 95188 59463
rect 96066 59392 96122 59401
rect 96066 59327 96122 59336
rect 95148 47592 95200 47598
rect 95148 47534 95200 47540
rect 96080 45554 96108 59327
rect 95896 45526 96108 45554
rect 94504 26920 94556 26926
rect 94504 26862 94556 26868
rect 93124 22772 93176 22778
rect 93124 22714 93176 22720
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 89628 11756 89680 11762
rect 89628 11698 89680 11704
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 93952 7676 94004 7682
rect 93952 7618 94004 7624
rect 92756 4820 92808 4826
rect 92756 4762 92808 4768
rect 92768 480 92796 4762
rect 93964 480 93992 7618
rect 95896 6526 95924 45526
rect 97276 17270 97304 59599
rect 98104 59401 98132 59735
rect 107750 59800 107806 59809
rect 100942 59735 100944 59744
rect 98828 59706 98880 59712
rect 100996 59735 100998 59744
rect 105544 59764 105596 59770
rect 100944 59706 100996 59712
rect 110694 59800 110750 59809
rect 107750 59735 107752 59744
rect 105544 59706 105596 59712
rect 107804 59735 107806 59744
rect 108488 59764 108540 59770
rect 107752 59706 107804 59712
rect 115570 59800 115626 59809
rect 110694 59735 110696 59744
rect 108488 59706 108540 59712
rect 110748 59735 110750 59744
rect 113824 59764 113876 59770
rect 110696 59706 110748 59712
rect 115570 59735 115572 59744
rect 113824 59706 113876 59712
rect 115624 59735 115626 59744
rect 119710 59800 119766 59809
rect 127254 59800 127310 59809
rect 119710 59735 119766 59744
rect 124864 59764 124916 59770
rect 115572 59706 115624 59712
rect 98090 59392 98146 59401
rect 98090 59327 98146 59336
rect 98642 59392 98698 59401
rect 98642 59327 98698 59336
rect 97264 17264 97316 17270
rect 97264 17206 97316 17212
rect 97448 10396 97500 10402
rect 97448 10338 97500 10344
rect 96252 8968 96304 8974
rect 96252 8910 96304 8916
rect 95884 6520 95936 6526
rect 95884 6462 95936 6468
rect 95148 5160 95200 5166
rect 95148 5102 95200 5108
rect 95160 480 95188 5102
rect 96264 480 96292 8910
rect 97460 480 97488 10338
rect 98656 6662 98684 59327
rect 98840 28286 98868 59706
rect 101586 59528 101642 59537
rect 101586 59463 101642 59472
rect 104898 59528 104954 59537
rect 104898 59463 104954 59472
rect 101402 59392 101458 59401
rect 101402 59327 101458 59336
rect 100022 59256 100078 59265
rect 100022 59191 100078 59200
rect 98828 28280 98880 28286
rect 98828 28222 98880 28228
rect 99840 14476 99892 14482
rect 99840 14418 99892 14424
rect 98644 6656 98696 6662
rect 98644 6598 98696 6604
rect 98644 5364 98696 5370
rect 98644 5306 98696 5312
rect 98656 4962 98684 5306
rect 98736 5228 98788 5234
rect 98736 5170 98788 5176
rect 98644 4956 98696 4962
rect 98644 4898 98696 4904
rect 98748 2666 98776 5170
rect 98656 2638 98776 2666
rect 98656 480 98684 2638
rect 99852 480 99880 14418
rect 100036 6730 100064 59191
rect 100760 57248 100812 57254
rect 100760 57190 100812 57196
rect 100024 6724 100076 6730
rect 100024 6666 100076 6672
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 100772 354 100800 57190
rect 101416 18630 101444 59327
rect 101600 46238 101628 59463
rect 104912 59430 104940 59463
rect 103520 59424 103572 59430
rect 102782 59392 102838 59401
rect 102782 59327 102838 59336
rect 103518 59392 103520 59401
rect 104900 59424 104952 59430
rect 103572 59392 103574 59401
rect 104900 59366 104952 59372
rect 103518 59327 103574 59336
rect 102796 49026 102824 59327
rect 104346 59256 104402 59265
rect 104346 59191 104402 59200
rect 104162 59120 104218 59129
rect 104162 59055 104218 59064
rect 102784 49020 102836 49026
rect 102784 48962 102836 48968
rect 102140 47592 102192 47598
rect 102140 47534 102192 47540
rect 101588 46232 101640 46238
rect 101588 46174 101640 46180
rect 101404 18624 101456 18630
rect 101404 18566 101456 18572
rect 102152 3262 102180 47534
rect 104072 15904 104124 15910
rect 104072 15846 104124 15852
rect 102232 5296 102284 5302
rect 102232 5238 102284 5244
rect 102140 3256 102192 3262
rect 102140 3198 102192 3204
rect 102244 480 102272 5238
rect 103336 3256 103388 3262
rect 103336 3198 103388 3204
rect 103348 480 103376 3198
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 15846
rect 104176 4894 104204 59055
rect 104360 19990 104388 59191
rect 104900 58676 104952 58682
rect 104900 58618 104952 58624
rect 104348 19984 104400 19990
rect 104348 19926 104400 19932
rect 104912 16574 104940 58618
rect 104912 16546 105492 16574
rect 104164 4888 104216 4894
rect 104164 4830 104216 4836
rect 105464 3482 105492 16546
rect 105556 5370 105584 59706
rect 108302 59528 108358 59537
rect 108302 59463 108358 59472
rect 107106 59256 107162 59265
rect 107106 59191 107162 59200
rect 107120 45554 107148 59191
rect 106936 45526 107148 45554
rect 106280 18624 106332 18630
rect 106280 18566 106332 18572
rect 106292 16574 106320 18566
rect 106292 16546 106504 16574
rect 105544 5364 105596 5370
rect 105544 5306 105596 5312
rect 105464 3454 105768 3482
rect 105740 480 105768 3454
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 106936 5030 106964 45526
rect 108120 9036 108172 9042
rect 108120 8978 108172 8984
rect 106924 5024 106976 5030
rect 106924 4966 106976 4972
rect 108132 480 108160 8978
rect 108316 5098 108344 59463
rect 108500 14550 108528 59706
rect 111246 59528 111302 59537
rect 111246 59463 111302 59472
rect 113272 59492 113324 59498
rect 109682 59392 109738 59401
rect 109682 59327 109738 59336
rect 111062 59392 111118 59401
rect 111062 59327 111118 59336
rect 109696 21418 109724 59327
rect 110420 50380 110472 50386
rect 110420 50322 110472 50328
rect 109684 21412 109736 21418
rect 109684 21354 109736 21360
rect 110432 16574 110460 50322
rect 110432 16546 110552 16574
rect 109040 15904 109092 15910
rect 109040 15846 109092 15852
rect 108488 14544 108540 14550
rect 108488 14486 108540 14492
rect 108304 5092 108356 5098
rect 108304 5034 108356 5040
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109052 354 109080 15846
rect 110524 480 110552 16546
rect 111076 10334 111104 59327
rect 111260 44878 111288 59463
rect 113272 59434 113324 59440
rect 113284 59401 113312 59434
rect 112442 59392 112498 59401
rect 112442 59327 112498 59336
rect 113270 59392 113326 59401
rect 113270 59327 113326 59336
rect 111248 44872 111300 44878
rect 111248 44814 111300 44820
rect 112456 24138 112484 59327
rect 113836 25566 113864 59706
rect 117502 59664 117558 59673
rect 118698 59664 118754 59673
rect 117502 59599 117558 59608
rect 118620 59622 118698 59650
rect 114650 59528 114706 59537
rect 114650 59463 114652 59472
rect 114704 59463 114706 59472
rect 116582 59528 116638 59537
rect 116582 59463 116638 59472
rect 114652 59434 114704 59440
rect 115202 59392 115258 59401
rect 115202 59327 115258 59336
rect 115754 59392 115810 59401
rect 115754 59327 115810 59336
rect 113824 25560 113876 25566
rect 113824 25502 113876 25508
rect 112444 24132 112496 24138
rect 112444 24074 112496 24080
rect 113180 19984 113232 19990
rect 113180 19926 113232 19932
rect 113192 16574 113220 19926
rect 113192 16546 114048 16574
rect 111064 10328 111116 10334
rect 111064 10270 111116 10276
rect 111616 7608 111668 7614
rect 111616 7550 111668 7556
rect 111628 480 111656 7550
rect 112812 4888 112864 4894
rect 112812 4830 112864 4836
rect 112824 480 112852 4830
rect 114020 480 114048 16546
rect 114744 11756 114796 11762
rect 114744 11698 114796 11704
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 114756 354 114784 11698
rect 115216 5166 115244 59327
rect 115768 45554 115796 59327
rect 115400 45526 115796 45554
rect 115400 5234 115428 45526
rect 116596 5302 116624 59463
rect 117516 59401 117544 59599
rect 117502 59392 117558 59401
rect 117502 59327 117558 59336
rect 117962 59392 118018 59401
rect 117962 59327 118018 59336
rect 117976 15910 118004 59327
rect 118620 58682 118648 59622
rect 118698 59599 118754 59608
rect 119434 59664 119490 59673
rect 119434 59599 119490 59608
rect 118608 58676 118660 58682
rect 118608 58618 118660 58624
rect 119448 45554 119476 59599
rect 119724 59401 119752 59735
rect 131118 59800 131174 59809
rect 127254 59735 127256 59744
rect 124864 59706 124916 59712
rect 127308 59735 127310 59744
rect 129004 59764 129056 59770
rect 127256 59706 127308 59712
rect 134062 59800 134118 59809
rect 131118 59735 131120 59744
rect 129004 59706 129056 59712
rect 131172 59735 131174 59744
rect 131764 59764 131816 59770
rect 131120 59706 131172 59712
rect 137006 59800 137062 59809
rect 134062 59735 134064 59744
rect 131764 59706 131816 59712
rect 134116 59735 134118 59744
rect 135168 59764 135220 59770
rect 134064 59706 134116 59712
rect 137006 59735 137008 59744
rect 135168 59706 135220 59712
rect 137060 59735 137062 59744
rect 140870 59800 140926 59809
rect 143814 59800 143870 59809
rect 140870 59735 140926 59744
rect 141424 59764 141476 59770
rect 137008 59706 137060 59712
rect 123484 59628 123536 59634
rect 123484 59570 123536 59576
rect 120906 59528 120962 59537
rect 120906 59463 120962 59472
rect 119710 59392 119766 59401
rect 119710 59327 119766 59336
rect 120722 59392 120778 59401
rect 120722 59327 120778 59336
rect 119356 45526 119476 45554
rect 117964 15904 118016 15910
rect 117964 15846 118016 15852
rect 118792 13116 118844 13122
rect 118792 13058 118844 13064
rect 117596 7608 117648 7614
rect 117596 7550 117648 7556
rect 116584 5296 116636 5302
rect 116584 5238 116636 5244
rect 115388 5228 115440 5234
rect 115388 5170 115440 5176
rect 115204 5160 115256 5166
rect 115204 5102 115256 5108
rect 116400 4276 116452 4282
rect 116400 4218 116452 4224
rect 116412 480 116440 4218
rect 117608 480 117636 7550
rect 118804 480 118832 13058
rect 119356 4894 119384 45526
rect 119344 4888 119396 4894
rect 119344 4830 119396 4836
rect 120736 4214 120764 59327
rect 120920 4282 120948 59463
rect 122746 59392 122802 59401
rect 122746 59327 122802 59336
rect 123022 59392 123078 59401
rect 123022 59327 123078 59336
rect 121460 17332 121512 17338
rect 121460 17274 121512 17280
rect 121472 16574 121500 17274
rect 121472 16546 122328 16574
rect 120908 4276 120960 4282
rect 120908 4218 120960 4224
rect 119896 4208 119948 4214
rect 119896 4150 119948 4156
rect 120724 4208 120776 4214
rect 120724 4150 120776 4156
rect 119908 480 119936 4150
rect 121092 3256 121144 3262
rect 121092 3198 121144 3204
rect 121104 480 121132 3198
rect 122300 480 122328 16546
rect 122760 4162 122788 59327
rect 123036 59242 123064 59327
rect 123298 59256 123354 59265
rect 123036 59214 123298 59242
rect 123298 59191 123354 59200
rect 123496 6186 123524 59570
rect 123484 6180 123536 6186
rect 123484 6122 123536 6128
rect 122760 4134 123064 4162
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123036 354 123064 4134
rect 124876 3466 124904 59706
rect 125322 59664 125378 59673
rect 125322 59599 125324 59608
rect 125376 59599 125378 59608
rect 125324 59570 125376 59576
rect 125322 59528 125378 59537
rect 125322 59463 125378 59472
rect 127806 59528 127862 59537
rect 127806 59463 127862 59472
rect 125336 45554 125364 59463
rect 126242 59392 126298 59401
rect 126242 59327 126298 59336
rect 127622 59392 127678 59401
rect 127622 59327 127678 59336
rect 125060 45526 125364 45554
rect 125060 6254 125088 45526
rect 125048 6248 125100 6254
rect 125048 6190 125100 6196
rect 125876 4888 125928 4894
rect 125876 4830 125928 4836
rect 124864 3460 124916 3466
rect 124864 3402 124916 3408
rect 124680 3188 124732 3194
rect 124680 3130 124732 3136
rect 124692 480 124720 3130
rect 125888 480 125916 4830
rect 126256 3534 126284 59327
rect 126980 28416 127032 28422
rect 126980 28358 127032 28364
rect 126244 3528 126296 3534
rect 126244 3470 126296 3476
rect 126992 480 127020 28358
rect 127532 13116 127584 13122
rect 127532 13058 127584 13064
rect 127544 3482 127572 13058
rect 127636 4010 127664 59327
rect 127624 4004 127676 4010
rect 127624 3946 127676 3952
rect 127820 3942 127848 59463
rect 129016 4078 129044 59706
rect 130474 59256 130530 59265
rect 130474 59191 130530 59200
rect 130488 45554 130516 59191
rect 130396 45526 130516 45554
rect 130292 10328 130344 10334
rect 130292 10270 130344 10276
rect 129372 4956 129424 4962
rect 129372 4898 129424 4904
rect 129004 4072 129056 4078
rect 129004 4014 129056 4020
rect 127808 3936 127860 3942
rect 127808 3878 127860 3884
rect 127544 3454 128216 3482
rect 128188 480 128216 3454
rect 129384 480 129412 4898
rect 130304 3482 130332 10270
rect 130396 4146 130424 45526
rect 131120 33856 131172 33862
rect 131120 33798 131172 33804
rect 131132 16574 131160 33798
rect 131132 16546 131344 16574
rect 130384 4140 130436 4146
rect 130384 4082 130436 4088
rect 130304 3454 130608 3482
rect 130580 480 130608 3454
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 131776 3330 131804 59706
rect 131946 59528 132002 59537
rect 131946 59463 132002 59472
rect 134522 59528 134578 59537
rect 134522 59463 134578 59472
rect 131960 3398 131988 59463
rect 133142 59392 133198 59401
rect 133142 59327 133198 59336
rect 133156 6322 133184 59327
rect 133880 11756 133932 11762
rect 133880 11698 133932 11704
rect 133144 6316 133196 6322
rect 133144 6258 133196 6264
rect 132960 5024 133012 5030
rect 132960 4966 133012 4972
rect 131948 3392 132000 3398
rect 131948 3334 132000 3340
rect 131764 3324 131816 3330
rect 131764 3266 131816 3272
rect 132972 480 133000 4966
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 133892 354 133920 11698
rect 134536 6390 134564 59463
rect 135180 55894 135208 59706
rect 140042 59664 140098 59673
rect 140042 59599 140098 59608
rect 137282 59528 137338 59537
rect 137282 59463 137338 59472
rect 135902 59392 135958 59401
rect 135902 59327 135958 59336
rect 135168 55888 135220 55894
rect 135168 55830 135220 55836
rect 135916 54534 135944 59327
rect 135904 54528 135956 54534
rect 135904 54470 135956 54476
rect 135260 49020 135312 49026
rect 135260 48962 135312 48968
rect 134524 6384 134576 6390
rect 134524 6326 134576 6332
rect 135272 480 135300 48962
rect 136640 25764 136692 25770
rect 136640 25706 136692 25712
rect 136652 16574 136680 25706
rect 136652 16546 137232 16574
rect 136456 7676 136508 7682
rect 136456 7618 136508 7624
rect 136468 480 136496 7618
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 137296 6458 137324 59463
rect 137466 59392 137522 59401
rect 137466 59327 137522 59336
rect 137480 29646 137508 59327
rect 138662 59256 138718 59265
rect 138662 59191 138718 59200
rect 138676 31074 138704 59191
rect 138664 31068 138716 31074
rect 138664 31010 138716 31016
rect 137468 29640 137520 29646
rect 137468 29582 137520 29588
rect 138848 15904 138900 15910
rect 138848 15846 138900 15852
rect 137284 6452 137336 6458
rect 137284 6394 137336 6400
rect 138860 480 138888 15846
rect 140056 6594 140084 59599
rect 140884 59401 140912 59735
rect 147678 59800 147734 59809
rect 143814 59735 143816 59744
rect 141424 59706 141476 59712
rect 143868 59735 143870 59744
rect 145564 59764 145616 59770
rect 143816 59706 143868 59712
rect 150622 59800 150678 59809
rect 147678 59735 147680 59744
rect 145564 59706 145616 59712
rect 147732 59735 147734 59744
rect 148324 59764 148376 59770
rect 147680 59706 147732 59712
rect 157430 59800 157486 59809
rect 150622 59735 150624 59744
rect 148324 59706 148376 59712
rect 150676 59735 150678 59744
rect 155224 59764 155276 59770
rect 150624 59706 150676 59712
rect 163318 59800 163374 59809
rect 157430 59735 157432 59744
rect 155224 59706 155276 59712
rect 157484 59735 157486 59744
rect 160744 59764 160796 59770
rect 157432 59706 157484 59712
rect 163318 59735 163320 59744
rect 160744 59706 160796 59712
rect 163372 59735 163374 59744
rect 168286 59800 168342 59809
rect 168286 59735 168342 59744
rect 170126 59800 170182 59809
rect 170126 59735 170182 59744
rect 173990 59800 174046 59809
rect 176934 59800 176990 59809
rect 173990 59735 174046 59744
rect 176396 59758 176934 59786
rect 163320 59706 163372 59712
rect 140870 59392 140926 59401
rect 140870 59327 140926 59336
rect 140780 31204 140832 31210
rect 140780 31146 140832 31152
rect 140792 16574 140820 31146
rect 141436 22846 141464 59706
rect 141606 59528 141662 59537
rect 141606 59463 141662 59472
rect 144366 59528 144422 59537
rect 144366 59463 144422 59472
rect 141620 32434 141648 59463
rect 142802 59392 142858 59401
rect 142802 59327 142858 59336
rect 144182 59392 144238 59401
rect 144182 59327 144238 59336
rect 142160 53168 142212 53174
rect 142160 53110 142212 53116
rect 141608 32428 141660 32434
rect 141608 32370 141660 32376
rect 141424 22840 141476 22846
rect 141424 22782 141476 22788
rect 140792 16546 141280 16574
rect 140044 6588 140096 6594
rect 140044 6530 140096 6536
rect 140044 5092 140096 5098
rect 140044 5034 140096 5040
rect 140056 480 140084 5034
rect 141252 480 141280 16546
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142172 354 142200 53110
rect 142816 35222 142844 59327
rect 143540 46368 143592 46374
rect 143540 46310 143592 46316
rect 142804 35216 142856 35222
rect 142804 35158 142856 35164
rect 143552 3942 143580 46310
rect 143632 9036 143684 9042
rect 143632 8978 143684 8984
rect 143540 3936 143592 3942
rect 143540 3878 143592 3884
rect 143644 3482 143672 8978
rect 144196 4758 144224 59327
rect 144380 36582 144408 59463
rect 144368 36576 144420 36582
rect 144368 36518 144420 36524
rect 144920 29640 144972 29646
rect 144920 29582 144972 29588
rect 144932 16574 144960 29582
rect 144932 16546 145512 16574
rect 144184 4752 144236 4758
rect 144184 4694 144236 4700
rect 144736 3936 144788 3942
rect 144736 3878 144788 3884
rect 143552 3454 143672 3482
rect 143552 480 143580 3454
rect 144748 480 144776 3878
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 145576 8974 145604 59706
rect 147034 59256 147090 59265
rect 147034 59191 147090 59200
rect 147048 45554 147076 59191
rect 146956 45526 147076 45554
rect 146956 14482 146984 45526
rect 147680 45008 147732 45014
rect 147680 44950 147732 44956
rect 147692 16574 147720 44950
rect 148336 18630 148364 59706
rect 148506 59528 148562 59537
rect 148506 59463 148562 59472
rect 151266 59528 151322 59537
rect 154486 59528 154542 59537
rect 151266 59463 151322 59472
rect 152464 59492 152516 59498
rect 148520 47598 148548 59463
rect 149702 59392 149758 59401
rect 149702 59327 149758 59336
rect 151082 59392 151138 59401
rect 151082 59327 151138 59336
rect 149716 50386 149744 59327
rect 150440 58676 150492 58682
rect 150440 58618 150492 58624
rect 149704 50380 149756 50386
rect 149704 50322 149756 50328
rect 148508 47592 148560 47598
rect 148508 47534 148560 47540
rect 148324 18624 148376 18630
rect 148324 18566 148376 18572
rect 150452 16574 150480 58618
rect 147692 16546 147904 16574
rect 150452 16546 150664 16574
rect 147128 14544 147180 14550
rect 147128 14486 147180 14492
rect 146944 14476 146996 14482
rect 146944 14418 146996 14424
rect 145564 8968 145616 8974
rect 145564 8910 145616 8916
rect 147140 480 147168 14486
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 149520 3460 149572 3466
rect 149520 3402 149572 3408
rect 149532 480 149560 3402
rect 150636 480 150664 16546
rect 151096 7614 151124 59327
rect 151280 19990 151308 59463
rect 154486 59463 154488 59472
rect 152464 59434 152516 59440
rect 154540 59463 154542 59472
rect 154488 59434 154540 59440
rect 151268 19984 151320 19990
rect 151268 19926 151320 19932
rect 151820 13320 151872 13326
rect 151820 13262 151872 13268
rect 151084 7608 151136 7614
rect 151084 7550 151136 7556
rect 151832 480 151860 13262
rect 152476 3262 152504 59434
rect 153842 59256 153898 59265
rect 153842 59191 153898 59200
rect 153016 3528 153068 3534
rect 153016 3470 153068 3476
rect 152464 3256 152516 3262
rect 152464 3198 152516 3204
rect 153028 480 153056 3470
rect 153856 3194 153884 59191
rect 154026 59120 154082 59129
rect 154026 59055 154082 59064
rect 154040 3602 154068 59055
rect 155132 13388 155184 13394
rect 155132 13330 155184 13336
rect 154212 6180 154264 6186
rect 154212 6122 154264 6128
rect 154028 3596 154080 3602
rect 154028 3538 154080 3544
rect 153844 3188 153896 3194
rect 153844 3130 153896 3136
rect 154224 480 154252 6122
rect 155144 3482 155172 13330
rect 155236 3738 155264 59706
rect 156602 59664 156658 59673
rect 156602 59599 156658 59608
rect 159364 59628 159416 59634
rect 156616 3806 156644 59599
rect 159364 59570 159416 59576
rect 157982 59528 158038 59537
rect 157982 59463 158038 59472
rect 157800 7608 157852 7614
rect 157800 7550 157852 7556
rect 156604 3800 156656 3806
rect 156604 3742 156656 3748
rect 155224 3732 155276 3738
rect 155224 3674 155276 3680
rect 156604 3596 156656 3602
rect 156604 3538 156656 3544
rect 155144 3454 155448 3482
rect 155420 480 155448 3454
rect 156616 480 156644 3538
rect 157812 480 157840 7550
rect 157996 3874 158024 59463
rect 158166 59392 158222 59401
rect 158166 59327 158222 59336
rect 157984 3868 158036 3874
rect 157984 3810 158036 3816
rect 158180 3670 158208 59327
rect 158904 13456 158956 13462
rect 158904 13398 158956 13404
rect 158168 3664 158220 3670
rect 158168 3606 158220 3612
rect 158916 480 158944 13398
rect 159376 3369 159404 59570
rect 160756 4962 160784 59706
rect 161294 59664 161350 59673
rect 161294 59599 161296 59608
rect 161348 59599 161350 59608
rect 161296 59570 161348 59576
rect 161294 59528 161350 59537
rect 161294 59463 161350 59472
rect 163502 59528 163558 59537
rect 167182 59528 167238 59537
rect 163502 59463 163558 59472
rect 165068 59492 165120 59498
rect 161308 45554 161336 59463
rect 162122 59392 162178 59401
rect 162122 59327 162178 59336
rect 161480 57384 161532 57390
rect 161480 57326 161532 57332
rect 160940 45526 161336 45554
rect 160744 4956 160796 4962
rect 160744 4898 160796 4904
rect 160940 4894 160968 45526
rect 161492 16574 161520 57326
rect 161492 16546 162072 16574
rect 161296 6248 161348 6254
rect 161296 6190 161348 6196
rect 160928 4888 160980 4894
rect 160928 4830 160980 4836
rect 160100 3664 160152 3670
rect 160100 3606 160152 3612
rect 159362 3360 159418 3369
rect 159362 3295 159418 3304
rect 160112 480 160140 3606
rect 161308 480 161336 6190
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 16546
rect 162136 5030 162164 59327
rect 163516 7682 163544 59463
rect 167182 59463 167184 59472
rect 165068 59434 165120 59440
rect 167236 59463 167238 59472
rect 167184 59434 167236 59440
rect 164882 59392 164938 59401
rect 164882 59327 164938 59336
rect 163688 13184 163740 13190
rect 163688 13126 163740 13132
rect 163504 7676 163556 7682
rect 163504 7618 163556 7624
rect 162124 5024 162176 5030
rect 162124 4966 162176 4972
rect 163700 480 163728 13126
rect 164896 5098 164924 59327
rect 165080 9042 165108 59434
rect 166446 59392 166502 59401
rect 166446 59327 166502 59336
rect 166460 51074 166488 59327
rect 167642 59256 167698 59265
rect 167642 59191 167698 59200
rect 166276 51046 166488 51074
rect 166276 14550 166304 51046
rect 167000 39364 167052 39370
rect 167000 39306 167052 39312
rect 167012 16574 167040 39306
rect 167012 16546 167224 16574
rect 166264 14544 166316 14550
rect 166264 14486 166316 14492
rect 166080 10396 166132 10402
rect 166080 10338 166132 10344
rect 165068 9036 165120 9042
rect 165068 8978 165120 8984
rect 164884 5092 164936 5098
rect 164884 5034 164936 5040
rect 164884 4208 164936 4214
rect 164884 4150 164936 4156
rect 164896 480 164924 4150
rect 166092 480 166120 10338
rect 167196 480 167224 16546
rect 167656 6186 167684 59191
rect 168300 58682 168328 59735
rect 169114 59664 169170 59673
rect 169114 59599 169170 59608
rect 168380 59356 168432 59362
rect 168380 59298 168432 59304
rect 168288 58676 168340 58682
rect 168288 58618 168340 58624
rect 167644 6180 167696 6186
rect 167644 6122 167696 6128
rect 168392 480 168420 59298
rect 169128 45554 169156 59599
rect 170140 59401 170168 59735
rect 173162 59664 173218 59673
rect 173162 59599 173218 59608
rect 170586 59528 170642 59537
rect 170586 59463 170642 59472
rect 170126 59392 170182 59401
rect 170126 59327 170182 59336
rect 170402 59392 170458 59401
rect 170402 59327 170458 59336
rect 169036 45526 169156 45554
rect 169036 7614 169064 45526
rect 169760 40724 169812 40730
rect 169760 40666 169812 40672
rect 169772 16574 169800 40666
rect 169772 16546 170352 16574
rect 169576 10532 169628 10538
rect 169576 10474 169628 10480
rect 169024 7608 169076 7614
rect 169024 7550 169076 7556
rect 169588 480 169616 10474
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 16546
rect 170416 4214 170444 59327
rect 170600 6254 170628 59463
rect 172704 10464 172756 10470
rect 172704 10406 172756 10412
rect 170588 6248 170640 6254
rect 170588 6190 170640 6196
rect 170404 4208 170456 4214
rect 170404 4150 170456 4156
rect 171968 4208 172020 4214
rect 171968 4150 172020 4156
rect 171980 480 172008 4150
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 172716 354 172744 10406
rect 173176 4214 173204 59599
rect 174004 59362 174032 59735
rect 175094 59528 175150 59537
rect 175094 59463 175150 59472
rect 174910 59392 174966 59401
rect 173992 59356 174044 59362
rect 174910 59327 174966 59336
rect 173992 59298 174044 59304
rect 173900 42084 173952 42090
rect 173900 42026 173952 42032
rect 173164 4208 173216 4214
rect 173164 4150 173216 4156
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173912 354 173940 42026
rect 174924 5574 174952 59327
rect 175108 9674 175136 59463
rect 176396 59401 176424 59758
rect 180798 59800 180854 59809
rect 176934 59735 176990 59744
rect 179328 59764 179380 59770
rect 186594 59800 186650 59809
rect 180798 59735 180800 59744
rect 179328 59706 179380 59712
rect 180852 59735 180854 59744
rect 184756 59764 184808 59770
rect 180800 59706 180852 59712
rect 186594 59735 186596 59744
rect 184756 59706 184808 59712
rect 186648 59735 186650 59744
rect 188342 59800 188398 59809
rect 188618 59800 188674 59809
rect 188398 59758 188618 59786
rect 188342 59735 188398 59744
rect 194598 59800 194654 59809
rect 188618 59735 188674 59744
rect 193140 59770 193260 59786
rect 193140 59764 193272 59770
rect 193140 59758 193220 59764
rect 186596 59706 186648 59712
rect 177762 59528 177818 59537
rect 177762 59463 177818 59472
rect 176382 59392 176438 59401
rect 176382 59327 176438 59336
rect 176566 59392 176622 59401
rect 176566 59327 176622 59336
rect 175108 9646 175320 9674
rect 175292 6914 175320 9646
rect 175292 6886 175504 6914
rect 174912 5568 174964 5574
rect 174912 5510 174964 5516
rect 175476 480 175504 6886
rect 176580 4894 176608 59327
rect 176660 32632 176712 32638
rect 176660 32574 176712 32580
rect 176568 4888 176620 4894
rect 176568 4830 176620 4836
rect 176672 480 176700 32574
rect 177776 6322 177804 59463
rect 177946 59392 178002 59401
rect 177946 59327 178002 59336
rect 177764 6316 177816 6322
rect 177764 6258 177816 6264
rect 177960 4826 177988 59327
rect 178684 37936 178736 37942
rect 178684 37878 178736 37884
rect 177948 4820 178000 4826
rect 177948 4762 178000 4768
rect 178696 3398 178724 37878
rect 179340 7750 179368 59706
rect 180706 59528 180762 59537
rect 180706 59463 180762 59472
rect 181810 59528 181866 59537
rect 181810 59463 181866 59472
rect 180248 10600 180300 10606
rect 180248 10542 180300 10548
rect 179328 7744 179380 7750
rect 179328 7686 179380 7692
rect 179052 5568 179104 5574
rect 179052 5510 179104 5516
rect 177856 3392 177908 3398
rect 177856 3334 177908 3340
rect 178684 3392 178736 3398
rect 178684 3334 178736 3340
rect 177868 480 177896 3334
rect 179064 480 179092 5510
rect 180260 480 180288 10542
rect 180720 9110 180748 59463
rect 180800 43444 180852 43450
rect 180800 43386 180852 43392
rect 180812 16574 180840 43386
rect 180812 16546 181024 16574
rect 180708 9104 180760 9110
rect 180708 9046 180760 9052
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 173134 -960 173246 326
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181824 6254 181852 59463
rect 181994 59392 182050 59401
rect 181994 59327 182050 59336
rect 182008 7682 182036 59327
rect 183466 59256 183522 59265
rect 183466 59191 183522 59200
rect 181996 7676 182048 7682
rect 181996 7618 182048 7624
rect 181812 6248 181864 6254
rect 181812 6190 181864 6196
rect 183480 6186 183508 59191
rect 184570 59120 184626 59129
rect 184570 59055 184626 59064
rect 183744 10668 183796 10674
rect 183744 10610 183796 10616
rect 183468 6180 183520 6186
rect 183468 6122 183520 6128
rect 182548 4888 182600 4894
rect 182548 4830 182600 4836
rect 182560 480 182588 4830
rect 183756 480 183784 10610
rect 184584 9042 184612 59055
rect 184768 17270 184796 59706
rect 187330 59664 187386 59673
rect 187330 59599 187386 59608
rect 193034 59664 193090 59673
rect 193034 59599 193090 59608
rect 186226 59392 186282 59401
rect 186226 59327 186282 59336
rect 186240 18630 186268 59327
rect 186964 55956 187016 55962
rect 186964 55898 187016 55904
rect 186228 18624 186280 18630
rect 186228 18566 186280 18572
rect 184756 17264 184808 17270
rect 184756 17206 184808 17212
rect 186872 10736 186924 10742
rect 186872 10678 186924 10684
rect 184572 9036 184624 9042
rect 184572 8978 184624 8984
rect 186136 6316 186188 6322
rect 186136 6258 186188 6264
rect 184940 3392 184992 3398
rect 184940 3334 184992 3340
rect 184952 480 184980 3334
rect 186148 480 186176 6258
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 181414 -960 181526 326
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 10678
rect 186976 3398 187004 55898
rect 187344 7614 187372 59599
rect 188986 59528 189042 59537
rect 188986 59463 189042 59472
rect 191470 59528 191526 59537
rect 191470 59463 191526 59472
rect 187514 59256 187570 59265
rect 187514 59191 187570 59200
rect 187528 19990 187556 59191
rect 187700 51808 187752 51814
rect 187700 51750 187752 51756
rect 187516 19984 187568 19990
rect 187516 19926 187568 19932
rect 187712 16574 187740 51750
rect 189000 21418 189028 59463
rect 190460 58812 190512 58818
rect 190460 58754 190512 58760
rect 188988 21412 189040 21418
rect 188988 21354 189040 21360
rect 187712 16546 188568 16574
rect 187332 7608 187384 7614
rect 187332 7550 187384 7556
rect 186964 3392 187016 3398
rect 186964 3334 187016 3340
rect 188540 480 188568 16546
rect 189724 4820 189776 4826
rect 189724 4762 189776 4768
rect 189736 480 189764 4762
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190472 354 190500 58754
rect 191484 5166 191512 59463
rect 191654 59392 191710 59401
rect 191654 59327 191710 59336
rect 191472 5160 191524 5166
rect 191472 5102 191524 5108
rect 191668 5098 191696 59327
rect 193048 58682 193076 59599
rect 193036 58676 193088 58682
rect 193036 58618 193088 58624
rect 191840 28348 191892 28354
rect 191840 28290 191892 28296
rect 191852 16574 191880 28290
rect 191852 16546 192064 16574
rect 191656 5092 191708 5098
rect 191656 5034 191708 5040
rect 192036 480 192064 16546
rect 193140 8974 193168 59758
rect 193220 59706 193272 59712
rect 193772 59764 193824 59770
rect 193772 59706 193824 59712
rect 194428 59758 194598 59786
rect 193784 59673 193812 59706
rect 193770 59664 193826 59673
rect 193770 59599 193826 59608
rect 193220 53304 193272 53310
rect 193220 53246 193272 53252
rect 193128 8968 193180 8974
rect 193128 8910 193180 8916
rect 193232 3738 193260 53246
rect 194428 51074 194456 59758
rect 204166 59800 204222 59809
rect 194598 59735 194654 59744
rect 202788 59764 202840 59770
rect 204166 59735 204168 59744
rect 202788 59706 202840 59712
rect 204220 59735 204222 59744
rect 206742 59800 206798 59809
rect 209962 59800 210018 59809
rect 209700 59770 209962 59786
rect 206742 59735 206798 59744
rect 208032 59764 208084 59770
rect 204168 59706 204220 59712
rect 194598 59664 194654 59673
rect 194598 59599 194654 59608
rect 195886 59664 195942 59673
rect 200302 59664 200358 59673
rect 200040 59634 200302 59650
rect 195886 59599 195942 59608
rect 198372 59628 198424 59634
rect 194612 57974 194640 59599
rect 194244 51046 194456 51074
rect 194520 57946 194640 57974
rect 194244 22778 194272 51046
rect 194520 45554 194548 57946
rect 194600 57316 194652 57322
rect 194600 57258 194652 57264
rect 194428 45526 194548 45554
rect 194428 24138 194456 45526
rect 194416 24132 194468 24138
rect 194416 24074 194468 24080
rect 194232 22772 194284 22778
rect 194232 22714 194284 22720
rect 194612 16574 194640 57258
rect 194612 16546 195192 16574
rect 193312 7744 193364 7750
rect 193312 7686 193364 7692
rect 193220 3732 193272 3738
rect 193220 3674 193272 3680
rect 193324 3482 193352 7686
rect 194416 3732 194468 3738
rect 194416 3674 194468 3680
rect 193232 3454 193352 3482
rect 193232 480 193260 3454
rect 194428 480 194456 3674
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 195900 5030 195928 59599
rect 198372 59570 198424 59576
rect 200028 59628 200302 59634
rect 200080 59622 200302 59628
rect 200302 59599 200358 59608
rect 200028 59570 200080 59576
rect 197266 59528 197322 59537
rect 197266 59463 197322 59472
rect 196808 9104 196860 9110
rect 196808 9046 196860 9052
rect 195888 5024 195940 5030
rect 195888 4966 195940 4972
rect 196820 480 196848 9046
rect 197280 4962 197308 59463
rect 197360 33992 197412 33998
rect 197360 33934 197412 33940
rect 197372 16574 197400 33934
rect 197372 16546 197952 16574
rect 197268 4956 197320 4962
rect 197268 4898 197320 4904
rect 197924 480 197952 16546
rect 198384 4894 198412 59570
rect 201314 59528 201370 59537
rect 201144 59486 201314 59514
rect 198554 59392 198610 59401
rect 198554 59327 198610 59336
rect 200026 59392 200082 59401
rect 200026 59327 200082 59336
rect 198568 25566 198596 59327
rect 198740 44872 198792 44878
rect 198740 44814 198792 44820
rect 198556 25560 198608 25566
rect 198556 25502 198608 25508
rect 198372 4888 198424 4894
rect 198372 4830 198424 4836
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 44814
rect 200040 26926 200068 59327
rect 200028 26920 200080 26926
rect 200028 26862 200080 26868
rect 200304 6248 200356 6254
rect 200304 6190 200356 6196
rect 200316 480 200344 6190
rect 201144 4826 201172 59486
rect 201314 59463 201370 59472
rect 201314 59392 201370 59401
rect 201314 59327 201370 59336
rect 201328 29714 201356 59327
rect 201500 51876 201552 51882
rect 201500 51818 201552 51824
rect 201316 29708 201368 29714
rect 201316 29650 201368 29656
rect 201132 4820 201184 4826
rect 201132 4762 201184 4768
rect 201512 480 201540 51818
rect 201592 32496 201644 32502
rect 201592 32438 201644 32444
rect 201604 16574 201632 32438
rect 202800 31074 202828 59706
rect 204166 59664 204222 59673
rect 204166 59599 204222 59608
rect 204180 51950 204208 59599
rect 205546 59528 205602 59537
rect 205546 59463 205602 59472
rect 204260 56024 204312 56030
rect 204260 55966 204312 55972
rect 204168 51944 204220 51950
rect 204168 51886 204220 51892
rect 202788 31068 202840 31074
rect 202788 31010 202840 31016
rect 204272 16574 204300 55966
rect 201604 16546 202736 16574
rect 204272 16546 205128 16574
rect 202708 480 202736 16546
rect 203892 7676 203944 7682
rect 203892 7618 203944 7624
rect 203904 480 203932 7618
rect 205100 480 205128 16546
rect 205560 6594 205588 59463
rect 206756 56098 206784 59735
rect 208032 59706 208084 59712
rect 209688 59764 209962 59770
rect 209740 59758 209962 59764
rect 212906 59800 212962 59809
rect 209962 59735 210018 59744
rect 210976 59764 211028 59770
rect 209688 59706 209740 59712
rect 212906 59735 212908 59744
rect 210976 59706 211028 59712
rect 212960 59735 212962 59744
rect 215850 59800 215906 59809
rect 215850 59735 215906 59744
rect 219530 59800 219586 59809
rect 222658 59800 222714 59809
rect 219530 59735 219586 59744
rect 220544 59764 220596 59770
rect 212908 59706 212960 59712
rect 206926 59392 206982 59401
rect 206926 59327 206982 59336
rect 206744 56092 206796 56098
rect 206744 56034 206796 56040
rect 206192 14476 206244 14482
rect 206192 14418 206244 14424
rect 205548 6588 205600 6594
rect 205548 6530 205600 6536
rect 206204 480 206232 14418
rect 206940 6526 206968 59327
rect 208044 47802 208072 59706
rect 209686 59392 209742 59401
rect 209686 59327 209742 59336
rect 208214 59256 208270 59265
rect 208214 59191 208270 59200
rect 208228 49230 208256 59191
rect 208400 54732 208452 54738
rect 208400 54674 208452 54680
rect 208216 49224 208268 49230
rect 208216 49166 208268 49172
rect 208032 47796 208084 47802
rect 208032 47738 208084 47744
rect 208412 16574 208440 54674
rect 208412 16546 208624 16574
rect 206928 6520 206980 6526
rect 206928 6462 206980 6468
rect 207388 6180 207440 6186
rect 207388 6122 207440 6128
rect 207400 480 207428 6122
rect 208596 480 208624 16546
rect 209700 6458 209728 59327
rect 210790 59256 210846 59265
rect 210790 59191 210846 59200
rect 209780 14544 209832 14550
rect 209780 14486 209832 14492
rect 209688 6452 209740 6458
rect 209688 6394 209740 6400
rect 209792 480 209820 14486
rect 210804 6390 210832 59191
rect 210792 6384 210844 6390
rect 210792 6326 210844 6332
rect 210988 6322 211016 59706
rect 215206 59664 215262 59673
rect 215206 59599 215262 59608
rect 213550 59528 213606 59537
rect 213550 59463 213606 59472
rect 212446 59256 212502 59265
rect 212446 59191 212502 59200
rect 211160 17400 211212 17406
rect 211160 17342 211212 17348
rect 211172 16574 211200 17342
rect 211172 16546 211752 16574
rect 211068 9036 211120 9042
rect 211068 8978 211120 8984
rect 210976 6316 211028 6322
rect 210976 6258 211028 6264
rect 211080 3482 211108 8978
rect 210988 3454 211108 3482
rect 210988 480 211016 3454
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 212460 6254 212488 59191
rect 213368 14612 213420 14618
rect 213368 14554 213420 14560
rect 212448 6248 212500 6254
rect 212448 6190 212500 6196
rect 213380 480 213408 14554
rect 213564 6186 213592 59463
rect 213734 59256 213790 59265
rect 213734 59191 213790 59200
rect 213748 43586 213776 59191
rect 213736 43580 213788 43586
rect 213736 43522 213788 43528
rect 215220 35358 215248 59599
rect 215864 59401 215892 59735
rect 219544 59537 219572 59735
rect 222658 59735 222660 59744
rect 220544 59706 220596 59712
rect 222712 59735 222714 59744
rect 223670 59800 223726 59809
rect 229466 59800 229522 59809
rect 223670 59735 223726 59744
rect 227536 59764 227588 59770
rect 222660 59706 222712 59712
rect 216586 59528 216642 59537
rect 216586 59463 216642 59472
rect 219530 59528 219586 59537
rect 219530 59463 219586 59472
rect 215850 59392 215906 59401
rect 215850 59327 215906 59336
rect 215300 57452 215352 57458
rect 215300 57394 215352 57400
rect 215208 35352 215260 35358
rect 215208 35294 215260 35300
rect 213920 17264 213972 17270
rect 213920 17206 213972 17212
rect 213932 16574 213960 17206
rect 213932 16546 214512 16574
rect 213552 6180 213604 6186
rect 213552 6122 213604 6128
rect 214484 480 214512 16546
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 57394
rect 216600 36718 216628 59463
rect 217874 59392 217930 59401
rect 217874 59327 217930 59336
rect 219346 59392 219402 59401
rect 219346 59327 219402 59336
rect 217690 59256 217746 59265
rect 217690 59191 217746 59200
rect 217704 38078 217732 59191
rect 217888 39574 217916 59327
rect 218060 50584 218112 50590
rect 218060 50526 218112 50532
rect 217876 39568 217928 39574
rect 217876 39510 217928 39516
rect 217692 38072 217744 38078
rect 217692 38014 217744 38020
rect 216588 36712 216640 36718
rect 216588 36654 216640 36660
rect 216864 14680 216916 14686
rect 216864 14622 216916 14628
rect 216876 480 216904 14622
rect 218072 11830 218100 50526
rect 219360 40934 219388 59327
rect 220556 45082 220584 59706
rect 220818 59664 220874 59673
rect 220818 59599 220874 59608
rect 223486 59664 223542 59673
rect 223486 59599 223542 59608
rect 220726 59528 220782 59537
rect 220726 59463 220782 59472
rect 220544 45076 220596 45082
rect 220544 45018 220596 45024
rect 220740 42294 220768 59463
rect 220832 59401 220860 59599
rect 220818 59392 220874 59401
rect 220818 59327 220874 59336
rect 222106 59392 222162 59401
rect 222106 59327 222162 59336
rect 222120 46442 222148 59327
rect 222108 46436 222160 46442
rect 222108 46378 222160 46384
rect 220728 42288 220780 42294
rect 220728 42230 220780 42236
rect 219348 40928 219400 40934
rect 219348 40870 219400 40876
rect 223500 33930 223528 59599
rect 223684 59401 223712 59735
rect 232410 59800 232466 59809
rect 229466 59735 229468 59744
rect 227536 59706 227588 59712
rect 229520 59735 229522 59744
rect 230112 59764 230164 59770
rect 229468 59706 229520 59712
rect 240138 59800 240194 59809
rect 232410 59735 232412 59744
rect 230112 59706 230164 59712
rect 232464 59735 232466 59744
rect 238668 59764 238720 59770
rect 232412 59706 232464 59712
rect 248970 59800 249026 59809
rect 240138 59735 240140 59744
rect 238668 59706 238720 59712
rect 240192 59735 240194 59744
rect 246672 59764 246724 59770
rect 240140 59706 240192 59712
rect 252834 59800 252890 59809
rect 248970 59735 248972 59744
rect 246672 59706 246724 59712
rect 249024 59735 249026 59744
rect 250996 59764 251048 59770
rect 248972 59706 249024 59712
rect 252834 59735 252836 59744
rect 250996 59706 251048 59712
rect 252888 59735 252890 59744
rect 254306 59800 254362 59809
rect 254306 59735 254362 59744
rect 257986 59800 258042 59809
rect 257986 59735 258042 59744
rect 259642 59800 259698 59809
rect 259642 59735 259698 59744
rect 264794 59800 264850 59809
rect 264794 59735 264850 59744
rect 264978 59800 265034 59809
rect 273258 59800 273314 59809
rect 264978 59735 265034 59744
rect 271788 59764 271840 59770
rect 252836 59706 252888 59712
rect 224774 59528 224830 59537
rect 226522 59528 226578 59537
rect 224774 59463 224830 59472
rect 226076 59486 226522 59514
rect 223670 59392 223726 59401
rect 223670 59327 223726 59336
rect 224590 59392 224646 59401
rect 224590 59327 224646 59336
rect 223488 33924 223540 33930
rect 223488 33866 223540 33872
rect 224604 32570 224632 59327
rect 224788 49162 224816 59463
rect 226076 59401 226104 59486
rect 226522 59463 226578 59472
rect 226062 59392 226118 59401
rect 226062 59327 226118 59336
rect 226246 59392 226302 59401
rect 226246 59327 226302 59336
rect 224776 49156 224828 49162
rect 224776 49098 224828 49104
rect 226260 47734 226288 59327
rect 227350 59256 227406 59265
rect 227350 59191 227406 59200
rect 226248 47728 226300 47734
rect 226248 47670 226300 47676
rect 224592 32564 224644 32570
rect 224592 32506 224644 32512
rect 227364 28490 227392 59191
rect 227548 50522 227576 59706
rect 229006 59392 229062 59401
rect 229006 59327 229062 59336
rect 227536 50516 227588 50522
rect 227536 50458 227588 50464
rect 227352 28484 227404 28490
rect 227352 28426 227404 28432
rect 226340 21616 226392 21622
rect 226340 21558 226392 21564
rect 222200 20120 222252 20126
rect 222200 20062 222252 20068
rect 218152 18624 218204 18630
rect 218152 18566 218204 18572
rect 218060 11824 218112 11830
rect 218060 11766 218112 11772
rect 218164 6914 218192 18566
rect 222212 16574 222240 20062
rect 224960 19984 225012 19990
rect 224960 19926 225012 19932
rect 224972 16574 225000 19926
rect 222212 16546 222792 16574
rect 224972 16546 225184 16574
rect 219992 14748 220044 14754
rect 219992 14690 220044 14696
rect 219256 11824 219308 11830
rect 219256 11766 219308 11772
rect 218072 6886 218192 6914
rect 218072 480 218100 6886
rect 219268 480 219296 11766
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 14690
rect 221556 7608 221608 7614
rect 221556 7550 221608 7556
rect 221568 480 221596 7550
rect 222764 480 222792 16546
rect 223580 14816 223632 14822
rect 223580 14758 223632 14764
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 220422 -960 220534 326
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223592 354 223620 14758
rect 225156 480 225184 16546
rect 226352 480 226380 21558
rect 227720 21412 227772 21418
rect 227720 21354 227772 21360
rect 227732 16574 227760 21354
rect 227732 16546 228312 16574
rect 227536 14884 227588 14890
rect 227536 14826 227588 14832
rect 227548 480 227576 14826
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16546
rect 229020 7682 229048 59327
rect 230124 35290 230152 59706
rect 233146 59664 233202 59673
rect 233146 59599 233202 59608
rect 230294 59256 230350 59265
rect 230294 59191 230350 59200
rect 231766 59256 231822 59265
rect 231766 59191 231822 59200
rect 230308 43518 230336 59191
rect 230296 43512 230348 43518
rect 230296 43454 230348 43460
rect 230112 35284 230164 35290
rect 230112 35226 230164 35232
rect 229100 18760 229152 18766
rect 229100 18702 229152 18708
rect 229112 16574 229140 18702
rect 229112 16546 229416 16574
rect 229008 7676 229060 7682
rect 229008 7618 229060 7624
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 16546
rect 231032 14952 231084 14958
rect 231032 14894 231084 14900
rect 231044 480 231072 14894
rect 231780 7614 231808 59191
rect 231860 58676 231912 58682
rect 231860 58618 231912 58624
rect 231768 7608 231820 7614
rect 231768 7550 231820 7556
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 58618
rect 233160 36650 233188 59599
rect 234250 59528 234306 59537
rect 237378 59528 237434 59537
rect 234250 59463 234306 59472
rect 235908 59492 235960 59498
rect 233148 36644 233200 36650
rect 233148 36586 233200 36592
rect 234264 17338 234292 59463
rect 237378 59463 237380 59472
rect 235908 59434 235960 59440
rect 237432 59463 237434 59472
rect 237380 59434 237432 59440
rect 234434 59392 234490 59401
rect 234434 59327 234490 59336
rect 234448 38010 234476 59327
rect 235920 39438 235948 59434
rect 237010 59256 237066 59265
rect 237010 59191 237066 59200
rect 237024 40798 237052 59191
rect 237286 59120 237342 59129
rect 237286 59055 237342 59064
rect 237300 45554 237328 59055
rect 237380 58744 237432 58750
rect 237380 58686 237432 58692
rect 237208 45526 237328 45554
rect 237208 42158 237236 45526
rect 237196 42152 237248 42158
rect 237196 42094 237248 42100
rect 237012 40792 237064 40798
rect 237012 40734 237064 40740
rect 235908 39432 235960 39438
rect 235908 39374 235960 39380
rect 234436 38004 234488 38010
rect 234436 37946 234488 37952
rect 236000 22976 236052 22982
rect 236000 22918 236052 22924
rect 234252 17332 234304 17338
rect 234252 17274 234304 17280
rect 236012 16574 236040 22918
rect 237392 16574 237420 58686
rect 238680 18698 238708 59706
rect 244094 59664 244150 59673
rect 242808 59628 242860 59634
rect 244094 59599 244096 59608
rect 242808 59570 242860 59576
rect 244148 59599 244150 59608
rect 244096 59570 244148 59576
rect 240046 59528 240102 59537
rect 240046 59463 240102 59472
rect 241426 59528 241482 59537
rect 241426 59463 241482 59472
rect 240060 44946 240088 59463
rect 241242 59392 241298 59401
rect 241242 59327 241298 59336
rect 240048 44940 240100 44946
rect 240048 44882 240100 44888
rect 241256 21486 241284 59327
rect 241244 21480 241296 21486
rect 241244 21422 241296 21428
rect 241440 20058 241468 59463
rect 242820 46306 242848 59570
rect 244094 59528 244150 59537
rect 246026 59528 246082 59537
rect 244094 59463 244150 59472
rect 244188 59492 244240 59498
rect 244108 51074 244136 59463
rect 246026 59463 246028 59472
rect 244188 59434 244240 59440
rect 246080 59463 246082 59472
rect 246028 59434 246080 59440
rect 244200 54670 244228 59434
rect 245566 59392 245622 59401
rect 245566 59327 245622 59336
rect 244188 54664 244240 54670
rect 244188 54606 244240 54612
rect 243924 51046 244136 51074
rect 242808 46300 242860 46306
rect 242808 46242 242860 46248
rect 241520 46232 241572 46238
rect 241520 46174 241572 46180
rect 241428 20052 241480 20058
rect 241428 19994 241480 20000
rect 238668 18692 238720 18698
rect 238668 18634 238720 18640
rect 241532 16574 241560 46174
rect 243924 22846 243952 51046
rect 244280 47660 244332 47666
rect 244280 47602 244332 47608
rect 243912 22840 243964 22846
rect 243912 22782 243964 22788
rect 244292 16574 244320 47602
rect 245580 24206 245608 59327
rect 245568 24200 245620 24206
rect 245568 24142 245620 24148
rect 245660 22772 245712 22778
rect 245660 22714 245712 22720
rect 245672 16574 245700 22714
rect 236012 16546 236592 16574
rect 237392 16546 237696 16574
rect 241532 16546 241744 16574
rect 244292 16546 245240 16574
rect 245672 16546 245976 16574
rect 234620 15020 234672 15026
rect 234620 14962 234672 14968
rect 233424 11824 233476 11830
rect 233424 11766 233476 11772
rect 233436 480 233464 11766
rect 234632 480 234660 14962
rect 235816 5160 235868 5166
rect 235816 5102 235868 5108
rect 235828 480 235856 5102
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 16546
rect 240140 11892 240192 11898
rect 240140 11834 240192 11840
rect 239312 5092 239364 5098
rect 239312 5034 239364 5040
rect 239324 480 239352 5034
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240152 354 240180 11834
rect 241716 480 241744 16546
rect 242900 8968 242952 8974
rect 242900 8910 242952 8916
rect 242912 480 242940 8910
rect 244096 7744 244148 7750
rect 244096 7686 244148 7692
rect 244108 480 244136 7686
rect 245212 480 245240 16546
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 16546
rect 246684 9110 246712 59706
rect 250902 59664 250958 59673
rect 250902 59599 250958 59608
rect 250810 59528 250866 59537
rect 250810 59463 250866 59472
rect 248326 59392 248382 59401
rect 248326 59327 248382 59336
rect 249706 59392 249762 59401
rect 249706 59327 249762 59336
rect 246854 59256 246910 59265
rect 246854 59191 246910 59200
rect 246868 25702 246896 59191
rect 248340 26994 248368 59327
rect 248328 26988 248380 26994
rect 248328 26930 248380 26936
rect 246856 25696 246908 25702
rect 246856 25638 246908 25644
rect 248420 25628 248472 25634
rect 248420 25570 248472 25576
rect 247040 24336 247092 24342
rect 247040 24278 247092 24284
rect 247052 16574 247080 24278
rect 247052 16546 247632 16574
rect 246672 9104 246724 9110
rect 246672 9046 246724 9052
rect 247604 480 247632 16546
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248432 354 248460 25570
rect 249720 9042 249748 59327
rect 249800 24132 249852 24138
rect 249800 24074 249852 24080
rect 249812 16574 249840 24074
rect 249812 16546 250024 16574
rect 249708 9036 249760 9042
rect 249708 8978 249760 8984
rect 249996 480 250024 16546
rect 250824 8974 250852 59463
rect 250916 59401 250944 59599
rect 250902 59392 250958 59401
rect 250902 59327 250958 59336
rect 251008 29782 251036 59706
rect 252466 59392 252522 59401
rect 252466 59327 252522 59336
rect 253754 59392 253810 59401
rect 253754 59327 253810 59336
rect 251180 54596 251232 54602
rect 251180 54538 251232 54544
rect 250996 29776 251048 29782
rect 250996 29718 251048 29724
rect 250812 8968 250864 8974
rect 250812 8910 250864 8916
rect 251192 3738 251220 54538
rect 252480 49094 252508 59327
rect 253572 58540 253624 58546
rect 253572 58482 253624 58488
rect 252468 49088 252520 49094
rect 252468 49030 252520 49036
rect 253584 31142 253612 58482
rect 253768 47598 253796 59327
rect 254320 58546 254348 59735
rect 255226 59664 255282 59673
rect 255226 59599 255282 59608
rect 254308 58540 254360 58546
rect 254308 58482 254360 58488
rect 253756 47592 253808 47598
rect 253756 47534 253808 47540
rect 255240 35222 255268 59599
rect 256606 59528 256662 59537
rect 256606 59463 256662 59472
rect 256620 36582 256648 59463
rect 257710 59392 257766 59401
rect 257710 59327 257766 59336
rect 256608 36576 256660 36582
rect 256608 36518 256660 36524
rect 255228 35216 255280 35222
rect 255228 35158 255280 35164
rect 253572 31136 253624 31142
rect 253572 31078 253624 31084
rect 257724 17270 257752 59327
rect 258000 53242 258028 59735
rect 259366 59664 259422 59673
rect 259366 59599 259422 59608
rect 257988 53236 258040 53242
rect 257988 53178 258040 53184
rect 259380 18630 259408 59599
rect 259656 59401 259684 59735
rect 263506 59664 263562 59673
rect 263336 59622 263506 59650
rect 260746 59528 260802 59537
rect 260746 59463 260802 59472
rect 259642 59392 259698 59401
rect 259642 59327 259698 59336
rect 260654 59392 260710 59401
rect 260654 59327 260710 59336
rect 260668 51074 260696 59327
rect 260576 51046 260696 51074
rect 259460 25560 259512 25566
rect 259460 25502 259512 25508
rect 259368 18624 259420 18630
rect 259368 18566 259420 18572
rect 257712 17264 257764 17270
rect 257712 17206 257764 17212
rect 255872 15972 255924 15978
rect 255872 15914 255924 15920
rect 254216 12028 254268 12034
rect 254216 11970 254268 11976
rect 251272 11960 251324 11966
rect 251272 11902 251324 11908
rect 251180 3732 251232 3738
rect 251180 3674 251232 3680
rect 251284 3482 251312 11902
rect 253480 5024 253532 5030
rect 253480 4966 253532 4972
rect 252376 3732 252428 3738
rect 252376 3674 252428 3680
rect 251192 3454 251312 3482
rect 251192 480 251220 3454
rect 252388 480 252416 3674
rect 253492 480 253520 4966
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 11970
rect 255884 480 255912 15914
rect 258264 12096 258316 12102
rect 258264 12038 258316 12044
rect 257068 4956 257120 4962
rect 257068 4898 257120 4904
rect 257080 480 257108 4898
rect 258276 480 258304 12038
rect 259472 11694 259500 25502
rect 260576 21418 260604 51046
rect 260564 21412 260616 21418
rect 260564 21354 260616 21360
rect 260760 19990 260788 59463
rect 260840 52012 260892 52018
rect 260840 51954 260892 51960
rect 260748 19984 260800 19990
rect 260748 19926 260800 19932
rect 260852 16574 260880 51954
rect 263336 24138 263364 59622
rect 263506 59599 263562 59608
rect 263506 59528 263562 59537
rect 263506 59463 263562 59472
rect 263324 24132 263376 24138
rect 263324 24074 263376 24080
rect 263520 22778 263548 59463
rect 264808 58682 264836 59735
rect 264992 59537 265020 59735
rect 280066 59800 280122 59809
rect 273258 59735 273260 59744
rect 271788 59706 271840 59712
rect 273312 59735 273314 59744
rect 278688 59764 278740 59770
rect 273260 59706 273312 59712
rect 280066 59735 280068 59744
rect 278688 59706 278740 59712
rect 280120 59735 280122 59744
rect 281078 59800 281134 59809
rect 289818 59800 289874 59809
rect 281078 59735 281134 59744
rect 287704 59764 287756 59770
rect 280068 59706 280120 59712
rect 267646 59664 267702 59673
rect 270314 59664 270370 59673
rect 267646 59599 267702 59608
rect 269028 59628 269080 59634
rect 264978 59528 265034 59537
rect 264978 59463 265034 59472
rect 267462 59528 267518 59537
rect 267462 59463 267518 59472
rect 264886 59392 264942 59401
rect 264886 59327 264942 59336
rect 264796 58676 264848 58682
rect 264796 58618 264848 58624
rect 264900 25566 264928 59327
rect 267476 45554 267504 59463
rect 267554 59392 267610 59401
rect 267554 59327 267610 59336
rect 267384 45526 267504 45554
rect 264980 27056 265032 27062
rect 264980 26998 265032 27004
rect 264888 25560 264940 25566
rect 264888 25502 264940 25508
rect 263508 22772 263560 22778
rect 263508 22714 263560 22720
rect 260852 16546 261800 16574
rect 259552 16040 259604 16046
rect 259552 15982 259604 15988
rect 259460 11688 259512 11694
rect 259460 11630 259512 11636
rect 259564 6914 259592 15982
rect 260656 11688 260708 11694
rect 260656 11630 260708 11636
rect 259472 6886 259592 6914
rect 259472 480 259500 6886
rect 260668 480 260696 11630
rect 261772 480 261800 16546
rect 262496 16108 262548 16114
rect 262496 16050 262548 16056
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16050
rect 264152 4888 264204 4894
rect 264152 4830 264204 4836
rect 264164 480 264192 4830
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 264992 354 265020 26998
rect 266544 16176 266596 16182
rect 266544 16118 266596 16124
rect 266556 480 266584 16118
rect 267384 5302 267412 45526
rect 267372 5296 267424 5302
rect 267372 5238 267424 5244
rect 267568 5234 267596 59327
rect 267660 57254 267688 59599
rect 270314 59599 270316 59608
rect 269028 59570 269080 59576
rect 270368 59599 270370 59608
rect 270316 59570 270368 59576
rect 267740 58880 267792 58886
rect 267740 58822 267792 58828
rect 267648 57248 267700 57254
rect 267648 57190 267700 57196
rect 267556 5228 267608 5234
rect 267556 5170 267608 5176
rect 267752 3738 267780 58822
rect 267832 26920 267884 26926
rect 267832 26862 267884 26868
rect 267740 3732 267792 3738
rect 267740 3674 267792 3680
rect 267844 3482 267872 26862
rect 269040 5166 269068 59570
rect 270314 59528 270370 59537
rect 270314 59463 270370 59472
rect 270130 59256 270186 59265
rect 270130 59191 270186 59200
rect 270040 16244 270092 16250
rect 270040 16186 270092 16192
rect 269028 5160 269080 5166
rect 269028 5102 269080 5108
rect 268476 3732 268528 3738
rect 268476 3674 268528 3680
rect 267752 3454 267872 3482
rect 267752 480 267780 3454
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268488 354 268516 3674
rect 270052 480 270080 16186
rect 270144 5098 270172 59191
rect 270328 26926 270356 59463
rect 270316 26920 270368 26926
rect 270316 26862 270368 26868
rect 270132 5092 270184 5098
rect 270132 5034 270184 5040
rect 271800 5030 271828 59706
rect 277122 59664 277178 59673
rect 275928 59628 275980 59634
rect 277122 59599 277124 59608
rect 275928 59570 275980 59576
rect 277176 59599 277178 59608
rect 277124 59570 277176 59576
rect 273166 59528 273222 59537
rect 273166 59463 273222 59472
rect 274454 59528 274510 59537
rect 274454 59463 274510 59472
rect 271880 29844 271932 29850
rect 271880 29786 271932 29792
rect 271892 16574 271920 29786
rect 273180 28286 273208 59463
rect 274270 59392 274326 59401
rect 274270 59327 274326 59336
rect 273168 28280 273220 28286
rect 273168 28222 273220 28228
rect 271892 16546 272472 16574
rect 271788 5024 271840 5030
rect 271788 4966 271840 4972
rect 271236 4820 271288 4826
rect 271236 4762 271288 4768
rect 271248 480 271276 4762
rect 272444 480 272472 16546
rect 273260 16312 273312 16318
rect 273260 16254 273312 16260
rect 268814 354 268926 480
rect 268488 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273272 354 273300 16254
rect 274284 4894 274312 59327
rect 274468 4962 274496 59463
rect 274640 29708 274692 29714
rect 274640 29650 274692 29656
rect 274652 16574 274680 29650
rect 274652 16546 274864 16574
rect 274456 4956 274508 4962
rect 274456 4898 274508 4904
rect 274272 4888 274324 4894
rect 274272 4830 274324 4836
rect 274836 480 274864 16546
rect 275940 4826 275968 59570
rect 277306 59528 277362 59537
rect 277306 59463 277362 59472
rect 277122 59392 277178 59401
rect 277122 59327 277178 59336
rect 276020 56160 276072 56166
rect 276020 56102 276072 56108
rect 275928 4820 275980 4826
rect 275928 4762 275980 4768
rect 276032 480 276060 56102
rect 277136 45554 277164 59327
rect 277320 55894 277348 59463
rect 277308 55888 277360 55894
rect 277308 55830 277360 55836
rect 277044 45526 277164 45554
rect 277044 29714 277072 45526
rect 278700 31074 278728 59706
rect 280066 59664 280122 59673
rect 280066 59599 280122 59608
rect 279882 59256 279938 59265
rect 279882 59191 279938 59200
rect 279896 54534 279924 59191
rect 279884 54528 279936 54534
rect 279884 54470 279936 54476
rect 280080 53106 280108 59599
rect 281092 59401 281120 59735
rect 292762 59800 292818 59809
rect 289818 59735 289820 59744
rect 287704 59706 287756 59712
rect 289872 59735 289874 59744
rect 290464 59764 290516 59770
rect 289820 59706 289872 59712
rect 292762 59735 292764 59744
rect 290464 59706 290516 59712
rect 292816 59735 292818 59744
rect 304998 59800 305054 59809
rect 304998 59735 305054 59744
rect 308954 59800 309010 59809
rect 308954 59735 309010 59744
rect 311990 59800 312046 59809
rect 311990 59735 312046 59744
rect 315762 59800 315818 59809
rect 319626 59800 319682 59809
rect 315762 59735 315764 59744
rect 292764 59706 292816 59712
rect 282826 59664 282882 59673
rect 286874 59664 286930 59673
rect 282826 59599 282882 59608
rect 284944 59628 284996 59634
rect 281446 59528 281502 59537
rect 281446 59463 281502 59472
rect 281078 59392 281134 59401
rect 281078 59327 281134 59336
rect 280068 53100 280120 53106
rect 280068 53042 280120 53048
rect 281460 32434 281488 59463
rect 281540 56092 281592 56098
rect 281540 56034 281592 56040
rect 281448 32428 281500 32434
rect 281448 32370 281500 32376
rect 278780 31272 278832 31278
rect 278780 31214 278832 31220
rect 277400 31068 277452 31074
rect 277400 31010 277452 31016
rect 278688 31068 278740 31074
rect 278688 31010 278740 31016
rect 277032 29708 277084 29714
rect 277032 29650 277084 29656
rect 277412 16574 277440 31010
rect 278792 16574 278820 31214
rect 277412 16546 278360 16574
rect 278792 16546 279096 16574
rect 276664 16380 276716 16386
rect 276664 16322 276716 16328
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276676 354 276704 16322
rect 278332 480 278360 16546
rect 277094 354 277206 480
rect 276676 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280712 16448 280764 16454
rect 280712 16390 280764 16396
rect 280724 480 280752 16390
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281552 354 281580 56034
rect 282840 33794 282868 59599
rect 286874 59599 286876 59608
rect 284944 59570 284996 59576
rect 286928 59599 286930 59608
rect 286876 59570 286928 59576
rect 284114 59528 284170 59537
rect 284114 59463 284170 59472
rect 283930 59392 283986 59401
rect 283930 59327 283986 59336
rect 283944 50386 283972 59327
rect 284128 51746 284156 59463
rect 284300 51944 284352 51950
rect 284300 51886 284352 51892
rect 284116 51740 284168 51746
rect 284116 51682 284168 51688
rect 283932 50380 283984 50386
rect 283932 50322 283984 50328
rect 282920 43648 282972 43654
rect 282920 43590 282972 43596
rect 282828 33788 282880 33794
rect 282828 33730 282880 33736
rect 282932 16574 282960 43590
rect 282932 16546 283144 16574
rect 283116 480 283144 16546
rect 284312 3738 284340 51886
rect 284956 28422 284984 59570
rect 286874 59528 286930 59537
rect 286336 59486 286874 59514
rect 284944 28416 284996 28422
rect 284944 28358 284996 28364
rect 284392 16516 284444 16522
rect 284392 16458 284444 16464
rect 284300 3732 284352 3738
rect 284300 3674 284352 3680
rect 284404 3482 284432 16458
rect 286336 10334 286364 59486
rect 286874 59463 286930 59472
rect 286874 59392 286930 59401
rect 286874 59327 286930 59336
rect 286888 45554 286916 59327
rect 286520 45526 286916 45554
rect 286520 11762 286548 45526
rect 287716 25770 287744 59706
rect 289082 59256 289138 59265
rect 289082 59191 289138 59200
rect 289096 31210 289124 59191
rect 290476 45014 290504 59706
rect 296626 59664 296682 59673
rect 295248 59628 295300 59634
rect 296626 59599 296628 59608
rect 295248 59570 295300 59576
rect 296680 59599 296682 59608
rect 303618 59664 303674 59673
rect 303618 59599 303674 59608
rect 296628 59570 296680 59576
rect 290646 59528 290702 59537
rect 290646 59463 290702 59472
rect 293222 59528 293278 59537
rect 293222 59463 293278 59472
rect 290660 46374 290688 59463
rect 291842 59392 291898 59401
rect 291842 59327 291898 59336
rect 290648 46368 290700 46374
rect 290648 46310 290700 46316
rect 290464 45008 290516 45014
rect 290464 44950 290516 44956
rect 289084 31204 289136 31210
rect 289084 31146 289136 31152
rect 287704 25764 287756 25770
rect 287704 25706 287756 25712
rect 287060 21548 287112 21554
rect 287060 21490 287112 21496
rect 287072 16574 287100 21490
rect 287072 16546 287376 16574
rect 286508 11756 286560 11762
rect 286508 11698 286560 11704
rect 286324 10328 286376 10334
rect 286324 10270 286376 10276
rect 286600 6656 286652 6662
rect 286600 6598 286652 6604
rect 285036 3732 285088 3738
rect 285036 3674 285088 3680
rect 284312 3454 284432 3482
rect 284312 480 284340 3454
rect 281878 354 281990 480
rect 281552 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285048 354 285076 3674
rect 286612 480 286640 6598
rect 285374 354 285486 480
rect 285048 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 291856 13326 291884 59327
rect 293236 13394 293264 59463
rect 293406 59392 293462 59401
rect 293406 59327 293462 59336
rect 293420 13462 293448 59327
rect 295260 57390 295288 59570
rect 296626 59528 296682 59537
rect 295996 59486 296626 59514
rect 295248 57384 295300 57390
rect 295248 57326 295300 57332
rect 295340 49224 295392 49230
rect 295340 49166 295392 49172
rect 295352 16574 295380 49166
rect 295352 16546 295656 16574
rect 293408 13456 293460 13462
rect 293408 13398 293460 13404
rect 293224 13388 293276 13394
rect 293224 13330 293276 13336
rect 291844 13320 291896 13326
rect 291844 13262 291896 13268
rect 294880 13320 294932 13326
rect 294880 13262 294932 13268
rect 291384 13252 291436 13258
rect 291384 13194 291436 13200
rect 288992 6588 289044 6594
rect 288992 6530 289044 6536
rect 290188 6588 290240 6594
rect 290188 6530 290240 6536
rect 289004 480 289032 6530
rect 290200 480 290228 6530
rect 291396 480 291424 13194
rect 292580 6520 292632 6526
rect 292580 6462 292632 6468
rect 293684 6520 293736 6526
rect 293684 6462 293736 6468
rect 292592 480 292620 6462
rect 293696 480 293724 6462
rect 294892 480 294920 13262
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 295628 354 295656 16546
rect 295996 10402 296024 59486
rect 296626 59463 296682 59472
rect 302238 59528 302294 59537
rect 302238 59463 302294 59472
rect 296166 59256 296222 59265
rect 296166 59191 296222 59200
rect 296180 10538 296208 59191
rect 299480 47796 299532 47802
rect 299480 47738 299532 47744
rect 299492 16574 299520 47738
rect 299492 16546 299704 16574
rect 298100 13388 298152 13394
rect 298100 13330 298152 13336
rect 296168 10532 296220 10538
rect 296168 10474 296220 10480
rect 295984 10396 296036 10402
rect 295984 10338 296036 10344
rect 297272 10328 297324 10334
rect 297272 10270 297324 10276
rect 297284 480 297312 10270
rect 296046 354 296158 480
rect 295628 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298112 354 298140 13330
rect 299676 480 299704 16546
rect 301504 13456 301556 13462
rect 301504 13398 301556 13404
rect 300768 6724 300820 6730
rect 300768 6666 300820 6672
rect 300780 480 300808 6666
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 13398
rect 302252 10470 302280 59463
rect 303632 32638 303660 59599
rect 305012 58818 305040 59735
rect 306378 59392 306434 59401
rect 306378 59327 306434 59336
rect 307942 59392 307998 59401
rect 307942 59327 307998 59336
rect 305274 59256 305330 59265
rect 305274 59191 305330 59200
rect 305090 59120 305146 59129
rect 305090 59055 305146 59064
rect 305000 58812 305052 58818
rect 305000 58754 305052 58760
rect 303620 32632 303672 32638
rect 303620 32574 303672 32580
rect 305104 10606 305132 59055
rect 305288 10674 305316 59191
rect 306392 10742 306420 59327
rect 307956 53310 307984 59327
rect 308968 56030 308996 59735
rect 309138 59528 309194 59537
rect 309138 59463 309194 59472
rect 308956 56024 309008 56030
rect 308956 55966 309008 55972
rect 307944 53304 307996 53310
rect 307944 53246 307996 53252
rect 309152 33998 309180 59463
rect 310518 59392 310574 59401
rect 310518 59327 310574 59336
rect 311898 59392 311954 59401
rect 311898 59327 311954 59336
rect 310532 51882 310560 59327
rect 311912 54738 311940 59327
rect 312004 57458 312032 59735
rect 315816 59735 315818 59744
rect 317604 59764 317656 59770
rect 315764 59706 315816 59712
rect 319626 59735 319682 59744
rect 322570 59800 322626 59809
rect 326158 59800 326214 59809
rect 322570 59735 322572 59744
rect 317604 59706 317656 59712
rect 314842 59528 314898 59537
rect 314842 59463 314898 59472
rect 317418 59528 317474 59537
rect 317418 59463 317474 59472
rect 313278 59392 313334 59401
rect 313278 59327 313334 59336
rect 311992 57452 312044 57458
rect 311992 57394 312044 57400
rect 311900 54732 311952 54738
rect 311900 54674 311952 54680
rect 310520 51876 310572 51882
rect 310520 51818 310572 51824
rect 311164 51876 311216 51882
rect 311164 51818 311216 51824
rect 309140 33992 309192 33998
rect 309140 33934 309192 33940
rect 307024 22908 307076 22914
rect 307024 22850 307076 22856
rect 306380 10736 306432 10742
rect 306380 10678 306432 10684
rect 305276 10668 305328 10674
rect 305276 10610 305328 10616
rect 305092 10600 305144 10606
rect 305092 10542 305144 10548
rect 302240 10464 302292 10470
rect 302240 10406 302292 10412
rect 303160 6452 303212 6458
rect 303160 6394 303212 6400
rect 304356 6452 304408 6458
rect 304356 6394 304408 6400
rect 303172 480 303200 6394
rect 304368 480 304396 6394
rect 306748 6384 306800 6390
rect 306748 6326 306800 6332
rect 305552 3256 305604 3262
rect 305552 3198 305604 3204
rect 305564 480 305592 3198
rect 306760 480 306788 6326
rect 307036 3262 307064 22850
rect 307944 10396 307996 10402
rect 307944 10338 307996 10344
rect 307024 3256 307076 3262
rect 307024 3198 307076 3204
rect 307956 480 307984 10338
rect 310244 6316 310296 6322
rect 310244 6258 310296 6264
rect 309048 3052 309100 3058
rect 309048 2994 309100 3000
rect 309060 480 309088 2994
rect 310256 480 310284 6258
rect 311176 3058 311204 51818
rect 311900 50448 311952 50454
rect 311900 50390 311952 50396
rect 311912 16574 311940 50390
rect 313292 17406 313320 59327
rect 314856 50590 314884 59463
rect 316130 59392 316186 59401
rect 316130 59327 316186 59336
rect 316040 56024 316092 56030
rect 316040 55966 316092 55972
rect 314844 50584 314896 50590
rect 314844 50526 314896 50532
rect 314660 38140 314712 38146
rect 314660 38082 314712 38088
rect 313280 17400 313332 17406
rect 313280 17342 313332 17348
rect 311912 16546 312216 16574
rect 311440 6316 311492 6322
rect 311440 6258 311492 6264
rect 311164 3052 311216 3058
rect 311164 2994 311216 3000
rect 311452 480 311480 6258
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 354 312216 16546
rect 313832 6248 313884 6254
rect 313832 6190 313884 6196
rect 313844 480 313872 6190
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314672 354 314700 38082
rect 316052 16574 316080 55966
rect 316144 20126 316172 59327
rect 316132 20120 316184 20126
rect 316132 20062 316184 20068
rect 317432 18766 317460 59463
rect 317616 21622 317644 59706
rect 318798 59664 318854 59673
rect 318798 59599 318854 59608
rect 317604 21616 317656 21622
rect 317604 21558 317656 21564
rect 317420 18760 317472 18766
rect 317420 18702 317472 18708
rect 316052 16546 316264 16574
rect 316236 480 316264 16546
rect 318812 11830 318840 59599
rect 319640 58818 319668 59735
rect 322624 59735 322626 59744
rect 324688 59764 324740 59770
rect 322572 59706 322624 59712
rect 326158 59735 326214 59744
rect 334346 59800 334402 59809
rect 339130 59800 339186 59809
rect 335280 59770 335492 59786
rect 334346 59735 334348 59744
rect 324688 59706 324740 59712
rect 320454 59664 320510 59673
rect 320454 59599 320510 59608
rect 324502 59664 324558 59673
rect 324502 59599 324504 59608
rect 320270 59528 320326 59537
rect 320270 59463 320326 59472
rect 319628 58812 319680 58818
rect 319628 58754 319680 58760
rect 320180 43580 320232 43586
rect 320180 43522 320232 43528
rect 320192 16574 320220 43522
rect 320284 22982 320312 59463
rect 320468 58546 320496 59599
rect 324556 59599 324558 59608
rect 324504 59570 324556 59576
rect 324502 59528 324558 59537
rect 324502 59463 324558 59472
rect 322938 59392 322994 59401
rect 322938 59327 322994 59336
rect 321744 58812 321796 58818
rect 321744 58754 321796 58760
rect 320456 58540 320508 58546
rect 320456 58482 320508 58488
rect 321560 57384 321612 57390
rect 321560 57326 321612 57332
rect 320824 24268 320876 24274
rect 320824 24210 320876 24216
rect 320272 22976 320324 22982
rect 320272 22918 320324 22924
rect 320192 16546 320496 16574
rect 318800 11824 318852 11830
rect 318800 11766 318852 11772
rect 317328 6180 317380 6186
rect 317328 6122 317380 6128
rect 318524 6180 318576 6186
rect 318524 6122 318576 6128
rect 317340 480 317368 6122
rect 318536 480 318564 6122
rect 319720 3324 319772 3330
rect 319720 3266 319772 3272
rect 319732 480 319760 3266
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 320836 3330 320864 24210
rect 321572 6914 321600 57326
rect 321756 11898 321784 58754
rect 321928 58540 321980 58546
rect 321928 58482 321980 58488
rect 321744 11892 321796 11898
rect 321744 11834 321796 11840
rect 321940 7750 321968 58482
rect 322952 24342 322980 59327
rect 324320 35352 324372 35358
rect 324320 35294 324372 35300
rect 322940 24336 322992 24342
rect 322940 24278 322992 24284
rect 322940 11756 322992 11762
rect 322940 11698 322992 11704
rect 321928 7744 321980 7750
rect 321928 7686 321980 7692
rect 321572 6886 322152 6914
rect 320824 3324 320876 3330
rect 320824 3266 320876 3272
rect 322124 480 322152 6886
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 322952 354 322980 11698
rect 324332 3210 324360 35294
rect 324516 12034 324544 59463
rect 324504 12028 324556 12034
rect 324504 11970 324556 11976
rect 324700 11966 324728 59706
rect 325700 59628 325752 59634
rect 325700 59570 325752 59576
rect 325712 12102 325740 59570
rect 326172 58886 326200 59735
rect 334400 59735 334402 59744
rect 335268 59764 335492 59770
rect 334348 59706 334400 59712
rect 335320 59758 335492 59764
rect 335268 59706 335320 59712
rect 327262 59664 327318 59673
rect 327262 59599 327318 59608
rect 334162 59664 334218 59673
rect 334162 59599 334218 59608
rect 327078 59392 327134 59401
rect 327078 59327 327134 59336
rect 326160 58880 326212 58886
rect 326160 58822 326212 58828
rect 327092 52018 327120 59327
rect 327080 52012 327132 52018
rect 327080 51954 327132 51960
rect 327080 36712 327132 36718
rect 327080 36654 327132 36660
rect 327092 16574 327120 36654
rect 327276 27062 327304 59599
rect 328550 59528 328606 59537
rect 328550 59463 328606 59472
rect 331402 59528 331458 59537
rect 331402 59463 331458 59472
rect 328564 56166 328592 59463
rect 329930 59392 329986 59401
rect 329930 59327 329986 59336
rect 328552 56160 328604 56166
rect 328552 56102 328604 56108
rect 329840 40860 329892 40866
rect 329840 40802 329892 40808
rect 329104 39500 329156 39506
rect 329104 39442 329156 39448
rect 327264 27056 327316 27062
rect 327264 26998 327316 27004
rect 327092 16546 328040 16574
rect 325700 12096 325752 12102
rect 325700 12038 325752 12044
rect 324688 11960 324740 11966
rect 324688 11902 324740 11908
rect 324412 11824 324464 11830
rect 324412 11766 324464 11772
rect 324424 3398 324452 11766
rect 324412 3392 324464 3398
rect 324412 3334 324464 3340
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 324332 3182 324452 3210
rect 324424 480 324452 3182
rect 325620 480 325648 3334
rect 326804 2916 326856 2922
rect 326804 2858 326856 2864
rect 326816 480 326844 2858
rect 328012 480 328040 16546
rect 329116 2922 329144 39442
rect 329852 16574 329880 40802
rect 329944 29850 329972 59327
rect 331220 38072 331272 38078
rect 331220 38014 331272 38020
rect 329932 29844 329984 29850
rect 329932 29786 329984 29792
rect 329852 16546 330432 16574
rect 329196 7744 329248 7750
rect 329196 7686 329248 7692
rect 329104 2916 329156 2922
rect 329104 2858 329156 2864
rect 329208 480 329236 7686
rect 330404 480 330432 16546
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331232 354 331260 38014
rect 331416 31278 331444 59463
rect 332598 59392 332654 59401
rect 332598 59327 332654 59336
rect 332612 43654 332640 59327
rect 332600 43648 332652 43654
rect 332600 43590 332652 43596
rect 333980 39568 334032 39574
rect 333980 39510 334032 39516
rect 331404 31272 331456 31278
rect 331404 31214 331456 31220
rect 332600 27056 332652 27062
rect 332600 26998 332652 27004
rect 332612 3398 332640 26998
rect 333992 16574 334020 39510
rect 333992 16546 334112 16574
rect 332692 10464 332744 10470
rect 332692 10406 332744 10412
rect 332600 3392 332652 3398
rect 332600 3334 332652 3340
rect 332704 480 332732 10406
rect 333888 3392 333940 3398
rect 333888 3334 333940 3340
rect 333900 480 333928 3334
rect 334084 490 334112 16546
rect 334176 6594 334204 59599
rect 334254 59392 334310 59401
rect 334254 59327 334310 59336
rect 334268 55214 334296 59327
rect 335360 58812 335412 58818
rect 335360 58754 335412 58760
rect 334268 55186 334388 55214
rect 334360 6662 334388 55186
rect 334348 6656 334400 6662
rect 334348 6598 334400 6604
rect 334164 6588 334216 6594
rect 334164 6530 334216 6536
rect 335372 3482 335400 58754
rect 335464 6526 335492 59758
rect 339130 59735 339132 59744
rect 339184 59735 339186 59744
rect 340878 59800 340934 59809
rect 345386 59800 345442 59809
rect 340878 59735 340934 59744
rect 340972 59764 341024 59770
rect 339132 59706 339184 59712
rect 338302 59528 338358 59537
rect 338302 59463 338358 59472
rect 336738 59256 336794 59265
rect 336738 59191 336794 59200
rect 336752 10334 336780 59191
rect 338120 40928 338172 40934
rect 338120 40870 338172 40876
rect 338132 16574 338160 40870
rect 338132 16546 338252 16574
rect 336740 10328 336792 10334
rect 336740 10270 336792 10276
rect 335452 6520 335504 6526
rect 335452 6462 335504 6468
rect 338224 3482 338252 16546
rect 338316 6458 338344 59463
rect 338486 59392 338542 59401
rect 338486 59327 338542 59336
rect 339498 59392 339554 59401
rect 339498 59327 339554 59336
rect 338500 6730 338528 59327
rect 339512 10402 339540 59327
rect 340892 57390 340920 59735
rect 345386 59735 345442 59744
rect 347686 59800 347742 59809
rect 347686 59735 347742 59744
rect 355598 59800 355654 59809
rect 360382 59800 360438 59809
rect 355598 59735 355600 59744
rect 340972 59706 341024 59712
rect 340880 57384 340932 57390
rect 340880 57326 340932 57332
rect 340880 42288 340932 42294
rect 340880 42230 340932 42236
rect 340144 42220 340196 42226
rect 340144 42162 340196 42168
rect 339592 10532 339644 10538
rect 339592 10474 339644 10480
rect 339500 10396 339552 10402
rect 339500 10338 339552 10344
rect 338488 6724 338540 6730
rect 338488 6666 338540 6672
rect 338304 6452 338356 6458
rect 338304 6394 338356 6400
rect 335372 3454 336320 3482
rect 338224 3454 338712 3482
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334084 462 334664 490
rect 336292 480 336320 3454
rect 337476 3392 337528 3398
rect 337476 3334 337528 3340
rect 337488 480 337516 3334
rect 338684 480 338712 3454
rect 334636 354 334664 462
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339604 354 339632 10474
rect 340156 3398 340184 42162
rect 340892 3398 340920 42230
rect 340984 6322 341012 59706
rect 341154 59528 341210 59537
rect 341154 59463 341210 59472
rect 341168 38146 341196 59463
rect 345018 59392 345074 59401
rect 345018 59327 345074 59336
rect 342258 59256 342314 59265
rect 342258 59191 342314 59200
rect 343822 59256 343878 59265
rect 343822 59191 343878 59200
rect 341156 38140 341208 38146
rect 341156 38082 341208 38088
rect 340972 6316 341024 6322
rect 340972 6258 341024 6264
rect 342272 6186 342300 59191
rect 342904 45008 342956 45014
rect 342904 44950 342956 44956
rect 342260 6180 342312 6186
rect 342260 6122 342312 6128
rect 340144 3392 340196 3398
rect 340144 3334 340196 3340
rect 340880 3392 340932 3398
rect 340880 3334 340932 3340
rect 342168 3392 342220 3398
rect 342168 3334 342220 3340
rect 340972 3324 341024 3330
rect 340972 3266 341024 3272
rect 340984 480 341012 3266
rect 342180 480 342208 3334
rect 342916 3330 342944 44950
rect 343836 11830 343864 59191
rect 345032 55214 345060 59327
rect 345400 58818 345428 59735
rect 346490 59528 346546 59537
rect 346490 59463 346546 59472
rect 346400 59356 346452 59362
rect 346400 59298 346452 59304
rect 345388 58812 345440 58818
rect 345388 58754 345440 58760
rect 345032 55186 345152 55214
rect 345020 45076 345072 45082
rect 345020 45018 345072 45024
rect 343824 11824 343876 11830
rect 343824 11766 343876 11772
rect 345032 6914 345060 45018
rect 345124 7750 345152 55186
rect 345664 35352 345716 35358
rect 345664 35294 345716 35300
rect 345112 7744 345164 7750
rect 345112 7686 345164 7692
rect 345032 6886 345336 6914
rect 343364 6316 343416 6322
rect 343364 6258 343416 6264
rect 342904 3324 342956 3330
rect 342904 3266 342956 3272
rect 343376 480 343404 6258
rect 344560 4140 344612 4146
rect 344560 4082 344612 4088
rect 344572 480 344600 4082
rect 339838 354 339950 480
rect 339604 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345308 354 345336 6886
rect 345676 4146 345704 35294
rect 346412 6914 346440 59298
rect 346504 10470 346532 59463
rect 347700 59401 347728 59735
rect 355652 59735 355654 59744
rect 358268 59764 358320 59770
rect 355600 59706 355652 59712
rect 360382 59735 360438 59744
rect 361486 59800 361542 59809
rect 361486 59735 361542 59744
rect 365350 59800 365406 59809
rect 369306 59800 369362 59809
rect 365350 59735 365352 59744
rect 358268 59706 358320 59712
rect 347870 59664 347926 59673
rect 347870 59599 347926 59608
rect 357622 59664 357678 59673
rect 357622 59599 357678 59608
rect 347778 59528 347834 59537
rect 347778 59463 347834 59472
rect 347686 59392 347742 59401
rect 347792 59362 347820 59463
rect 347686 59327 347742 59336
rect 347780 59356 347832 59362
rect 347780 59298 347832 59304
rect 347884 55214 347912 59599
rect 349158 59528 349214 59537
rect 349158 59463 349214 59472
rect 352746 59528 352802 59537
rect 355322 59528 355378 59537
rect 352746 59463 352748 59472
rect 347884 55186 348004 55214
rect 347780 17400 347832 17406
rect 347780 17342 347832 17348
rect 346492 10464 346544 10470
rect 346492 10406 346544 10412
rect 347792 6914 347820 17342
rect 347976 10538 348004 55186
rect 347964 10532 348016 10538
rect 347964 10474 348016 10480
rect 346412 6886 346992 6914
rect 347792 6886 348096 6914
rect 345664 4140 345716 4146
rect 345664 4082 345716 4088
rect 346964 480 346992 6886
rect 348068 480 348096 6886
rect 349172 3398 349200 59463
rect 352800 59463 352802 59472
rect 354680 59492 354732 59498
rect 352748 59434 352800 59440
rect 355322 59463 355378 59472
rect 354680 59434 354732 59440
rect 349342 59392 349398 59401
rect 349342 59327 349398 59336
rect 353942 59392 353998 59401
rect 353942 59327 353998 59336
rect 349252 46436 349304 46442
rect 349252 46378 349304 46384
rect 349160 3392 349212 3398
rect 349160 3334 349212 3340
rect 349264 480 349292 46378
rect 349356 6322 349384 59327
rect 352562 59256 352618 59265
rect 352562 59191 352618 59200
rect 351920 33924 351972 33930
rect 351920 33866 351972 33872
rect 351932 16574 351960 33866
rect 351932 16546 352512 16574
rect 349344 6316 349396 6322
rect 349344 6258 349396 6264
rect 352484 3482 352512 16546
rect 352576 5574 352604 59191
rect 353956 16574 353984 59327
rect 354692 58002 354720 59434
rect 354680 57996 354732 58002
rect 354680 57938 354732 57944
rect 354036 36712 354088 36718
rect 354036 36654 354088 36660
rect 353864 16546 353984 16574
rect 353864 6186 353892 16546
rect 354048 6914 354076 36654
rect 355336 10334 355364 59463
rect 357636 59401 357664 59599
rect 358082 59528 358138 59537
rect 358082 59463 358138 59472
rect 356702 59392 356758 59401
rect 356702 59327 356758 59336
rect 357622 59392 357678 59401
rect 357622 59327 357678 59336
rect 356060 49156 356112 49162
rect 356060 49098 356112 49104
rect 356072 16574 356100 49098
rect 356072 16546 356376 16574
rect 355324 10328 355376 10334
rect 355324 10270 355376 10276
rect 353956 6886 354076 6914
rect 353852 6180 353904 6186
rect 353852 6122 353904 6128
rect 352564 5568 352616 5574
rect 352564 5510 352616 5516
rect 352484 3454 352880 3482
rect 350448 3392 350500 3398
rect 350448 3334 350500 3340
rect 351644 3392 351696 3398
rect 351644 3334 351696 3340
rect 350460 480 350488 3334
rect 351656 480 351684 3334
rect 352852 480 352880 3454
rect 353956 3398 353984 6886
rect 354036 5568 354088 5574
rect 354036 5510 354088 5516
rect 353944 3392 353996 3398
rect 353944 3334 353996 3340
rect 354048 480 354076 5510
rect 355232 3392 355284 3398
rect 355232 3334 355284 3340
rect 355244 480 355272 3334
rect 356348 480 356376 16546
rect 356716 6730 356744 59327
rect 356796 31204 356848 31210
rect 356796 31146 356848 31152
rect 356704 6724 356756 6730
rect 356704 6666 356756 6672
rect 356808 3398 356836 31146
rect 357440 11824 357492 11830
rect 357440 11766 357492 11772
rect 357452 3398 357480 11766
rect 358096 6594 358124 59463
rect 358280 6662 358308 59706
rect 360396 59401 360424 59735
rect 360474 59528 360530 59537
rect 360474 59463 360530 59472
rect 361026 59528 361082 59537
rect 361026 59463 361082 59472
rect 359462 59392 359518 59401
rect 359462 59327 359518 59336
rect 360382 59392 360438 59401
rect 360382 59327 360438 59336
rect 358820 32564 358872 32570
rect 358820 32506 358872 32512
rect 358832 6914 358860 32506
rect 359476 16574 359504 59327
rect 360200 57996 360252 58002
rect 360200 57938 360252 57944
rect 360212 16574 360240 57938
rect 360488 51074 360516 59463
rect 360488 51046 360884 51074
rect 359476 16546 359596 16574
rect 360212 16546 360792 16574
rect 358832 6886 359504 6914
rect 358268 6656 358320 6662
rect 358268 6598 358320 6604
rect 358084 6588 358136 6594
rect 358084 6530 358136 6536
rect 357532 6180 357584 6186
rect 357532 6122 357584 6128
rect 356796 3392 356848 3398
rect 356796 3334 356848 3340
rect 357440 3392 357492 3398
rect 357440 3334 357492 3340
rect 357544 480 357572 6122
rect 358728 3392 358780 3398
rect 358728 3334 358780 3340
rect 358740 480 358768 3334
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 6886
rect 359568 6526 359596 16546
rect 359556 6520 359608 6526
rect 359556 6462 359608 6468
rect 360764 3482 360792 16546
rect 360856 6458 360884 51046
rect 360844 6452 360896 6458
rect 360844 6394 360896 6400
rect 361040 6390 361068 59463
rect 361500 59401 361528 59735
rect 365404 59735 365406 59744
rect 367744 59764 367796 59770
rect 365352 59706 365404 59712
rect 378046 59800 378102 59809
rect 369306 59735 369308 59744
rect 367744 59706 367796 59712
rect 369360 59735 369362 59744
rect 371976 59764 372028 59770
rect 369308 59706 369360 59712
rect 381910 59800 381912 59809
rect 383292 59832 383344 59838
rect 381964 59800 381966 59809
rect 378102 59758 378456 59786
rect 378046 59735 378102 59744
rect 371976 59706 372028 59712
rect 363326 59664 363382 59673
rect 363382 59622 363828 59650
rect 363326 59599 363382 59608
rect 362222 59528 362278 59537
rect 362222 59463 362278 59472
rect 361486 59392 361542 59401
rect 361486 59327 361542 59336
rect 361028 6384 361080 6390
rect 361028 6326 361080 6332
rect 362236 6322 362264 59463
rect 363800 59401 363828 59622
rect 365166 59528 365222 59537
rect 365166 59463 365222 59472
rect 363602 59392 363658 59401
rect 363602 59327 363658 59336
rect 363786 59392 363842 59401
rect 363786 59327 363842 59336
rect 364982 59392 365038 59401
rect 364982 59327 365038 59336
rect 362960 47728 363012 47734
rect 362960 47670 363012 47676
rect 362972 16574 363000 47670
rect 362972 16546 363552 16574
rect 362224 6316 362276 6322
rect 362224 6258 362276 6264
rect 360764 3454 361160 3482
rect 361132 480 361160 3454
rect 362316 3392 362368 3398
rect 362316 3334 362368 3340
rect 362328 480 362356 3334
rect 363524 480 363552 16546
rect 363616 6254 363644 59327
rect 363696 18828 363748 18834
rect 363696 18770 363748 18776
rect 363604 6248 363656 6254
rect 363604 6190 363656 6196
rect 363708 3398 363736 18770
rect 364616 10328 364668 10334
rect 364616 10270 364668 10276
rect 363696 3392 363748 3398
rect 363696 3334 363748 3340
rect 364628 480 364656 10270
rect 364996 6186 365024 59327
rect 365180 7954 365208 59463
rect 366362 59256 366418 59265
rect 366362 59191 366418 59200
rect 365720 28484 365772 28490
rect 365720 28426 365772 28432
rect 365168 7948 365220 7954
rect 365168 7890 365220 7896
rect 364984 6180 365036 6186
rect 364984 6122 365036 6128
rect 365732 3398 365760 28426
rect 366376 7886 366404 59191
rect 366364 7880 366416 7886
rect 366364 7822 366416 7828
rect 367756 7818 367784 59706
rect 369122 59528 369178 59537
rect 369122 59463 369178 59472
rect 371146 59528 371202 59537
rect 371146 59463 371202 59472
rect 367926 59256 367982 59265
rect 367926 59191 367982 59200
rect 367744 7812 367796 7818
rect 367744 7754 367796 7760
rect 367940 7750 367968 59191
rect 369136 8294 369164 59463
rect 370502 59256 370558 59265
rect 370502 59191 370558 59200
rect 369860 50516 369912 50522
rect 369860 50458 369912 50464
rect 369872 16574 369900 50458
rect 369872 16546 370176 16574
rect 369124 8288 369176 8294
rect 369124 8230 369176 8236
rect 367928 7744 367980 7750
rect 367928 7686 367980 7692
rect 368204 6724 368256 6730
rect 368204 6666 368256 6672
rect 365812 3732 365864 3738
rect 365812 3674 365864 3680
rect 365720 3392 365772 3398
rect 365720 3334 365772 3340
rect 365824 480 365852 3674
rect 367008 3392 367060 3398
rect 367008 3334 367060 3340
rect 367020 480 367048 3334
rect 368216 480 368244 6666
rect 369400 3392 369452 3398
rect 369400 3334 369452 3340
rect 369412 480 369440 3334
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370148 354 370176 16546
rect 370516 8226 370544 59191
rect 371160 58886 371188 59463
rect 371148 58880 371200 58886
rect 371148 58822 371200 58828
rect 371884 49224 371936 49230
rect 371884 49166 371936 49172
rect 370596 46436 370648 46442
rect 370596 46378 370648 46384
rect 370504 8220 370556 8226
rect 370504 8162 370556 8168
rect 370608 3398 370636 46378
rect 371700 6656 371752 6662
rect 371700 6598 371752 6604
rect 370596 3392 370648 3398
rect 370596 3334 370648 3340
rect 371712 480 371740 6598
rect 371896 3738 371924 49166
rect 371988 28490 372016 59706
rect 374090 59664 374146 59673
rect 374090 59599 374092 59608
rect 374144 59599 374146 59608
rect 376024 59628 376076 59634
rect 374092 59570 374144 59576
rect 376024 59570 376076 59576
rect 374090 59528 374146 59537
rect 374146 59486 374224 59514
rect 374090 59463 374146 59472
rect 374090 59392 374146 59401
rect 374196 59378 374224 59486
rect 374196 59350 374776 59378
rect 374090 59327 374146 59336
rect 372158 59256 372214 59265
rect 372158 59191 372214 59200
rect 372172 32638 372200 59191
rect 374104 55214 374132 59327
rect 374748 55214 374776 59350
rect 374104 55186 374684 55214
rect 374748 55186 374868 55214
rect 372160 32632 372212 32638
rect 372160 32574 372212 32580
rect 371976 28484 372028 28490
rect 371976 28426 372028 28432
rect 374656 10810 374684 55186
rect 374644 10804 374696 10810
rect 374644 10746 374696 10752
rect 374840 10742 374868 55186
rect 374828 10736 374880 10742
rect 374828 10678 374880 10684
rect 376036 10674 376064 59570
rect 378428 59537 378456 59758
rect 381910 59735 381966 59744
rect 383290 59800 383292 59809
rect 383344 59800 383346 59809
rect 383290 59735 383346 59744
rect 383842 59800 383898 59809
rect 384854 59800 384910 59809
rect 383898 59758 383976 59786
rect 383842 59735 383898 59744
rect 377586 59528 377642 59537
rect 377586 59463 377642 59472
rect 378414 59528 378470 59537
rect 378414 59463 378470 59472
rect 381542 59528 381598 59537
rect 381542 59463 381598 59472
rect 383842 59528 383898 59537
rect 383842 59463 383898 59472
rect 377402 59392 377458 59401
rect 377402 59327 377458 59336
rect 376760 43512 376812 43518
rect 376760 43454 376812 43460
rect 376116 28416 376168 28422
rect 376116 28358 376168 28364
rect 376024 10668 376076 10674
rect 376024 10610 376076 10616
rect 374092 7676 374144 7682
rect 374092 7618 374144 7624
rect 372896 4004 372948 4010
rect 372896 3946 372948 3952
rect 371884 3732 371936 3738
rect 371884 3674 371936 3680
rect 372908 480 372936 3946
rect 374104 480 374132 7618
rect 375288 6588 375340 6594
rect 375288 6530 375340 6536
rect 375300 480 375328 6530
rect 376128 4010 376156 28358
rect 376772 6914 376800 43454
rect 377416 10606 377444 59327
rect 377404 10600 377456 10606
rect 377404 10542 377456 10548
rect 377600 10538 377628 59463
rect 380162 59392 380218 59401
rect 380162 59327 380218 59336
rect 378598 59256 378654 59265
rect 378598 59191 378654 59200
rect 378612 55214 378640 59191
rect 378612 55186 378824 55214
rect 377588 10532 377640 10538
rect 377588 10474 377640 10480
rect 378796 10470 378824 55186
rect 380176 43654 380204 59327
rect 380164 43648 380216 43654
rect 380164 43590 380216 43596
rect 380900 35284 380952 35290
rect 380900 35226 380952 35232
rect 378876 32564 378928 32570
rect 378876 32506 378928 32512
rect 378784 10464 378836 10470
rect 378784 10406 378836 10412
rect 378888 6914 378916 32506
rect 380912 16574 380940 35226
rect 380912 16546 381216 16574
rect 376772 6886 377720 6914
rect 376116 4004 376168 4010
rect 376116 3946 376168 3952
rect 376484 3392 376536 3398
rect 376484 3334 376536 3340
rect 376496 480 376524 3334
rect 377692 480 377720 6886
rect 378796 6886 378916 6914
rect 378796 3398 378824 6886
rect 378876 6520 378928 6526
rect 378876 6462 378928 6468
rect 378784 3392 378836 3398
rect 378784 3334 378836 3340
rect 378888 480 378916 6462
rect 379980 3392 380032 3398
rect 379980 3334 380032 3340
rect 379992 480 380020 3334
rect 381188 480 381216 16546
rect 381556 10334 381584 59463
rect 381726 59392 381782 59401
rect 381726 59327 381782 59336
rect 383014 59392 383070 59401
rect 383014 59327 383070 59336
rect 381740 10402 381768 59327
rect 382924 43512 382976 43518
rect 382924 43454 382976 43460
rect 381728 10396 381780 10402
rect 381728 10338 381780 10344
rect 381544 10328 381596 10334
rect 381544 10270 381596 10276
rect 382372 6452 382424 6458
rect 382372 6394 382424 6400
rect 382384 480 382412 6394
rect 382936 3398 382964 43454
rect 383028 33998 383056 59327
rect 383856 57390 383884 59463
rect 383844 57384 383896 57390
rect 383844 57326 383896 57332
rect 383948 50522 383976 59758
rect 384854 59735 384910 59744
rect 385958 59800 386014 59809
rect 388718 59800 388774 59809
rect 385958 59735 385960 59744
rect 384868 59401 384896 59735
rect 386012 59735 386014 59744
rect 388628 59764 388680 59770
rect 385960 59706 386012 59712
rect 391662 59800 391718 59809
rect 388718 59735 388720 59744
rect 388628 59706 388680 59712
rect 388772 59735 388774 59744
rect 391388 59764 391440 59770
rect 388720 59706 388772 59712
rect 394606 59800 394662 59809
rect 391662 59735 391664 59744
rect 391388 59706 391440 59712
rect 391716 59735 391718 59744
rect 394148 59764 394200 59770
rect 391664 59706 391716 59712
rect 394606 59735 394662 59744
rect 395710 59800 395766 59809
rect 398470 59800 398526 59809
rect 395710 59735 395712 59744
rect 394148 59706 394200 59712
rect 385682 59664 385738 59673
rect 385682 59599 385738 59608
rect 384854 59392 384910 59401
rect 384854 59327 384910 59336
rect 383936 50516 383988 50522
rect 383936 50458 383988 50464
rect 383016 33992 383068 33998
rect 383016 33934 383068 33940
rect 385696 20126 385724 59599
rect 388442 59528 388498 59537
rect 388442 59463 388498 59472
rect 387062 59392 387118 59401
rect 387062 59327 387118 59336
rect 387076 38146 387104 59327
rect 387064 38140 387116 38146
rect 387064 38082 387116 38088
rect 387800 36644 387852 36650
rect 387800 36586 387852 36592
rect 385776 21616 385828 21622
rect 385776 21558 385828 21564
rect 385684 20120 385736 20126
rect 385684 20062 385736 20068
rect 384764 7608 384816 7614
rect 384764 7550 384816 7556
rect 383568 3800 383620 3806
rect 383568 3742 383620 3748
rect 382924 3392 382976 3398
rect 382924 3334 382976 3340
rect 383580 480 383608 3742
rect 384776 480 384804 7550
rect 385788 3806 385816 21558
rect 386696 11892 386748 11898
rect 386696 11834 386748 11840
rect 385960 6384 386012 6390
rect 385960 6326 386012 6332
rect 385776 3800 385828 3806
rect 385776 3742 385828 3748
rect 385972 480 386000 6326
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 370566 -960 370678 326
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 386708 354 386736 11834
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 36586
rect 388456 6458 388484 59463
rect 388640 6526 388668 59706
rect 391202 59528 391258 59537
rect 391202 59463 391258 59472
rect 389822 59392 389878 59401
rect 389822 59327 389878 59336
rect 388628 6520 388680 6526
rect 388628 6462 388680 6468
rect 388444 6452 388496 6458
rect 388444 6394 388496 6400
rect 389836 6390 389864 59327
rect 391216 38078 391244 59463
rect 391400 43586 391428 59706
rect 393594 59528 393650 59537
rect 393594 59463 393650 59472
rect 392674 59392 392730 59401
rect 392674 59327 392730 59336
rect 392584 58812 392636 58818
rect 392584 58754 392636 58760
rect 391388 43580 391440 43586
rect 391388 43522 391440 43528
rect 391204 38072 391256 38078
rect 391204 38014 391256 38020
rect 390560 17332 390612 17338
rect 390560 17274 390612 17280
rect 389824 6384 389876 6390
rect 389824 6326 389876 6332
rect 389456 6316 389508 6322
rect 389456 6258 389508 6264
rect 389468 480 389496 6258
rect 390572 3194 390600 17274
rect 390560 3188 390612 3194
rect 390560 3130 390612 3136
rect 391848 3188 391900 3194
rect 391848 3130 391900 3136
rect 390652 2916 390704 2922
rect 390652 2858 390704 2864
rect 390664 480 390692 2858
rect 391860 480 391888 3130
rect 392596 2922 392624 58754
rect 392688 39574 392716 59327
rect 393608 55214 393636 59463
rect 393608 55186 394004 55214
rect 392676 39568 392728 39574
rect 392676 39510 392728 39516
rect 393976 6254 394004 55186
rect 394160 6322 394188 59706
rect 394620 59401 394648 59735
rect 395764 59735 395766 59744
rect 398104 59764 398156 59770
rect 395712 59706 395764 59712
rect 402426 59800 402482 59809
rect 398470 59735 398472 59744
rect 398104 59706 398156 59712
rect 398524 59735 398526 59744
rect 401048 59764 401100 59770
rect 398472 59706 398524 59712
rect 405278 59800 405334 59809
rect 402426 59735 402428 59744
rect 401048 59706 401100 59712
rect 402480 59735 402482 59744
rect 405188 59764 405240 59770
rect 402428 59706 402480 59712
rect 408406 59800 408462 59809
rect 405278 59735 405280 59744
rect 405188 59706 405240 59712
rect 405332 59735 405334 59744
rect 407948 59764 408000 59770
rect 405280 59706 405332 59712
rect 410154 59800 410210 59809
rect 408462 59758 408724 59786
rect 408406 59735 408462 59744
rect 407948 59706 408000 59712
rect 395342 59664 395398 59673
rect 395342 59599 395398 59608
rect 394606 59392 394662 59401
rect 394606 59327 394662 59336
rect 394700 38004 394752 38010
rect 394700 37946 394752 37952
rect 394712 16574 394740 37946
rect 395356 17338 395384 59599
rect 396722 59392 396778 59401
rect 396722 59327 396778 59336
rect 395344 17332 395396 17338
rect 395344 17274 395396 17280
rect 394712 16546 395384 16574
rect 394240 9172 394292 9178
rect 394240 9114 394292 9120
rect 394148 6316 394200 6322
rect 394148 6258 394200 6264
rect 393044 6248 393096 6254
rect 393044 6190 393096 6196
rect 393964 6248 394016 6254
rect 393964 6190 394016 6196
rect 392584 2916 392636 2922
rect 392584 2858 392636 2864
rect 393056 480 393084 6190
rect 394252 480 394280 9114
rect 395356 480 395384 16546
rect 396736 6186 396764 59327
rect 398116 40934 398144 59706
rect 398286 59528 398342 59537
rect 398286 59463 398342 59472
rect 398300 42294 398328 59463
rect 399390 59392 399446 59401
rect 400862 59392 400918 59401
rect 399446 59350 399524 59378
rect 399390 59327 399446 59336
rect 399496 45082 399524 59350
rect 400862 59327 400918 59336
rect 399484 45076 399536 45082
rect 399484 45018 399536 45024
rect 398288 42288 398340 42294
rect 398288 42230 398340 42236
rect 398104 40928 398156 40934
rect 398104 40870 398156 40876
rect 398840 39432 398892 39438
rect 398840 39374 398892 39380
rect 398852 16574 398880 39374
rect 400876 18766 400904 59327
rect 401060 46374 401088 59706
rect 402334 59664 402390 59673
rect 402334 59599 402390 59608
rect 402242 59528 402298 59537
rect 402242 59463 402298 59472
rect 402256 49162 402284 59463
rect 402348 59401 402376 59599
rect 405002 59528 405058 59537
rect 405002 59463 405058 59472
rect 402334 59392 402390 59401
rect 402334 59327 402390 59336
rect 403622 59392 403678 59401
rect 403622 59327 403678 59336
rect 402244 49156 402296 49162
rect 402244 49098 402296 49104
rect 401048 46368 401100 46374
rect 401048 46310 401100 46316
rect 401600 40792 401652 40798
rect 401600 40734 401652 40740
rect 400956 29844 401008 29850
rect 400956 29786 401008 29792
rect 400864 18760 400916 18766
rect 400864 18702 400916 18708
rect 398852 16546 398972 16574
rect 396540 6180 396592 6186
rect 396540 6122 396592 6128
rect 396724 6180 396776 6186
rect 396724 6122 396776 6128
rect 396552 480 396580 6122
rect 397736 3188 397788 3194
rect 397736 3130 397788 3136
rect 397748 480 397776 3130
rect 398944 480 398972 16546
rect 400128 7948 400180 7954
rect 400128 7890 400180 7896
rect 400140 480 400168 7890
rect 400968 3194 400996 29786
rect 401612 16574 401640 40734
rect 403636 35290 403664 59327
rect 405016 36650 405044 59463
rect 405200 47734 405228 59706
rect 407762 59528 407818 59537
rect 407762 59463 407818 59472
rect 406382 59392 406438 59401
rect 406382 59327 406438 59336
rect 405188 47728 405240 47734
rect 405188 47670 405240 47676
rect 405740 42152 405792 42158
rect 405740 42094 405792 42100
rect 405004 36644 405056 36650
rect 405004 36586 405056 36592
rect 403624 35284 403676 35290
rect 403624 35226 403676 35232
rect 403624 33924 403676 33930
rect 403624 33866 403676 33872
rect 401612 16546 402560 16574
rect 401324 3800 401376 3806
rect 401324 3742 401376 3748
rect 400956 3188 401008 3194
rect 400956 3130 401008 3136
rect 401336 480 401364 3742
rect 402532 480 402560 16546
rect 403636 3806 403664 33866
rect 404360 20188 404412 20194
rect 404360 20130 404412 20136
rect 403716 7880 403768 7886
rect 403716 7822 403768 7828
rect 403624 3800 403676 3806
rect 403624 3742 403676 3748
rect 403728 3482 403756 7822
rect 403636 3454 403756 3482
rect 403636 480 403664 3454
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 20130
rect 405752 16574 405780 42094
rect 405752 16546 406056 16574
rect 406028 480 406056 16546
rect 406396 8158 406424 59327
rect 406384 8152 406436 8158
rect 406384 8094 406436 8100
rect 407776 8022 407804 59463
rect 407960 8090 407988 59706
rect 408696 59673 408724 59758
rect 412086 59800 412142 59809
rect 410154 59735 410156 59744
rect 410208 59735 410210 59744
rect 411904 59764 411956 59770
rect 410156 59706 410208 59712
rect 412454 59800 412510 59809
rect 412142 59758 412454 59786
rect 412086 59735 412142 59744
rect 412454 59735 412510 59744
rect 413098 59800 413154 59809
rect 427450 59800 427506 59809
rect 413098 59735 413100 59744
rect 411904 59706 411956 59712
rect 413152 59735 413154 59744
rect 414664 59764 414716 59770
rect 413100 59706 413152 59712
rect 427450 59735 427506 59744
rect 427634 59800 427690 59809
rect 427634 59735 427690 59744
rect 434442 59800 434498 59809
rect 438030 59800 438086 59809
rect 434498 59758 434944 59786
rect 434442 59735 434498 59744
rect 414664 59706 414716 59712
rect 408682 59664 408738 59673
rect 408682 59599 408738 59608
rect 410154 59664 410210 59673
rect 410154 59599 410210 59608
rect 410168 59401 410196 59599
rect 410522 59528 410578 59537
rect 410522 59463 410578 59472
rect 409142 59392 409198 59401
rect 409142 59327 409198 59336
rect 410154 59392 410210 59401
rect 410154 59327 410210 59336
rect 408500 18692 408552 18698
rect 408500 18634 408552 18640
rect 407948 8084 408000 8090
rect 407948 8026 408000 8032
rect 407764 8016 407816 8022
rect 407764 7958 407816 7964
rect 407212 7812 407264 7818
rect 407212 7754 407264 7760
rect 407224 480 407252 7754
rect 408512 6914 408540 18634
rect 409156 7954 409184 59327
rect 409144 7948 409196 7954
rect 409144 7890 409196 7896
rect 410536 7818 410564 59463
rect 410706 59392 410762 59401
rect 410706 59327 410762 59336
rect 410720 7886 410748 59327
rect 410708 7880 410760 7886
rect 410708 7822 410760 7828
rect 410524 7812 410576 7818
rect 410524 7754 410576 7760
rect 411916 7750 411944 59706
rect 413926 59664 413982 59673
rect 413926 59599 413982 59608
rect 413940 59401 413968 59599
rect 414018 59528 414074 59537
rect 414018 59463 414074 59472
rect 413098 59392 413154 59401
rect 413098 59327 413154 59336
rect 413926 59392 413982 59401
rect 413926 59327 413982 59336
rect 413112 55214 413140 59327
rect 413112 55186 413324 55214
rect 412640 44940 412692 44946
rect 412640 44882 412692 44888
rect 412272 9240 412324 9246
rect 412272 9182 412324 9188
rect 410800 7744 410852 7750
rect 410800 7686 410852 7692
rect 411904 7744 411956 7750
rect 411904 7686 411956 7692
rect 408512 6886 409184 6914
rect 408408 3800 408460 3806
rect 408408 3742 408460 3748
rect 408420 480 408448 3742
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 6886
rect 410812 480 410840 7686
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 354 411986 480
rect 412284 354 412312 9182
rect 411874 326 412312 354
rect 412652 354 412680 44882
rect 413296 7682 413324 55186
rect 414032 13122 414060 59463
rect 414020 13116 414072 13122
rect 414020 13058 414072 13064
rect 414296 8288 414348 8294
rect 414296 8230 414348 8236
rect 413284 7676 413336 7682
rect 413284 7618 413336 7624
rect 414308 480 414336 8230
rect 414676 7614 414704 59706
rect 418158 59664 418214 59673
rect 418158 59599 418214 59608
rect 419814 59664 419870 59673
rect 419814 59599 419816 59608
rect 415030 59528 415086 59537
rect 417054 59528 417110 59537
rect 415086 59486 415624 59514
rect 415030 59463 415086 59472
rect 415596 59401 415624 59486
rect 417054 59463 417110 59472
rect 415398 59392 415454 59401
rect 415398 59327 415454 59336
rect 415582 59392 415638 59401
rect 415582 59327 415638 59336
rect 416870 59392 416926 59401
rect 416870 59327 416926 59336
rect 415412 33862 415440 59327
rect 416884 49026 416912 59327
rect 416872 49020 416924 49026
rect 416872 48962 416924 48968
rect 415400 33856 415452 33862
rect 415400 33798 415452 33804
rect 415400 20052 415452 20058
rect 415400 19994 415452 20000
rect 414664 7608 414716 7614
rect 414664 7550 414716 7556
rect 415412 3534 415440 19994
rect 417068 15910 417096 59463
rect 418172 53174 418200 59599
rect 419868 59599 419870 59608
rect 421104 59628 421156 59634
rect 419816 59570 419868 59576
rect 421104 59570 421156 59576
rect 419538 59528 419594 59537
rect 419538 59463 419594 59472
rect 418804 54732 418856 54738
rect 418804 54674 418856 54680
rect 418160 53168 418212 53174
rect 418160 53110 418212 53116
rect 417056 15904 417108 15910
rect 417056 15846 417108 15852
rect 417884 8220 417936 8226
rect 417884 8162 417936 8168
rect 415492 3732 415544 3738
rect 415492 3674 415544 3680
rect 415400 3528 415452 3534
rect 415400 3470 415452 3476
rect 415504 480 415532 3674
rect 416688 3528 416740 3534
rect 416688 3470 416740 3476
rect 416700 480 416728 3470
rect 417896 480 417924 8162
rect 418816 3806 418844 54674
rect 419552 29646 419580 59463
rect 419540 29640 419592 29646
rect 419540 29582 419592 29588
rect 420920 28484 420972 28490
rect 420920 28426 420972 28432
rect 419540 21480 419592 21486
rect 419540 21422 419592 21428
rect 419552 16574 419580 21422
rect 419552 16546 420224 16574
rect 418804 3800 418856 3806
rect 418804 3742 418856 3748
rect 418986 3360 419042 3369
rect 418986 3295 419042 3304
rect 419000 480 419028 3295
rect 420196 480 420224 16546
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 411874 -960 411986 326
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 420932 354 420960 28426
rect 421116 3398 421144 59570
rect 421838 59528 421894 59537
rect 421838 59463 421894 59472
rect 424782 59528 424838 59537
rect 426530 59528 426586 59537
rect 424838 59486 425284 59514
rect 424782 59463 424838 59472
rect 421852 59129 421880 59463
rect 425256 59401 425284 59486
rect 426530 59463 426586 59472
rect 425058 59392 425114 59401
rect 425058 59327 425114 59336
rect 425242 59392 425298 59401
rect 425242 59327 425298 59336
rect 422390 59256 422446 59265
rect 422390 59191 422446 59200
rect 423954 59256 424010 59265
rect 423954 59191 424010 59200
rect 421286 59120 421342 59129
rect 421286 59055 421342 59064
rect 421838 59120 421894 59129
rect 421838 59055 421894 59064
rect 421300 3466 421328 59055
rect 422404 3602 422432 59191
rect 423680 46300 423732 46306
rect 423680 46242 423732 46248
rect 422576 8220 422628 8226
rect 422576 8162 422628 8168
rect 422392 3596 422444 3602
rect 422392 3538 422444 3544
rect 421288 3460 421340 3466
rect 421288 3402 421340 3408
rect 421104 3392 421156 3398
rect 421104 3334 421156 3340
rect 422588 480 422616 8162
rect 423692 3346 423720 46242
rect 423772 32632 423824 32638
rect 423772 32574 423824 32580
rect 423784 3534 423812 32574
rect 423968 13190 423996 59191
rect 424138 59120 424194 59129
rect 424138 59055 424194 59064
rect 423956 13184 424008 13190
rect 423956 13126 424008 13132
rect 424152 3670 424180 59055
rect 425072 39370 425100 59327
rect 426544 42090 426572 59463
rect 427464 59401 427492 59735
rect 426714 59392 426770 59401
rect 426714 59327 426770 59336
rect 427450 59392 427506 59401
rect 427450 59327 427506 59336
rect 426532 42084 426584 42090
rect 426532 42026 426584 42032
rect 426728 40730 426756 59327
rect 427648 55962 427676 59735
rect 427910 59664 427966 59673
rect 427910 59599 427966 59608
rect 427820 58880 427872 58886
rect 427820 58822 427872 58828
rect 427636 55956 427688 55962
rect 427636 55898 427688 55904
rect 426716 40724 426768 40730
rect 426716 40666 426768 40672
rect 425060 39364 425112 39370
rect 425060 39306 425112 39312
rect 426440 22840 426492 22846
rect 426440 22782 426492 22788
rect 426452 16574 426480 22782
rect 427832 16574 427860 58822
rect 427924 37942 427952 59599
rect 430578 59528 430634 59537
rect 430578 59463 430634 59472
rect 433522 59528 433578 59537
rect 433522 59463 433578 59472
rect 429198 59256 429254 59265
rect 429198 59191 429254 59200
rect 429212 43450 429240 59191
rect 430592 57322 430620 59463
rect 432050 59392 432106 59401
rect 432050 59327 432106 59336
rect 430670 59256 430726 59265
rect 430670 59191 430726 59200
rect 430580 57316 430632 57322
rect 430580 57258 430632 57264
rect 430580 54664 430632 54670
rect 430580 54606 430632 54612
rect 429200 43444 429252 43450
rect 429200 43386 429252 43392
rect 427912 37936 427964 37942
rect 427912 37878 427964 37884
rect 430592 16574 430620 54606
rect 430684 51814 430712 59191
rect 430672 51808 430724 51814
rect 430672 51750 430724 51756
rect 432064 45554 432092 59327
rect 431972 45526 432092 45554
rect 431972 28354 432000 45526
rect 433536 44878 433564 59463
rect 434916 59401 434944 59758
rect 441986 59800 442042 59809
rect 438030 59735 438032 59744
rect 438084 59735 438086 59744
rect 438860 59764 438912 59770
rect 438032 59706 438084 59712
rect 441986 59735 442042 59744
rect 446402 59800 446458 59809
rect 446402 59735 446458 59744
rect 448150 59800 448206 59809
rect 448150 59735 448206 59744
rect 453946 59800 454002 59809
rect 461582 59800 461638 59809
rect 454002 59758 454264 59786
rect 453946 59735 454002 59744
rect 438860 59706 438912 59712
rect 437570 59664 437626 59673
rect 437570 59599 437626 59608
rect 436190 59528 436246 59537
rect 436190 59463 436246 59472
rect 434718 59392 434774 59401
rect 434718 59327 434774 59336
rect 434902 59392 434958 59401
rect 434902 59327 434958 59336
rect 433524 44872 433576 44878
rect 433524 44814 433576 44820
rect 434732 32502 434760 59327
rect 434720 32496 434772 32502
rect 434720 32438 434772 32444
rect 431960 28348 432012 28354
rect 431960 28290 432012 28296
rect 433340 24200 433392 24206
rect 433340 24142 433392 24148
rect 433352 16574 433380 24142
rect 426452 16546 426848 16574
rect 427832 16546 428504 16574
rect 430592 16546 430896 16574
rect 433352 16546 434024 16574
rect 424140 3664 424192 3670
rect 424140 3606 424192 3612
rect 423772 3528 423824 3534
rect 423772 3470 423824 3476
rect 424968 3528 425020 3534
rect 424968 3470 425020 3476
rect 423692 3318 423812 3346
rect 423784 480 423812 3318
rect 424980 480 425008 3470
rect 426164 3460 426216 3466
rect 426164 3402 426216 3408
rect 426176 480 426204 3402
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 426820 354 426848 16546
rect 428476 480 428504 16546
rect 429660 9308 429712 9314
rect 429660 9250 429712 9256
rect 429672 480 429700 9250
rect 430868 480 430896 16546
rect 432052 10804 432104 10810
rect 432052 10746 432104 10752
rect 432064 480 432092 10746
rect 433248 3528 433300 3534
rect 433248 3470 433300 3476
rect 433260 480 433288 3470
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 436204 14550 436232 59463
rect 436374 59392 436430 59401
rect 436374 59327 436430 59336
rect 436192 14544 436244 14550
rect 436192 14486 436244 14492
rect 436388 14482 436416 59327
rect 437480 25696 437532 25702
rect 437480 25638 437532 25644
rect 436376 14476 436428 14482
rect 436376 14418 436428 14424
rect 435088 10736 435140 10742
rect 435088 10678 435140 10684
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 10678
rect 436744 3596 436796 3602
rect 436744 3538 436796 3544
rect 436756 480 436784 3538
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 25638
rect 437584 14618 437612 59599
rect 438872 14686 438900 59706
rect 441066 59664 441122 59673
rect 441066 59599 441122 59608
rect 441080 59401 441108 59599
rect 440514 59392 440570 59401
rect 440514 59327 440570 59336
rect 441066 59392 441122 59401
rect 441066 59327 441122 59336
rect 441618 59392 441674 59401
rect 441618 59327 441674 59336
rect 440330 59120 440386 59129
rect 440330 59055 440386 59064
rect 440344 14754 440372 59055
rect 440528 14822 440556 59327
rect 441632 14890 441660 59327
rect 442000 58750 442028 59735
rect 443090 59664 443146 59673
rect 443090 59599 443146 59608
rect 441988 58744 442040 58750
rect 441988 58686 442040 58692
rect 443104 15026 443132 59599
rect 445758 59528 445814 59537
rect 445758 59463 445814 59472
rect 443274 59392 443330 59401
rect 443274 59327 443330 59336
rect 443092 15020 443144 15026
rect 443092 14962 443144 14968
rect 443288 14958 443316 59327
rect 445772 46238 445800 59463
rect 446416 58138 446444 59735
rect 446954 59664 447010 59673
rect 446954 59599 447010 59608
rect 447138 59664 447194 59673
rect 447138 59599 447194 59608
rect 446404 58132 446456 58138
rect 446404 58074 446456 58080
rect 446968 57974 446996 59599
rect 447152 58954 447180 59599
rect 447140 58948 447192 58954
rect 447140 58890 447192 58896
rect 448164 58410 448192 59735
rect 449990 59528 450046 59537
rect 449990 59463 450046 59472
rect 453026 59528 453082 59537
rect 453026 59463 453082 59472
rect 448520 58948 448572 58954
rect 448520 58890 448572 58896
rect 448152 58404 448204 58410
rect 448152 58346 448204 58352
rect 447416 58132 447468 58138
rect 447416 58074 447468 58080
rect 446968 57946 447180 57974
rect 447152 47666 447180 57946
rect 447140 47660 447192 47666
rect 447140 47602 447192 47608
rect 445760 46232 445812 46238
rect 445760 46174 445812 46180
rect 444380 26988 444432 26994
rect 444380 26930 444432 26936
rect 444392 16574 444420 26930
rect 447428 25634 447456 58074
rect 448532 54602 448560 58890
rect 448520 54596 448572 54602
rect 448520 54538 448572 54544
rect 447416 25628 447468 25634
rect 447416 25570 447468 25576
rect 444392 16546 445064 16574
rect 443276 14952 443328 14958
rect 443276 14894 443328 14900
rect 441620 14884 441672 14890
rect 441620 14826 441672 14832
rect 440516 14816 440568 14822
rect 440516 14758 440568 14764
rect 440332 14748 440384 14754
rect 440332 14690 440384 14696
rect 438860 14680 438912 14686
rect 438860 14622 438912 14628
rect 437572 14612 437624 14618
rect 437572 14554 437624 14560
rect 440884 14476 440936 14482
rect 440884 14418 440936 14424
rect 439136 10668 439188 10674
rect 439136 10610 439188 10616
rect 439148 480 439176 10610
rect 440896 3738 440924 14418
rect 442632 10600 442684 10606
rect 442632 10542 442684 10548
rect 441528 9104 441580 9110
rect 441528 9046 441580 9052
rect 440884 3732 440936 3738
rect 440884 3674 440936 3680
rect 440332 3664 440384 3670
rect 440332 3606 440384 3612
rect 440344 480 440372 3606
rect 441540 480 441568 9046
rect 442644 480 442672 10542
rect 443828 3732 443880 3738
rect 443828 3674 443880 3680
rect 443840 480 443868 3674
rect 445036 480 445064 16546
rect 450004 16046 450032 59463
rect 452842 59392 452898 59401
rect 452842 59327 452898 59336
rect 451278 59256 451334 59265
rect 451278 59191 451334 59200
rect 450176 58404 450228 58410
rect 450176 58346 450228 58352
rect 449992 16040 450044 16046
rect 449992 15982 450044 15988
rect 450188 15978 450216 58346
rect 451292 16114 451320 59191
rect 452660 43648 452712 43654
rect 452660 43590 452712 43596
rect 451280 16108 451332 16114
rect 451280 16050 451332 16056
rect 450176 15972 450228 15978
rect 450176 15914 450228 15920
rect 445760 10532 445812 10538
rect 445760 10474 445812 10480
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 354 445800 10474
rect 448520 10464 448572 10470
rect 448520 10406 448572 10412
rect 447416 3800 447468 3806
rect 447416 3742 447468 3748
rect 447428 480 447456 3742
rect 448532 3398 448560 10406
rect 448612 9036 448664 9042
rect 448612 8978 448664 8984
rect 448520 3392 448572 3398
rect 448520 3334 448572 3340
rect 448624 480 448652 8978
rect 452108 8968 452160 8974
rect 452108 8910 452160 8916
rect 450912 3868 450964 3874
rect 450912 3810 450964 3816
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 449820 480 449848 3334
rect 450924 480 450952 3810
rect 452120 480 452148 8910
rect 452672 6914 452700 43590
rect 452856 16182 452884 59327
rect 453040 16250 453068 59463
rect 454236 59401 454264 59758
rect 456616 59764 456668 59770
rect 456616 59706 456668 59712
rect 457076 59764 457128 59770
rect 463606 59800 463662 59809
rect 461582 59735 461584 59744
rect 457076 59706 457128 59712
rect 461636 59735 461638 59744
rect 462412 59764 462464 59770
rect 461584 59706 461636 59712
rect 463606 59735 463662 59744
rect 467562 59800 467618 59809
rect 470598 59800 470654 59809
rect 467618 59758 468064 59786
rect 467562 59735 467618 59744
rect 462412 59706 462464 59712
rect 455878 59664 455934 59673
rect 455878 59599 455934 59608
rect 455892 59401 455920 59599
rect 456628 59537 456656 59706
rect 456890 59664 456946 59673
rect 456890 59599 456892 59608
rect 456944 59599 456946 59608
rect 456892 59570 456944 59576
rect 456614 59528 456670 59537
rect 456614 59463 456670 59472
rect 456890 59528 456946 59537
rect 456890 59463 456946 59472
rect 454038 59392 454094 59401
rect 454038 59327 454094 59336
rect 454222 59392 454278 59401
rect 454222 59327 454278 59336
rect 455510 59392 455566 59401
rect 455510 59327 455566 59336
rect 455878 59392 455934 59401
rect 455878 59327 455934 59336
rect 454052 16318 454080 59327
rect 455420 29776 455472 29782
rect 455420 29718 455472 29724
rect 454040 16312 454092 16318
rect 454040 16254 454092 16260
rect 453028 16244 453080 16250
rect 453028 16186 453080 16192
rect 452844 16176 452896 16182
rect 452844 16118 452896 16124
rect 455432 6914 455460 29718
rect 455524 16386 455552 59327
rect 456904 16522 456932 59463
rect 456892 16516 456944 16522
rect 456892 16458 456944 16464
rect 457088 16454 457116 59706
rect 460938 59664 460994 59673
rect 458272 59628 458324 59634
rect 460938 59599 460994 59608
rect 458272 59570 458324 59576
rect 458180 49088 458232 49094
rect 458180 49030 458232 49036
rect 458192 16574 458220 49030
rect 458284 21554 458312 59570
rect 459834 59528 459890 59537
rect 459834 59463 459890 59472
rect 459650 59392 459706 59401
rect 459650 59327 459706 59336
rect 458272 21548 458324 21554
rect 458272 21490 458324 21496
rect 458192 16546 459232 16574
rect 457076 16448 457128 16454
rect 457076 16390 457128 16396
rect 455512 16380 455564 16386
rect 455512 16322 455564 16328
rect 456892 10396 456944 10402
rect 456892 10338 456944 10344
rect 452672 6886 453344 6914
rect 455432 6886 455736 6914
rect 453316 480 453344 6886
rect 454500 3936 454552 3942
rect 454500 3878 454552 3884
rect 454512 480 454540 3878
rect 455708 480 455736 6886
rect 456904 480 456932 10338
rect 458088 4004 458140 4010
rect 458088 3946 458140 3952
rect 458100 480 458128 3946
rect 459204 480 459232 16546
rect 459664 13258 459692 59327
rect 459848 13326 459876 59463
rect 460952 13394 460980 59599
rect 462320 31136 462372 31142
rect 462320 31078 462372 31084
rect 460940 13388 460992 13394
rect 460940 13330 460992 13336
rect 459836 13320 459888 13326
rect 459836 13262 459888 13268
rect 459652 13252 459704 13258
rect 459652 13194 459704 13200
rect 459928 10328 459980 10334
rect 459928 10270 459980 10276
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 10270
rect 461584 8968 461636 8974
rect 461584 8910 461636 8916
rect 461596 480 461624 8910
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 31078
rect 462424 13462 462452 59706
rect 463620 56030 463648 59735
rect 463698 59528 463754 59537
rect 463698 59463 463754 59472
rect 466642 59528 466698 59537
rect 466642 59463 466698 59472
rect 463608 56024 463660 56030
rect 463608 55966 463660 55972
rect 463712 51882 463740 59463
rect 463882 59392 463938 59401
rect 463882 59327 463938 59336
rect 465078 59392 465134 59401
rect 465078 59327 465134 59336
rect 463700 51876 463752 51882
rect 463700 51818 463752 51824
rect 463700 33992 463752 33998
rect 463700 33934 463752 33940
rect 463712 16574 463740 33934
rect 463896 22914 463924 59327
rect 465092 50454 465120 59327
rect 466460 50516 466512 50522
rect 466460 50458 466512 50464
rect 465080 50448 465132 50454
rect 465080 50390 465132 50396
rect 465080 47592 465132 47598
rect 465080 47534 465132 47540
rect 463884 22908 463936 22914
rect 463884 22850 463936 22856
rect 465092 16574 465120 47534
rect 466472 16574 466500 50458
rect 466656 24274 466684 59463
rect 468036 59401 468064 59758
rect 474370 59800 474426 59809
rect 470598 59735 470600 59744
rect 470652 59735 470654 59744
rect 471980 59764 472032 59770
rect 470600 59706 470652 59712
rect 480258 59800 480314 59809
rect 474370 59735 474372 59744
rect 471980 59706 472032 59712
rect 474424 59735 474426 59744
rect 476396 59764 476448 59770
rect 474372 59706 474424 59712
rect 483294 59800 483350 59809
rect 480258 59735 480260 59744
rect 476396 59706 476448 59712
rect 480312 59735 480314 59744
rect 481640 59764 481692 59770
rect 480260 59706 480312 59712
rect 483294 59735 483350 59744
rect 483478 59800 483534 59809
rect 483478 59735 483534 59744
rect 488446 59800 488502 59809
rect 488446 59735 488502 59744
rect 488630 59800 488686 59809
rect 488630 59735 488686 59744
rect 495898 59800 495954 59809
rect 500682 59800 500738 59809
rect 495898 59735 495900 59744
rect 481640 59706 481692 59712
rect 470552 59664 470608 59673
rect 470608 59622 470732 59650
rect 470552 59599 470608 59608
rect 469310 59528 469366 59537
rect 469310 59463 469366 59472
rect 467838 59392 467894 59401
rect 467838 59327 467894 59336
rect 468022 59392 468078 59401
rect 468022 59327 468078 59336
rect 466644 24268 466696 24274
rect 466644 24210 466696 24216
rect 463712 16546 464016 16574
rect 465092 16546 465856 16574
rect 466472 16546 467512 16574
rect 462412 13456 462464 13462
rect 462412 13398 462464 13404
rect 463988 480 464016 16546
rect 465172 4072 465224 4078
rect 465172 4014 465224 4020
rect 465184 480 465212 4014
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 354 465856 16546
rect 467484 480 467512 16546
rect 467852 11762 467880 59327
rect 469324 40866 469352 59463
rect 469494 59392 469550 59401
rect 469494 59327 469550 59336
rect 469312 40860 469364 40866
rect 469312 40802 469364 40808
rect 469508 39506 469536 59327
rect 470600 57384 470652 57390
rect 470600 57326 470652 57332
rect 469496 39500 469548 39506
rect 469496 39442 469548 39448
rect 469220 35216 469272 35222
rect 469220 35158 469272 35164
rect 469232 16574 469260 35158
rect 469232 16546 469904 16574
rect 467840 11756 467892 11762
rect 467840 11698 467892 11704
rect 468668 4140 468720 4146
rect 468668 4082 468720 4088
rect 468680 480 468708 4082
rect 469876 480 469904 16546
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 354 470640 57326
rect 470704 27062 470732 59622
rect 471992 42226 472020 59706
rect 476302 59664 476358 59673
rect 476302 59599 476358 59608
rect 473634 59528 473690 59537
rect 473634 59463 473690 59472
rect 476210 59528 476266 59537
rect 476210 59463 476266 59472
rect 473450 59392 473506 59401
rect 473450 59327 473506 59336
rect 473464 45014 473492 59327
rect 473452 45008 473504 45014
rect 473452 44950 473504 44956
rect 471980 42220 472032 42226
rect 471980 42162 472032 42168
rect 473360 36576 473412 36582
rect 473360 36518 473412 36524
rect 470692 27056 470744 27062
rect 470692 26998 470744 27004
rect 473372 6914 473400 36518
rect 473648 35358 473676 59463
rect 474738 59392 474794 59401
rect 474738 59327 474794 59336
rect 473636 35352 473688 35358
rect 473636 35294 473688 35300
rect 473452 20120 473504 20126
rect 473452 20062 473504 20068
rect 473464 16574 473492 20062
rect 474752 17406 474780 59327
rect 476120 53236 476172 53242
rect 476120 53178 476172 53184
rect 474740 17400 474792 17406
rect 474740 17342 474792 17348
rect 476132 16574 476160 53178
rect 476224 31210 476252 59463
rect 476316 59401 476344 59599
rect 476302 59392 476358 59401
rect 476302 59327 476358 59336
rect 476408 36718 476436 59706
rect 478326 59664 478382 59673
rect 478326 59599 478382 59608
rect 480258 59664 480314 59673
rect 480314 59622 480484 59650
rect 480258 59599 480314 59608
rect 478340 59401 478368 59599
rect 478878 59528 478934 59537
rect 478878 59463 478934 59472
rect 477590 59392 477646 59401
rect 477590 59327 477646 59336
rect 478326 59392 478382 59401
rect 478326 59327 478382 59336
rect 477500 38140 477552 38146
rect 477500 38082 477552 38088
rect 476396 36712 476448 36718
rect 476396 36654 476448 36660
rect 476212 31204 476264 31210
rect 476212 31146 476264 31152
rect 473464 16546 474136 16574
rect 476132 16546 476528 16574
rect 473372 6886 473492 6914
rect 472256 3392 472308 3398
rect 472256 3334 472308 3340
rect 472268 480 472296 3334
rect 473464 480 473492 6886
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 16546
rect 475752 3324 475804 3330
rect 475752 3266 475804 3272
rect 475764 480 475792 3266
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 477512 6914 477540 38082
rect 477604 11830 477632 59327
rect 478892 18834 478920 59463
rect 480350 59256 480406 59265
rect 480350 59191 480406 59200
rect 480364 49230 480392 59191
rect 480352 49224 480404 49230
rect 480352 49166 480404 49172
rect 480456 46442 480484 59622
rect 480444 46436 480496 46442
rect 480444 46378 480496 46384
rect 481652 28422 481680 59706
rect 483110 59528 483166 59537
rect 483110 59463 483166 59472
rect 483124 43518 483152 59463
rect 483308 59401 483336 59735
rect 483294 59392 483350 59401
rect 483294 59327 483350 59336
rect 483294 59256 483350 59265
rect 483294 59191 483350 59200
rect 483112 43512 483164 43518
rect 483112 43454 483164 43460
rect 483308 32570 483336 59191
rect 483492 58818 483520 59735
rect 484398 59664 484454 59673
rect 484398 59599 484454 59608
rect 487066 59664 487122 59673
rect 487066 59599 487122 59608
rect 483480 58812 483532 58818
rect 483480 58754 483532 58760
rect 483296 32564 483348 32570
rect 483296 32506 483348 32512
rect 481640 28416 481692 28422
rect 481640 28358 481692 28364
rect 484412 21622 484440 59599
rect 487080 59401 487108 59599
rect 488460 59537 488488 59735
rect 487250 59528 487306 59537
rect 487250 59463 487306 59472
rect 488446 59528 488502 59537
rect 488446 59463 488502 59472
rect 485962 59392 486018 59401
rect 485962 59327 486018 59336
rect 487066 59392 487122 59401
rect 487066 59327 487122 59336
rect 484400 21616 484452 21622
rect 484400 21558 484452 21564
rect 478880 18828 478932 18834
rect 478880 18770 478932 18776
rect 483020 18624 483072 18630
rect 483020 18566 483072 18572
rect 480260 17264 480312 17270
rect 480260 17206 480312 17212
rect 480272 16574 480300 17206
rect 483032 16574 483060 18566
rect 480272 16546 480576 16574
rect 483032 16546 484072 16574
rect 477592 11824 477644 11830
rect 477592 11766 477644 11772
rect 477512 6886 478184 6914
rect 478156 480 478184 6886
rect 479340 3256 479392 3262
rect 479340 3198 479392 3204
rect 479352 480 479380 3198
rect 480548 480 480576 16546
rect 482376 10328 482428 10334
rect 482376 10270 482428 10276
rect 481732 6520 481784 6526
rect 481732 6462 481784 6468
rect 481744 480 481772 6462
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 354 482416 10270
rect 484044 480 484072 16546
rect 485976 11898 486004 59327
rect 487160 19984 487212 19990
rect 487160 19926 487212 19932
rect 486424 13116 486476 13122
rect 486424 13058 486476 13064
rect 485964 11892 486016 11898
rect 485964 11834 486016 11840
rect 485228 6452 485280 6458
rect 485228 6394 485280 6400
rect 485240 480 485268 6394
rect 486436 480 486464 13058
rect 482806 354 482918 480
rect 482388 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487172 354 487200 19926
rect 487264 9178 487292 59463
rect 488538 59392 488594 59401
rect 488538 59327 488594 59336
rect 488552 29850 488580 59327
rect 488644 54738 488672 59735
rect 495952 59735 495954 59744
rect 496912 59764 496964 59770
rect 495900 59706 495952 59712
rect 503626 59800 503682 59809
rect 500682 59735 500684 59744
rect 496912 59706 496964 59712
rect 500736 59735 500738 59744
rect 502616 59764 502668 59770
rect 500684 59706 500736 59712
rect 514298 59800 514354 59809
rect 503626 59735 503628 59744
rect 502616 59706 502668 59712
rect 503680 59735 503682 59744
rect 505192 59764 505244 59770
rect 503628 59706 503680 59712
rect 517242 59800 517298 59809
rect 514354 59758 514984 59786
rect 514298 59735 514354 59744
rect 505192 59706 505244 59712
rect 489918 59664 489974 59673
rect 489918 59599 489974 59608
rect 492862 59664 492918 59673
rect 492862 59599 492864 59608
rect 488632 54732 488684 54738
rect 488632 54674 488684 54680
rect 489932 51074 489960 59599
rect 492916 59599 492918 59608
rect 494152 59628 494204 59634
rect 492864 59570 492916 59576
rect 494152 59570 494204 59576
rect 490010 59528 490066 59537
rect 492954 59528 493010 59537
rect 490066 59486 490236 59514
rect 490010 59463 490066 59472
rect 489932 51046 490052 51074
rect 490024 33930 490052 51046
rect 490012 33924 490064 33930
rect 490012 33866 490064 33872
rect 488540 29844 488592 29850
rect 488540 29786 488592 29792
rect 489920 21412 489972 21418
rect 489920 21354 489972 21360
rect 487252 9172 487304 9178
rect 487252 9114 487304 9120
rect 488816 6384 488868 6390
rect 488816 6326 488868 6332
rect 488828 480 488856 6326
rect 489932 3194 489960 21354
rect 490208 20194 490236 59486
rect 492954 59463 493010 59472
rect 492770 59392 492826 59401
rect 492770 59327 492826 59336
rect 491300 43580 491352 43586
rect 491300 43522 491352 43528
rect 490196 20188 490248 20194
rect 490196 20130 490248 20136
rect 491312 16574 491340 43522
rect 491312 16546 492352 16574
rect 490012 11756 490064 11762
rect 490012 11698 490064 11704
rect 489920 3188 489972 3194
rect 489920 3130 489972 3136
rect 490024 3074 490052 11698
rect 490748 3188 490800 3194
rect 490748 3130 490800 3136
rect 489932 3046 490052 3074
rect 489932 480 489960 3046
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490760 354 490788 3130
rect 492324 480 492352 16546
rect 492784 9246 492812 59327
rect 492968 14482 492996 59463
rect 494060 58676 494112 58682
rect 494060 58618 494112 58624
rect 493048 14612 493100 14618
rect 493048 14554 493100 14560
rect 492956 14476 493008 14482
rect 492956 14418 493008 14424
rect 492772 9240 492824 9246
rect 492772 9182 492824 9188
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 14554
rect 494072 3482 494100 58618
rect 494164 3641 494192 59570
rect 495530 59392 495586 59401
rect 495530 59327 495586 59336
rect 495440 38072 495492 38078
rect 495440 38014 495492 38020
rect 494150 3632 494206 3641
rect 494150 3567 494206 3576
rect 494072 3454 494744 3482
rect 494716 480 494744 3454
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 38014
rect 495544 8226 495572 59327
rect 496924 9314 496952 59706
rect 497738 59528 497794 59537
rect 499854 59528 499910 59537
rect 497738 59463 497740 59472
rect 497792 59463 497794 59472
rect 499672 59492 499724 59498
rect 497740 59434 497792 59440
rect 499854 59463 499910 59472
rect 502430 59528 502486 59537
rect 502430 59463 502486 59472
rect 499672 59434 499724 59440
rect 498382 59392 498438 59401
rect 498382 59327 498438 59336
rect 497094 59256 497150 59265
rect 497094 59191 497150 59200
rect 496912 9308 496964 9314
rect 496912 9250 496964 9256
rect 495532 8220 495584 8226
rect 495532 8162 495584 8168
rect 497108 3466 497136 59191
rect 498200 39568 498252 39574
rect 498200 39510 498252 39516
rect 498212 3534 498240 39510
rect 498292 22772 498344 22778
rect 498292 22714 498344 22720
rect 498200 3528 498252 3534
rect 498200 3470 498252 3476
rect 497096 3460 497148 3466
rect 497096 3402 497148 3408
rect 498304 3346 498332 22714
rect 498396 3466 498424 59327
rect 499684 3602 499712 59434
rect 499868 3670 499896 59463
rect 501050 59392 501106 59401
rect 501050 59327 501106 59336
rect 500960 24132 501012 24138
rect 500960 24074 501012 24080
rect 499856 3664 499908 3670
rect 499856 3606 499908 3612
rect 499672 3596 499724 3602
rect 499672 3538 499724 3544
rect 499028 3528 499080 3534
rect 499028 3470 499080 3476
rect 498384 3460 498436 3466
rect 498384 3402 498436 3408
rect 498212 3318 498332 3346
rect 497096 3188 497148 3194
rect 497096 3130 497148 3136
rect 497108 480 497136 3130
rect 498212 480 498240 3318
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499040 354 499068 3470
rect 500592 3460 500644 3466
rect 500592 3402 500644 3408
rect 500604 480 500632 3402
rect 500972 490 501000 24074
rect 501064 3738 501092 59327
rect 502444 3874 502472 59463
rect 502432 3868 502484 3874
rect 502432 3810 502484 3816
rect 502628 3806 502656 59706
rect 503626 59664 503682 59673
rect 503682 59622 503760 59650
rect 503626 59599 503682 59608
rect 502984 6316 503036 6322
rect 502984 6258 503036 6264
rect 502616 3800 502668 3806
rect 502616 3742 502668 3748
rect 501052 3732 501104 3738
rect 501052 3674 501104 3680
rect 499366 354 499478 480
rect 499040 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 500972 462 501368 490
rect 502996 480 503024 6258
rect 503732 3942 503760 59622
rect 505100 25560 505152 25566
rect 505100 25502 505152 25508
rect 503720 3936 503772 3942
rect 503720 3878 503772 3884
rect 504180 3528 504232 3534
rect 504180 3470 504232 3476
rect 505112 3482 505140 25502
rect 505204 4010 505232 59706
rect 511998 59664 512054 59673
rect 511998 59599 512054 59608
rect 507490 59528 507546 59537
rect 510618 59528 510674 59537
rect 507490 59463 507492 59472
rect 507544 59463 507546 59472
rect 509424 59492 509476 59498
rect 507492 59434 507544 59440
rect 510618 59463 510674 59472
rect 509424 59434 509476 59440
rect 506754 59256 506810 59265
rect 506754 59191 506810 59200
rect 507950 59256 508006 59265
rect 507950 59191 508006 59200
rect 506570 59120 506626 59129
rect 506570 59055 506626 59064
rect 506584 8974 506612 59055
rect 506572 8968 506624 8974
rect 506572 8910 506624 8916
rect 506480 6248 506532 6254
rect 506480 6190 506532 6196
rect 505192 4004 505244 4010
rect 505192 3946 505244 3952
rect 504192 480 504220 3470
rect 505112 3454 505416 3482
rect 505388 480 505416 3454
rect 506492 480 506520 6190
rect 506768 4078 506796 59191
rect 507860 57248 507912 57254
rect 507860 57190 507912 57196
rect 506756 4072 506808 4078
rect 506756 4014 506808 4020
rect 507676 3596 507728 3602
rect 507676 3538 507728 3544
rect 507688 480 507716 3538
rect 507872 3482 507900 57190
rect 507964 4146 507992 59191
rect 509240 17332 509292 17338
rect 509240 17274 509292 17280
rect 509252 16574 509280 17274
rect 509252 16546 509372 16574
rect 507952 4140 508004 4146
rect 507952 4082 508004 4088
rect 507872 3454 508912 3482
rect 508884 480 508912 3454
rect 509344 490 509372 16546
rect 509436 3398 509464 59434
rect 509606 59392 509662 59401
rect 509606 59327 509662 59336
rect 509620 16574 509648 59327
rect 509620 16546 509740 16574
rect 509424 3392 509476 3398
rect 509424 3334 509476 3340
rect 509712 3330 509740 16546
rect 509700 3324 509752 3330
rect 509700 3266 509752 3272
rect 510632 3262 510660 59463
rect 512012 10334 512040 59599
rect 514956 59401 514984 59758
rect 522118 59800 522174 59809
rect 517242 59735 517244 59744
rect 517296 59735 517298 59744
rect 519176 59764 519228 59770
rect 517244 59706 517296 59712
rect 524050 59800 524106 59809
rect 522118 59735 522120 59744
rect 519176 59706 519228 59712
rect 522172 59735 522174 59744
rect 523684 59764 523736 59770
rect 522120 59706 522172 59712
rect 526994 59800 527050 59809
rect 524050 59735 524052 59744
rect 523684 59706 523736 59712
rect 524104 59735 524106 59744
rect 526444 59764 526496 59770
rect 524052 59706 524104 59712
rect 530858 59800 530914 59809
rect 526994 59735 526996 59744
rect 526444 59706 526496 59712
rect 527048 59735 527050 59744
rect 529204 59764 529256 59770
rect 526996 59706 527048 59712
rect 533802 59800 533858 59809
rect 530858 59735 530860 59744
rect 529204 59706 529256 59712
rect 530912 59735 530914 59744
rect 533528 59764 533580 59770
rect 530860 59706 530912 59712
rect 533802 59735 533804 59744
rect 533528 59706 533580 59712
rect 533856 59735 533858 59744
rect 536288 59764 536340 59770
rect 533804 59706 533856 59712
rect 536288 59706 536340 59712
rect 516322 59528 516378 59537
rect 516322 59463 516378 59472
rect 518990 59528 519046 59537
rect 518990 59463 519046 59472
rect 514758 59392 514814 59401
rect 514758 59327 514814 59336
rect 514942 59392 514998 59401
rect 514942 59327 514998 59336
rect 513654 59256 513710 59265
rect 513654 59191 513710 59200
rect 513470 59120 513526 59129
rect 513470 59055 513526 59064
rect 513484 13122 513512 59055
rect 513472 13116 513524 13122
rect 513472 13058 513524 13064
rect 513668 11762 513696 59191
rect 514772 14618 514800 59327
rect 516140 40928 516192 40934
rect 516140 40870 516192 40876
rect 516152 16574 516180 40870
rect 516152 16546 516272 16574
rect 514760 14612 514812 14618
rect 514760 14554 514812 14560
rect 513656 11756 513708 11762
rect 513656 11698 513708 11704
rect 512000 10328 512052 10334
rect 512000 10270 512052 10276
rect 513564 6180 513616 6186
rect 513564 6122 513616 6128
rect 512460 5296 512512 5302
rect 512460 5238 512512 5244
rect 511264 3664 511316 3670
rect 511264 3606 511316 3612
rect 510620 3256 510672 3262
rect 510620 3198 510672 3204
rect 501340 354 501368 462
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 509344 462 509648 490
rect 511276 480 511304 3606
rect 512472 480 512500 5238
rect 513576 480 513604 6122
rect 515956 5228 516008 5234
rect 515956 5170 516008 5176
rect 514760 3188 514812 3194
rect 514760 3130 514812 3136
rect 514772 480 514800 3130
rect 515968 480 515996 5170
rect 516140 3732 516192 3738
rect 516140 3674 516192 3680
rect 516152 3466 516180 3674
rect 516140 3460 516192 3466
rect 516140 3402 516192 3408
rect 516244 3074 516272 16546
rect 516336 3738 516364 59463
rect 516506 59392 516562 59401
rect 516506 59327 516562 59336
rect 517518 59392 517574 59401
rect 517518 59327 517574 59336
rect 516324 3732 516376 3738
rect 516324 3674 516376 3680
rect 516520 3262 516548 59327
rect 517532 3534 517560 59327
rect 518348 3800 518400 3806
rect 518348 3742 518400 3748
rect 517520 3528 517572 3534
rect 517520 3470 517572 3476
rect 516508 3256 516560 3262
rect 516508 3198 516560 3204
rect 516244 3046 517192 3074
rect 517164 480 517192 3046
rect 518360 480 518388 3742
rect 519004 3670 519032 59463
rect 518992 3664 519044 3670
rect 518992 3606 519044 3612
rect 519188 3602 519216 59706
rect 521658 59528 521714 59537
rect 521658 59463 521714 59472
rect 520370 59392 520426 59401
rect 520370 59327 520426 59336
rect 520280 42288 520332 42294
rect 520280 42230 520332 42236
rect 519544 5160 519596 5166
rect 519544 5102 519596 5108
rect 519176 3596 519228 3602
rect 519176 3538 519228 3544
rect 519556 480 519584 5102
rect 509620 354 509648 462
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520292 354 520320 42230
rect 520384 3194 520412 59327
rect 521672 3806 521700 59463
rect 523130 59256 523186 59265
rect 523130 59191 523186 59200
rect 522304 45076 522356 45082
rect 522304 45018 522356 45024
rect 521660 3800 521712 3806
rect 521660 3742 521712 3748
rect 521844 3528 521896 3534
rect 521844 3470 521896 3476
rect 520372 3188 520424 3194
rect 520372 3130 520424 3136
rect 521856 480 521884 3470
rect 522316 3058 522344 45018
rect 523144 3534 523172 59191
rect 523224 26920 523276 26926
rect 523224 26862 523276 26868
rect 523132 3528 523184 3534
rect 523132 3470 523184 3476
rect 522304 3052 522356 3058
rect 522304 2994 522356 3000
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 520710 -960 520822 326
rect 521814 -960 521926 480
rect 523010 354 523122 480
rect 523236 354 523264 26862
rect 523696 2990 523724 59706
rect 525062 59392 525118 59401
rect 525062 59327 525118 59336
rect 525076 4146 525104 59327
rect 525156 46368 525208 46374
rect 525156 46310 525208 46316
rect 525064 4140 525116 4146
rect 525064 4082 525116 4088
rect 525168 3194 525196 46310
rect 526456 3602 526484 59706
rect 526626 59528 526682 59537
rect 526626 59463 526682 59472
rect 526640 16574 526668 59463
rect 527822 59256 527878 59265
rect 527822 59191 527878 59200
rect 527836 16574 527864 59191
rect 526640 16546 526760 16574
rect 527836 16546 527956 16574
rect 526628 5092 526680 5098
rect 526628 5034 526680 5040
rect 526444 3596 526496 3602
rect 526444 3538 526496 3544
rect 525156 3188 525208 3194
rect 525156 3130 525208 3136
rect 524236 3052 524288 3058
rect 524236 2994 524288 3000
rect 523684 2984 523736 2990
rect 523684 2926 523736 2932
rect 524248 480 524276 2994
rect 525432 2984 525484 2990
rect 525432 2926 525484 2932
rect 525444 480 525472 2926
rect 526640 480 526668 5034
rect 526732 3534 526760 16546
rect 526720 3528 526772 3534
rect 526720 3470 526772 3476
rect 527928 3466 527956 16546
rect 529020 4140 529072 4146
rect 529020 4082 529072 4088
rect 527916 3460 527968 3466
rect 527916 3402 527968 3408
rect 527824 3188 527876 3194
rect 527824 3130 527876 3136
rect 527836 480 527864 3130
rect 529032 480 529060 4082
rect 529216 3330 529244 59706
rect 530766 59528 530822 59537
rect 530766 59463 530822 59472
rect 533342 59528 533398 59537
rect 533342 59463 533398 59472
rect 530582 59392 530638 59401
rect 530582 59327 530638 59336
rect 530124 5024 530176 5030
rect 530124 4966 530176 4972
rect 529204 3324 529256 3330
rect 529204 3266 529256 3272
rect 530136 480 530164 4966
rect 530596 3398 530624 59327
rect 530780 4146 530808 59463
rect 531962 59392 532018 59401
rect 531962 59327 532018 59336
rect 531412 18760 531464 18766
rect 531412 18702 531464 18708
rect 531424 6914 531452 18702
rect 531332 6886 531452 6914
rect 530768 4140 530820 4146
rect 530768 4082 530820 4088
rect 530584 3392 530636 3398
rect 530584 3334 530636 3340
rect 531332 480 531360 6886
rect 531976 4078 532004 59327
rect 532700 28280 532752 28286
rect 532700 28222 532752 28228
rect 532712 16574 532740 28222
rect 532712 16546 533292 16574
rect 531964 4072 532016 4078
rect 531964 4014 532016 4020
rect 532516 3596 532568 3602
rect 532516 3538 532568 3544
rect 532528 480 532556 3538
rect 533264 3482 533292 16546
rect 533356 3942 533384 59463
rect 533540 4010 533568 59706
rect 535734 59528 535790 59537
rect 535734 59463 535790 59472
rect 534722 59392 534778 59401
rect 534722 59327 534778 59336
rect 534080 49156 534132 49162
rect 534080 49098 534132 49104
rect 534092 16574 534120 49098
rect 534092 16546 534488 16574
rect 533528 4004 533580 4010
rect 533528 3946 533580 3952
rect 533344 3936 533396 3942
rect 533344 3878 533396 3884
rect 533264 3454 533752 3482
rect 533724 480 533752 3454
rect 523010 326 523264 354
rect 523010 -960 523122 326
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 534736 3874 534764 59327
rect 535748 55214 535776 59463
rect 535748 55186 536144 55214
rect 534724 3868 534776 3874
rect 534724 3810 534776 3816
rect 536116 3738 536144 55186
rect 536300 3806 536328 59706
rect 537482 59664 537538 59673
rect 537482 59599 537538 59608
rect 541622 59664 541678 59673
rect 541622 59599 541678 59608
rect 537208 4956 537260 4962
rect 537208 4898 537260 4904
rect 536288 3800 536340 3806
rect 536288 3742 536340 3748
rect 536104 3732 536156 3738
rect 536104 3674 536156 3680
rect 536104 3528 536156 3534
rect 536104 3470 536156 3476
rect 536116 480 536144 3470
rect 537220 480 537248 4898
rect 537496 3670 537524 59599
rect 538678 59528 538734 59537
rect 538734 59486 538996 59514
rect 538678 59463 538734 59472
rect 538862 59392 538918 59401
rect 538968 59378 538996 59486
rect 539046 59392 539102 59401
rect 538968 59350 539046 59378
rect 538862 59327 538918 59336
rect 539046 59327 539102 59336
rect 540242 59392 540298 59401
rect 540242 59327 540298 59336
rect 538220 35284 538272 35290
rect 538220 35226 538272 35232
rect 537484 3664 537536 3670
rect 537484 3606 537536 3612
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 35226
rect 538876 3534 538904 59327
rect 538864 3528 538916 3534
rect 538864 3470 538916 3476
rect 540256 3466 540284 59327
rect 540980 47728 541032 47734
rect 540980 47670 541032 47676
rect 540992 16574 541020 47670
rect 540992 16546 541572 16574
rect 540796 4888 540848 4894
rect 540796 4830 540848 4836
rect 539600 3460 539652 3466
rect 539600 3402 539652 3408
rect 540244 3460 540296 3466
rect 540244 3402 540296 3408
rect 539612 480 539640 3402
rect 540808 480 540836 4830
rect 541544 3482 541572 16546
rect 541636 3602 541664 59599
rect 542266 59528 542322 59537
rect 542266 59463 542322 59472
rect 542280 59430 542308 59463
rect 542268 59424 542320 59430
rect 542268 59366 542320 59372
rect 582380 59424 582432 59430
rect 582380 59366 582432 59372
rect 547880 55888 547932 55894
rect 547880 55830 547932 55836
rect 545120 36644 545172 36650
rect 545120 36586 545172 36592
rect 545132 16574 545160 36586
rect 545132 16546 545528 16574
rect 544384 4820 544436 4826
rect 544384 4762 544436 4768
rect 541624 3596 541676 3602
rect 541624 3538 541676 3544
rect 541544 3454 542032 3482
rect 542004 480 542032 3454
rect 543188 3324 543240 3330
rect 543188 3266 543240 3272
rect 543200 480 543228 3266
rect 544396 480 544424 4762
rect 545500 480 545528 16546
rect 546684 3392 546736 3398
rect 546684 3334 546736 3340
rect 546696 480 546724 3334
rect 547892 480 547920 55830
rect 557540 54528 557592 54534
rect 557540 54470 557592 54476
rect 554780 31068 554832 31074
rect 554780 31010 554832 31016
rect 550640 29708 550692 29714
rect 550640 29650 550692 29656
rect 550652 16574 550680 29650
rect 550652 16546 551048 16574
rect 549076 8152 549128 8158
rect 549076 8094 549128 8100
rect 549088 480 549116 8094
rect 550272 4140 550324 4146
rect 550272 4082 550324 4088
rect 550284 480 550312 4082
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 552664 8084 552716 8090
rect 552664 8026 552716 8032
rect 552676 480 552704 8026
rect 553768 4072 553820 4078
rect 553768 4014 553820 4020
rect 553780 480 553808 4014
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 31010
rect 557552 16574 557580 54470
rect 561680 53100 561732 53106
rect 561680 53042 561732 53048
rect 561692 16574 561720 53042
rect 572720 51740 572772 51746
rect 572720 51682 572772 51688
rect 568580 33788 568632 33794
rect 568580 33730 568632 33736
rect 564532 32428 564584 32434
rect 564532 32370 564584 32376
rect 564544 16574 564572 32370
rect 568592 16574 568620 33730
rect 557552 16546 558592 16574
rect 561692 16546 562088 16574
rect 564544 16546 565216 16574
rect 568592 16546 568712 16574
rect 556160 8016 556212 8022
rect 556160 7958 556212 7964
rect 556172 480 556200 7958
rect 557356 4004 557408 4010
rect 557356 3946 557408 3952
rect 557368 480 557396 3946
rect 558564 480 558592 16546
rect 559748 7948 559800 7954
rect 559748 7890 559800 7896
rect 559760 480 559788 7890
rect 560852 3936 560904 3942
rect 560852 3878 560904 3884
rect 560864 480 560892 3878
rect 562060 480 562088 16546
rect 563244 7880 563296 7886
rect 563244 7822 563296 7828
rect 563256 480 563284 7822
rect 564440 3868 564492 3874
rect 564440 3810 564492 3816
rect 564452 480 564480 3810
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565188 354 565216 16546
rect 566832 7812 566884 7818
rect 566832 7754 566884 7760
rect 566844 480 566872 7754
rect 568028 3800 568080 3806
rect 568028 3742 568080 3748
rect 568040 480 568068 3742
rect 565606 354 565718 480
rect 565188 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 568684 354 568712 16546
rect 570328 7744 570380 7750
rect 570328 7686 570380 7692
rect 570340 480 570368 7686
rect 571524 3732 571576 3738
rect 571524 3674 571576 3680
rect 571536 480 571564 3674
rect 572732 480 572760 51682
rect 575480 50380 575532 50386
rect 575480 50322 575532 50328
rect 575492 16574 575520 50322
rect 582392 16574 582420 59366
rect 575492 16546 575888 16574
rect 582392 16546 583432 16574
rect 573916 7676 573968 7682
rect 573916 7618 573968 7624
rect 573928 480 573956 7618
rect 575112 3664 575164 3670
rect 575112 3606 575164 3612
rect 575124 480 575152 3606
rect 569102 354 569214 480
rect 568684 326 569214 354
rect 569102 -960 569214 326
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 575860 354 575888 16546
rect 577412 7608 577464 7614
rect 577412 7550 577464 7556
rect 577424 480 577452 7550
rect 582196 3596 582248 3602
rect 582196 3538 582248 3544
rect 578608 3528 578660 3534
rect 578608 3470 578660 3476
rect 578620 480 578648 3470
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 581012 480 581040 3402
rect 582208 480 582236 3538
rect 583404 480 583432 16546
rect 576278 354 576390 480
rect 575860 326 576390 354
rect 576278 -960 576390 326
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 57426 559408 57482 559464
rect 6458 3304 6514 3360
rect 57978 59744 58034 59800
rect 65890 59764 65946 59800
rect 65890 59744 65892 59764
rect 65892 59744 65944 59764
rect 65944 59744 65946 59764
rect 67914 59744 67970 59800
rect 68834 59744 68890 59800
rect 69846 59744 69902 59800
rect 58622 59608 58678 59664
rect 62026 59608 62082 59664
rect 61382 59472 61438 59528
rect 59358 59372 59360 59392
rect 59360 59372 59412 59392
rect 59412 59372 59414 59392
rect 59358 59336 59414 59372
rect 63958 59492 64014 59528
rect 63958 59472 63960 59492
rect 63960 59472 64012 59492
rect 64012 59472 64014 59492
rect 62026 59336 62082 59392
rect 62762 59336 62818 59392
rect 65982 59608 66038 59664
rect 65890 59336 65946 59392
rect 66902 59472 66958 59528
rect 68466 59608 68522 59664
rect 67914 59336 67970 59392
rect 68282 59336 68338 59392
rect 71042 59608 71098 59664
rect 74998 59608 75054 59664
rect 68834 59472 68890 59528
rect 69846 59472 69902 59528
rect 69662 59336 69718 59392
rect 71778 59472 71834 59528
rect 75642 59744 75698 59800
rect 85026 59744 85082 59800
rect 85210 59744 85266 59800
rect 87970 59744 88026 59800
rect 92294 59744 92350 59800
rect 94134 59744 94190 59800
rect 75642 59608 75698 59664
rect 77574 59608 77630 59664
rect 75458 59472 75514 59528
rect 72422 59336 72478 59392
rect 73802 59336 73858 59392
rect 74998 59336 75054 59392
rect 75182 59200 75238 59256
rect 76562 59472 76618 59528
rect 77574 59336 77630 59392
rect 78770 59608 78826 59664
rect 79966 59608 80022 59664
rect 84106 59608 84162 59664
rect 78586 59336 78642 59392
rect 81346 59472 81402 59528
rect 82542 59336 82598 59392
rect 85394 59472 85450 59528
rect 86866 59472 86922 59528
rect 85210 59336 85266 59392
rect 89626 59472 89682 59528
rect 88246 59336 88302 59392
rect 89442 59336 89498 59392
rect 91282 59472 91338 59528
rect 90822 59336 90878 59392
rect 92386 59472 92442 59528
rect 93214 59336 93270 59392
rect 97078 59764 97134 59800
rect 97078 59744 97080 59764
rect 97080 59744 97132 59764
rect 97132 59744 97134 59764
rect 98090 59744 98146 59800
rect 97262 59608 97318 59664
rect 95146 59472 95202 59528
rect 96066 59336 96122 59392
rect 100942 59764 100998 59800
rect 100942 59744 100944 59764
rect 100944 59744 100996 59764
rect 100996 59744 100998 59764
rect 107750 59764 107806 59800
rect 107750 59744 107752 59764
rect 107752 59744 107804 59764
rect 107804 59744 107806 59764
rect 110694 59764 110750 59800
rect 110694 59744 110696 59764
rect 110696 59744 110748 59764
rect 110748 59744 110750 59764
rect 115570 59764 115626 59800
rect 115570 59744 115572 59764
rect 115572 59744 115624 59764
rect 115624 59744 115626 59764
rect 119710 59744 119766 59800
rect 98090 59336 98146 59392
rect 98642 59336 98698 59392
rect 101586 59472 101642 59528
rect 104898 59472 104954 59528
rect 101402 59336 101458 59392
rect 100022 59200 100078 59256
rect 102782 59336 102838 59392
rect 103518 59372 103520 59392
rect 103520 59372 103572 59392
rect 103572 59372 103574 59392
rect 103518 59336 103574 59372
rect 104346 59200 104402 59256
rect 104162 59064 104218 59120
rect 108302 59472 108358 59528
rect 107106 59200 107162 59256
rect 111246 59472 111302 59528
rect 109682 59336 109738 59392
rect 111062 59336 111118 59392
rect 112442 59336 112498 59392
rect 113270 59336 113326 59392
rect 117502 59608 117558 59664
rect 114650 59492 114706 59528
rect 114650 59472 114652 59492
rect 114652 59472 114704 59492
rect 114704 59472 114706 59492
rect 116582 59472 116638 59528
rect 115202 59336 115258 59392
rect 115754 59336 115810 59392
rect 117502 59336 117558 59392
rect 117962 59336 118018 59392
rect 118698 59608 118754 59664
rect 119434 59608 119490 59664
rect 127254 59764 127310 59800
rect 127254 59744 127256 59764
rect 127256 59744 127308 59764
rect 127308 59744 127310 59764
rect 131118 59764 131174 59800
rect 131118 59744 131120 59764
rect 131120 59744 131172 59764
rect 131172 59744 131174 59764
rect 134062 59764 134118 59800
rect 134062 59744 134064 59764
rect 134064 59744 134116 59764
rect 134116 59744 134118 59764
rect 137006 59764 137062 59800
rect 137006 59744 137008 59764
rect 137008 59744 137060 59764
rect 137060 59744 137062 59764
rect 140870 59744 140926 59800
rect 120906 59472 120962 59528
rect 119710 59336 119766 59392
rect 120722 59336 120778 59392
rect 122746 59336 122802 59392
rect 123022 59336 123078 59392
rect 123298 59200 123354 59256
rect 125322 59628 125378 59664
rect 125322 59608 125324 59628
rect 125324 59608 125376 59628
rect 125376 59608 125378 59628
rect 125322 59472 125378 59528
rect 127806 59472 127862 59528
rect 126242 59336 126298 59392
rect 127622 59336 127678 59392
rect 130474 59200 130530 59256
rect 131946 59472 132002 59528
rect 134522 59472 134578 59528
rect 133142 59336 133198 59392
rect 140042 59608 140098 59664
rect 137282 59472 137338 59528
rect 135902 59336 135958 59392
rect 137466 59336 137522 59392
rect 138662 59200 138718 59256
rect 143814 59764 143870 59800
rect 143814 59744 143816 59764
rect 143816 59744 143868 59764
rect 143868 59744 143870 59764
rect 147678 59764 147734 59800
rect 147678 59744 147680 59764
rect 147680 59744 147732 59764
rect 147732 59744 147734 59764
rect 150622 59764 150678 59800
rect 150622 59744 150624 59764
rect 150624 59744 150676 59764
rect 150676 59744 150678 59764
rect 157430 59764 157486 59800
rect 157430 59744 157432 59764
rect 157432 59744 157484 59764
rect 157484 59744 157486 59764
rect 163318 59764 163374 59800
rect 163318 59744 163320 59764
rect 163320 59744 163372 59764
rect 163372 59744 163374 59764
rect 168286 59744 168342 59800
rect 170126 59744 170182 59800
rect 173990 59744 174046 59800
rect 140870 59336 140926 59392
rect 141606 59472 141662 59528
rect 144366 59472 144422 59528
rect 142802 59336 142858 59392
rect 144182 59336 144238 59392
rect 147034 59200 147090 59256
rect 148506 59472 148562 59528
rect 151266 59472 151322 59528
rect 149702 59336 149758 59392
rect 151082 59336 151138 59392
rect 154486 59492 154542 59528
rect 154486 59472 154488 59492
rect 154488 59472 154540 59492
rect 154540 59472 154542 59492
rect 153842 59200 153898 59256
rect 154026 59064 154082 59120
rect 156602 59608 156658 59664
rect 157982 59472 158038 59528
rect 158166 59336 158222 59392
rect 161294 59628 161350 59664
rect 161294 59608 161296 59628
rect 161296 59608 161348 59628
rect 161348 59608 161350 59628
rect 161294 59472 161350 59528
rect 163502 59472 163558 59528
rect 162122 59336 162178 59392
rect 159362 3304 159418 3360
rect 167182 59492 167238 59528
rect 167182 59472 167184 59492
rect 167184 59472 167236 59492
rect 167236 59472 167238 59492
rect 164882 59336 164938 59392
rect 166446 59336 166502 59392
rect 167642 59200 167698 59256
rect 169114 59608 169170 59664
rect 173162 59608 173218 59664
rect 170586 59472 170642 59528
rect 170126 59336 170182 59392
rect 170402 59336 170458 59392
rect 175094 59472 175150 59528
rect 174910 59336 174966 59392
rect 176934 59744 176990 59800
rect 180798 59764 180854 59800
rect 180798 59744 180800 59764
rect 180800 59744 180852 59764
rect 180852 59744 180854 59764
rect 186594 59764 186650 59800
rect 186594 59744 186596 59764
rect 186596 59744 186648 59764
rect 186648 59744 186650 59764
rect 188342 59744 188398 59800
rect 188618 59744 188674 59800
rect 177762 59472 177818 59528
rect 176382 59336 176438 59392
rect 176566 59336 176622 59392
rect 177946 59336 178002 59392
rect 180706 59472 180762 59528
rect 181810 59472 181866 59528
rect 181994 59336 182050 59392
rect 183466 59200 183522 59256
rect 184570 59064 184626 59120
rect 187330 59608 187386 59664
rect 193034 59608 193090 59664
rect 186226 59336 186282 59392
rect 188986 59472 189042 59528
rect 191470 59472 191526 59528
rect 187514 59200 187570 59256
rect 191654 59336 191710 59392
rect 193770 59608 193826 59664
rect 194598 59744 194654 59800
rect 204166 59764 204222 59800
rect 204166 59744 204168 59764
rect 204168 59744 204220 59764
rect 204220 59744 204222 59764
rect 206742 59744 206798 59800
rect 194598 59608 194654 59664
rect 195886 59608 195942 59664
rect 200302 59608 200358 59664
rect 197266 59472 197322 59528
rect 198554 59336 198610 59392
rect 200026 59336 200082 59392
rect 201314 59472 201370 59528
rect 201314 59336 201370 59392
rect 204166 59608 204222 59664
rect 205546 59472 205602 59528
rect 209962 59744 210018 59800
rect 212906 59764 212962 59800
rect 212906 59744 212908 59764
rect 212908 59744 212960 59764
rect 212960 59744 212962 59764
rect 215850 59744 215906 59800
rect 219530 59744 219586 59800
rect 206926 59336 206982 59392
rect 209686 59336 209742 59392
rect 208214 59200 208270 59256
rect 210790 59200 210846 59256
rect 215206 59608 215262 59664
rect 213550 59472 213606 59528
rect 212446 59200 212502 59256
rect 213734 59200 213790 59256
rect 222658 59764 222714 59800
rect 222658 59744 222660 59764
rect 222660 59744 222712 59764
rect 222712 59744 222714 59764
rect 223670 59744 223726 59800
rect 216586 59472 216642 59528
rect 219530 59472 219586 59528
rect 215850 59336 215906 59392
rect 217874 59336 217930 59392
rect 219346 59336 219402 59392
rect 217690 59200 217746 59256
rect 220818 59608 220874 59664
rect 223486 59608 223542 59664
rect 220726 59472 220782 59528
rect 220818 59336 220874 59392
rect 222106 59336 222162 59392
rect 229466 59764 229522 59800
rect 229466 59744 229468 59764
rect 229468 59744 229520 59764
rect 229520 59744 229522 59764
rect 232410 59764 232466 59800
rect 232410 59744 232412 59764
rect 232412 59744 232464 59764
rect 232464 59744 232466 59764
rect 240138 59764 240194 59800
rect 240138 59744 240140 59764
rect 240140 59744 240192 59764
rect 240192 59744 240194 59764
rect 248970 59764 249026 59800
rect 248970 59744 248972 59764
rect 248972 59744 249024 59764
rect 249024 59744 249026 59764
rect 252834 59764 252890 59800
rect 252834 59744 252836 59764
rect 252836 59744 252888 59764
rect 252888 59744 252890 59764
rect 254306 59744 254362 59800
rect 257986 59744 258042 59800
rect 259642 59744 259698 59800
rect 264794 59744 264850 59800
rect 264978 59744 265034 59800
rect 224774 59472 224830 59528
rect 223670 59336 223726 59392
rect 224590 59336 224646 59392
rect 226522 59472 226578 59528
rect 226062 59336 226118 59392
rect 226246 59336 226302 59392
rect 227350 59200 227406 59256
rect 229006 59336 229062 59392
rect 233146 59608 233202 59664
rect 230294 59200 230350 59256
rect 231766 59200 231822 59256
rect 234250 59472 234306 59528
rect 237378 59492 237434 59528
rect 237378 59472 237380 59492
rect 237380 59472 237432 59492
rect 237432 59472 237434 59492
rect 234434 59336 234490 59392
rect 237010 59200 237066 59256
rect 237286 59064 237342 59120
rect 244094 59628 244150 59664
rect 244094 59608 244096 59628
rect 244096 59608 244148 59628
rect 244148 59608 244150 59628
rect 240046 59472 240102 59528
rect 241426 59472 241482 59528
rect 241242 59336 241298 59392
rect 244094 59472 244150 59528
rect 246026 59492 246082 59528
rect 246026 59472 246028 59492
rect 246028 59472 246080 59492
rect 246080 59472 246082 59492
rect 245566 59336 245622 59392
rect 250902 59608 250958 59664
rect 250810 59472 250866 59528
rect 248326 59336 248382 59392
rect 249706 59336 249762 59392
rect 246854 59200 246910 59256
rect 250902 59336 250958 59392
rect 252466 59336 252522 59392
rect 253754 59336 253810 59392
rect 255226 59608 255282 59664
rect 256606 59472 256662 59528
rect 257710 59336 257766 59392
rect 259366 59608 259422 59664
rect 260746 59472 260802 59528
rect 259642 59336 259698 59392
rect 260654 59336 260710 59392
rect 263506 59608 263562 59664
rect 263506 59472 263562 59528
rect 273258 59764 273314 59800
rect 273258 59744 273260 59764
rect 273260 59744 273312 59764
rect 273312 59744 273314 59764
rect 280066 59764 280122 59800
rect 280066 59744 280068 59764
rect 280068 59744 280120 59764
rect 280120 59744 280122 59764
rect 281078 59744 281134 59800
rect 267646 59608 267702 59664
rect 264978 59472 265034 59528
rect 267462 59472 267518 59528
rect 264886 59336 264942 59392
rect 267554 59336 267610 59392
rect 270314 59628 270370 59664
rect 270314 59608 270316 59628
rect 270316 59608 270368 59628
rect 270368 59608 270370 59628
rect 270314 59472 270370 59528
rect 270130 59200 270186 59256
rect 277122 59628 277178 59664
rect 277122 59608 277124 59628
rect 277124 59608 277176 59628
rect 277176 59608 277178 59628
rect 273166 59472 273222 59528
rect 274454 59472 274510 59528
rect 274270 59336 274326 59392
rect 277306 59472 277362 59528
rect 277122 59336 277178 59392
rect 280066 59608 280122 59664
rect 279882 59200 279938 59256
rect 289818 59764 289874 59800
rect 289818 59744 289820 59764
rect 289820 59744 289872 59764
rect 289872 59744 289874 59764
rect 292762 59764 292818 59800
rect 292762 59744 292764 59764
rect 292764 59744 292816 59764
rect 292816 59744 292818 59764
rect 304998 59744 305054 59800
rect 308954 59744 309010 59800
rect 311990 59744 312046 59800
rect 315762 59764 315818 59800
rect 315762 59744 315764 59764
rect 315764 59744 315816 59764
rect 315816 59744 315818 59764
rect 282826 59608 282882 59664
rect 281446 59472 281502 59528
rect 281078 59336 281134 59392
rect 286874 59628 286930 59664
rect 286874 59608 286876 59628
rect 286876 59608 286928 59628
rect 286928 59608 286930 59628
rect 284114 59472 284170 59528
rect 283930 59336 283986 59392
rect 286874 59472 286930 59528
rect 286874 59336 286930 59392
rect 289082 59200 289138 59256
rect 296626 59628 296682 59664
rect 296626 59608 296628 59628
rect 296628 59608 296680 59628
rect 296680 59608 296682 59628
rect 303618 59608 303674 59664
rect 290646 59472 290702 59528
rect 293222 59472 293278 59528
rect 291842 59336 291898 59392
rect 293406 59336 293462 59392
rect 296626 59472 296682 59528
rect 302238 59472 302294 59528
rect 296166 59200 296222 59256
rect 306378 59336 306434 59392
rect 307942 59336 307998 59392
rect 305274 59200 305330 59256
rect 305090 59064 305146 59120
rect 309138 59472 309194 59528
rect 310518 59336 310574 59392
rect 311898 59336 311954 59392
rect 319626 59744 319682 59800
rect 322570 59764 322626 59800
rect 322570 59744 322572 59764
rect 322572 59744 322624 59764
rect 322624 59744 322626 59764
rect 314842 59472 314898 59528
rect 317418 59472 317474 59528
rect 313278 59336 313334 59392
rect 316130 59336 316186 59392
rect 318798 59608 318854 59664
rect 326158 59744 326214 59800
rect 334346 59764 334402 59800
rect 334346 59744 334348 59764
rect 334348 59744 334400 59764
rect 334400 59744 334402 59764
rect 320454 59608 320510 59664
rect 324502 59628 324558 59664
rect 324502 59608 324504 59628
rect 324504 59608 324556 59628
rect 324556 59608 324558 59628
rect 320270 59472 320326 59528
rect 324502 59472 324558 59528
rect 322938 59336 322994 59392
rect 327262 59608 327318 59664
rect 334162 59608 334218 59664
rect 327078 59336 327134 59392
rect 328550 59472 328606 59528
rect 331402 59472 331458 59528
rect 329930 59336 329986 59392
rect 332598 59336 332654 59392
rect 334254 59336 334310 59392
rect 339130 59764 339186 59800
rect 339130 59744 339132 59764
rect 339132 59744 339184 59764
rect 339184 59744 339186 59764
rect 340878 59744 340934 59800
rect 338302 59472 338358 59528
rect 336738 59200 336794 59256
rect 338486 59336 338542 59392
rect 339498 59336 339554 59392
rect 345386 59744 345442 59800
rect 347686 59744 347742 59800
rect 355598 59764 355654 59800
rect 355598 59744 355600 59764
rect 355600 59744 355652 59764
rect 355652 59744 355654 59764
rect 341154 59472 341210 59528
rect 345018 59336 345074 59392
rect 342258 59200 342314 59256
rect 343822 59200 343878 59256
rect 346490 59472 346546 59528
rect 360382 59744 360438 59800
rect 361486 59744 361542 59800
rect 365350 59764 365406 59800
rect 365350 59744 365352 59764
rect 365352 59744 365404 59764
rect 365404 59744 365406 59764
rect 347870 59608 347926 59664
rect 357622 59608 357678 59664
rect 347778 59472 347834 59528
rect 347686 59336 347742 59392
rect 349158 59472 349214 59528
rect 352746 59492 352802 59528
rect 352746 59472 352748 59492
rect 352748 59472 352800 59492
rect 352800 59472 352802 59492
rect 355322 59472 355378 59528
rect 349342 59336 349398 59392
rect 353942 59336 353998 59392
rect 352562 59200 352618 59256
rect 358082 59472 358138 59528
rect 356702 59336 356758 59392
rect 357622 59336 357678 59392
rect 360474 59472 360530 59528
rect 361026 59472 361082 59528
rect 359462 59336 359518 59392
rect 360382 59336 360438 59392
rect 369306 59764 369362 59800
rect 369306 59744 369308 59764
rect 369308 59744 369360 59764
rect 369360 59744 369362 59764
rect 378046 59744 378102 59800
rect 363326 59608 363382 59664
rect 362222 59472 362278 59528
rect 361486 59336 361542 59392
rect 365166 59472 365222 59528
rect 363602 59336 363658 59392
rect 363786 59336 363842 59392
rect 364982 59336 365038 59392
rect 366362 59200 366418 59256
rect 369122 59472 369178 59528
rect 371146 59472 371202 59528
rect 367926 59200 367982 59256
rect 370502 59200 370558 59256
rect 374090 59628 374146 59664
rect 374090 59608 374092 59628
rect 374092 59608 374144 59628
rect 374144 59608 374146 59628
rect 374090 59472 374146 59528
rect 374090 59336 374146 59392
rect 372158 59200 372214 59256
rect 381910 59780 381912 59800
rect 381912 59780 381964 59800
rect 381964 59780 381966 59800
rect 381910 59744 381966 59780
rect 383290 59780 383292 59800
rect 383292 59780 383344 59800
rect 383344 59780 383346 59800
rect 383290 59744 383346 59780
rect 383842 59744 383898 59800
rect 377586 59472 377642 59528
rect 378414 59472 378470 59528
rect 381542 59472 381598 59528
rect 383842 59472 383898 59528
rect 377402 59336 377458 59392
rect 380162 59336 380218 59392
rect 378598 59200 378654 59256
rect 381726 59336 381782 59392
rect 383014 59336 383070 59392
rect 384854 59744 384910 59800
rect 385958 59764 386014 59800
rect 385958 59744 385960 59764
rect 385960 59744 386012 59764
rect 386012 59744 386014 59764
rect 388718 59764 388774 59800
rect 388718 59744 388720 59764
rect 388720 59744 388772 59764
rect 388772 59744 388774 59764
rect 391662 59764 391718 59800
rect 391662 59744 391664 59764
rect 391664 59744 391716 59764
rect 391716 59744 391718 59764
rect 394606 59744 394662 59800
rect 395710 59764 395766 59800
rect 395710 59744 395712 59764
rect 395712 59744 395764 59764
rect 395764 59744 395766 59764
rect 385682 59608 385738 59664
rect 384854 59336 384910 59392
rect 388442 59472 388498 59528
rect 387062 59336 387118 59392
rect 391202 59472 391258 59528
rect 389822 59336 389878 59392
rect 393594 59472 393650 59528
rect 392674 59336 392730 59392
rect 398470 59764 398526 59800
rect 398470 59744 398472 59764
rect 398472 59744 398524 59764
rect 398524 59744 398526 59764
rect 402426 59764 402482 59800
rect 402426 59744 402428 59764
rect 402428 59744 402480 59764
rect 402480 59744 402482 59764
rect 405278 59764 405334 59800
rect 405278 59744 405280 59764
rect 405280 59744 405332 59764
rect 405332 59744 405334 59764
rect 408406 59744 408462 59800
rect 395342 59608 395398 59664
rect 394606 59336 394662 59392
rect 396722 59336 396778 59392
rect 398286 59472 398342 59528
rect 399390 59336 399446 59392
rect 400862 59336 400918 59392
rect 402334 59608 402390 59664
rect 402242 59472 402298 59528
rect 405002 59472 405058 59528
rect 402334 59336 402390 59392
rect 403622 59336 403678 59392
rect 407762 59472 407818 59528
rect 406382 59336 406438 59392
rect 410154 59764 410210 59800
rect 410154 59744 410156 59764
rect 410156 59744 410208 59764
rect 410208 59744 410210 59764
rect 412086 59744 412142 59800
rect 412454 59744 412510 59800
rect 413098 59764 413154 59800
rect 413098 59744 413100 59764
rect 413100 59744 413152 59764
rect 413152 59744 413154 59764
rect 427450 59744 427506 59800
rect 427634 59744 427690 59800
rect 434442 59744 434498 59800
rect 408682 59608 408738 59664
rect 410154 59608 410210 59664
rect 410522 59472 410578 59528
rect 409142 59336 409198 59392
rect 410154 59336 410210 59392
rect 410706 59336 410762 59392
rect 413926 59608 413982 59664
rect 414018 59472 414074 59528
rect 413098 59336 413154 59392
rect 413926 59336 413982 59392
rect 418158 59608 418214 59664
rect 419814 59628 419870 59664
rect 419814 59608 419816 59628
rect 419816 59608 419868 59628
rect 419868 59608 419870 59628
rect 415030 59472 415086 59528
rect 417054 59472 417110 59528
rect 415398 59336 415454 59392
rect 415582 59336 415638 59392
rect 416870 59336 416926 59392
rect 419538 59472 419594 59528
rect 418986 3304 419042 3360
rect 421838 59472 421894 59528
rect 424782 59472 424838 59528
rect 426530 59472 426586 59528
rect 425058 59336 425114 59392
rect 425242 59336 425298 59392
rect 422390 59200 422446 59256
rect 423954 59200 424010 59256
rect 421286 59064 421342 59120
rect 421838 59064 421894 59120
rect 424138 59064 424194 59120
rect 426714 59336 426770 59392
rect 427450 59336 427506 59392
rect 427910 59608 427966 59664
rect 430578 59472 430634 59528
rect 433522 59472 433578 59528
rect 429198 59200 429254 59256
rect 432050 59336 432106 59392
rect 430670 59200 430726 59256
rect 438030 59764 438086 59800
rect 438030 59744 438032 59764
rect 438032 59744 438084 59764
rect 438084 59744 438086 59764
rect 441986 59744 442042 59800
rect 446402 59744 446458 59800
rect 448150 59744 448206 59800
rect 453946 59744 454002 59800
rect 437570 59608 437626 59664
rect 436190 59472 436246 59528
rect 434718 59336 434774 59392
rect 434902 59336 434958 59392
rect 436374 59336 436430 59392
rect 441066 59608 441122 59664
rect 440514 59336 440570 59392
rect 441066 59336 441122 59392
rect 441618 59336 441674 59392
rect 440330 59064 440386 59120
rect 443090 59608 443146 59664
rect 445758 59472 445814 59528
rect 443274 59336 443330 59392
rect 446954 59608 447010 59664
rect 447138 59608 447194 59664
rect 449990 59472 450046 59528
rect 453026 59472 453082 59528
rect 452842 59336 452898 59392
rect 451278 59200 451334 59256
rect 461582 59764 461638 59800
rect 461582 59744 461584 59764
rect 461584 59744 461636 59764
rect 461636 59744 461638 59764
rect 463606 59744 463662 59800
rect 467562 59744 467618 59800
rect 455878 59608 455934 59664
rect 456890 59628 456946 59664
rect 456890 59608 456892 59628
rect 456892 59608 456944 59628
rect 456944 59608 456946 59628
rect 456614 59472 456670 59528
rect 456890 59472 456946 59528
rect 454038 59336 454094 59392
rect 454222 59336 454278 59392
rect 455510 59336 455566 59392
rect 455878 59336 455934 59392
rect 460938 59608 460994 59664
rect 459834 59472 459890 59528
rect 459650 59336 459706 59392
rect 463698 59472 463754 59528
rect 466642 59472 466698 59528
rect 463882 59336 463938 59392
rect 465078 59336 465134 59392
rect 470598 59764 470654 59800
rect 470598 59744 470600 59764
rect 470600 59744 470652 59764
rect 470652 59744 470654 59764
rect 474370 59764 474426 59800
rect 474370 59744 474372 59764
rect 474372 59744 474424 59764
rect 474424 59744 474426 59764
rect 480258 59764 480314 59800
rect 480258 59744 480260 59764
rect 480260 59744 480312 59764
rect 480312 59744 480314 59764
rect 483294 59744 483350 59800
rect 483478 59744 483534 59800
rect 488446 59744 488502 59800
rect 488630 59744 488686 59800
rect 495898 59764 495954 59800
rect 495898 59744 495900 59764
rect 495900 59744 495952 59764
rect 495952 59744 495954 59764
rect 470552 59608 470608 59664
rect 469310 59472 469366 59528
rect 467838 59336 467894 59392
rect 468022 59336 468078 59392
rect 469494 59336 469550 59392
rect 476302 59608 476358 59664
rect 473634 59472 473690 59528
rect 476210 59472 476266 59528
rect 473450 59336 473506 59392
rect 474738 59336 474794 59392
rect 476302 59336 476358 59392
rect 478326 59608 478382 59664
rect 480258 59608 480314 59664
rect 478878 59472 478934 59528
rect 477590 59336 477646 59392
rect 478326 59336 478382 59392
rect 480350 59200 480406 59256
rect 483110 59472 483166 59528
rect 483294 59336 483350 59392
rect 483294 59200 483350 59256
rect 484398 59608 484454 59664
rect 487066 59608 487122 59664
rect 487250 59472 487306 59528
rect 488446 59472 488502 59528
rect 485962 59336 486018 59392
rect 487066 59336 487122 59392
rect 488538 59336 488594 59392
rect 500682 59764 500738 59800
rect 500682 59744 500684 59764
rect 500684 59744 500736 59764
rect 500736 59744 500738 59764
rect 503626 59764 503682 59800
rect 503626 59744 503628 59764
rect 503628 59744 503680 59764
rect 503680 59744 503682 59764
rect 514298 59744 514354 59800
rect 489918 59608 489974 59664
rect 492862 59628 492918 59664
rect 492862 59608 492864 59628
rect 492864 59608 492916 59628
rect 492916 59608 492918 59628
rect 490010 59472 490066 59528
rect 492954 59472 493010 59528
rect 492770 59336 492826 59392
rect 495530 59336 495586 59392
rect 494150 3576 494206 3632
rect 497738 59492 497794 59528
rect 497738 59472 497740 59492
rect 497740 59472 497792 59492
rect 497792 59472 497794 59492
rect 499854 59472 499910 59528
rect 502430 59472 502486 59528
rect 498382 59336 498438 59392
rect 497094 59200 497150 59256
rect 501050 59336 501106 59392
rect 503626 59608 503682 59664
rect 511998 59608 512054 59664
rect 507490 59492 507546 59528
rect 507490 59472 507492 59492
rect 507492 59472 507544 59492
rect 507544 59472 507546 59492
rect 510618 59472 510674 59528
rect 506754 59200 506810 59256
rect 507950 59200 508006 59256
rect 506570 59064 506626 59120
rect 509606 59336 509662 59392
rect 517242 59764 517298 59800
rect 517242 59744 517244 59764
rect 517244 59744 517296 59764
rect 517296 59744 517298 59764
rect 522118 59764 522174 59800
rect 522118 59744 522120 59764
rect 522120 59744 522172 59764
rect 522172 59744 522174 59764
rect 524050 59764 524106 59800
rect 524050 59744 524052 59764
rect 524052 59744 524104 59764
rect 524104 59744 524106 59764
rect 526994 59764 527050 59800
rect 526994 59744 526996 59764
rect 526996 59744 527048 59764
rect 527048 59744 527050 59764
rect 530858 59764 530914 59800
rect 530858 59744 530860 59764
rect 530860 59744 530912 59764
rect 530912 59744 530914 59764
rect 533802 59764 533858 59800
rect 533802 59744 533804 59764
rect 533804 59744 533856 59764
rect 533856 59744 533858 59764
rect 516322 59472 516378 59528
rect 518990 59472 519046 59528
rect 514758 59336 514814 59392
rect 514942 59336 514998 59392
rect 513654 59200 513710 59256
rect 513470 59064 513526 59120
rect 516506 59336 516562 59392
rect 517518 59336 517574 59392
rect 521658 59472 521714 59528
rect 520370 59336 520426 59392
rect 523130 59200 523186 59256
rect 525062 59336 525118 59392
rect 526626 59472 526682 59528
rect 527822 59200 527878 59256
rect 530766 59472 530822 59528
rect 533342 59472 533398 59528
rect 530582 59336 530638 59392
rect 531962 59336 532018 59392
rect 535734 59472 535790 59528
rect 534722 59336 534778 59392
rect 537482 59608 537538 59664
rect 541622 59608 541678 59664
rect 538678 59472 538734 59528
rect 538862 59336 538918 59392
rect 539046 59336 539102 59392
rect 540242 59336 540298 59392
rect 542266 59472 542322 59528
<< metal3 >>
rect 583520 697084 584960 697324
rect -960 692052 480 692292
rect 583520 683756 584960 683996
rect 583520 670564 584960 670804
rect -960 668524 480 668764
rect 583520 657236 584960 657476
rect -960 645132 480 645372
rect 583520 643908 584960 644148
rect 583520 630716 584960 630956
rect -960 621604 480 621844
rect 583520 617388 584960 617628
rect 583520 604060 584960 604300
rect -960 598212 480 598452
rect 583520 590868 584960 591108
rect 583520 577540 584960 577780
rect -960 574684 480 574924
rect 583520 564212 584960 564452
rect 57421 559466 57487 559469
rect 57421 559464 59554 559466
rect 57421 559408 57426 559464
rect 57482 559430 59554 559464
rect 57482 559408 60076 559430
rect 57421 559406 60076 559408
rect 57421 559403 57487 559406
rect 59494 559370 60076 559406
rect -960 551292 480 551532
rect 583520 551020 584960 551260
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect 583520 511172 584960 511412
rect -960 504372 480 504612
rect 583520 497844 584960 498084
rect 583520 484516 584960 484756
rect -960 480844 480 481084
rect 583520 471324 584960 471564
rect 583520 457996 584960 458236
rect -960 457452 480 457692
rect 583520 444668 584960 444908
rect -960 433924 480 434164
rect 583520 431476 584960 431716
rect 583520 418148 584960 418388
rect -960 410532 480 410772
rect 583520 404820 584960 405060
rect 583520 391628 584960 391868
rect -960 387004 480 387244
rect 583520 378300 584960 378540
rect 583520 364972 584960 365212
rect -960 363612 480 363852
rect 583520 351780 584960 352020
rect -960 340084 480 340324
rect 583520 338452 584960 338692
rect 583520 325124 584960 325364
rect -960 316556 480 316796
rect 583520 311932 584960 312172
rect 583520 298604 584960 298844
rect -960 293164 480 293404
rect 583520 285276 584960 285516
rect 583520 272084 584960 272324
rect -960 269636 480 269876
rect 583520 258756 584960 258996
rect -960 246244 480 246484
rect 583520 245428 584960 245668
rect 583520 232236 584960 232476
rect -960 222716 480 222956
rect 583520 218908 584960 219148
rect 583520 205580 584960 205820
rect -960 199324 480 199564
rect 583520 192388 584960 192628
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 152404 480 152644
rect 583520 152540 584960 152780
rect 583520 139212 584960 139452
rect -960 128876 480 129116
rect 583520 125884 584960 126124
rect 583520 112692 584960 112932
rect -960 105484 480 105724
rect 583520 99364 584960 99604
rect 583520 86036 584960 86276
rect -960 81956 480 82196
rect 583520 72844 584960 73084
rect 57973 59802 58039 59805
rect 60936 59802 60996 60044
rect 57973 59800 60996 59802
rect 57973 59744 57978 59800
rect 58034 59744 60996 59800
rect 57973 59742 60996 59744
rect 57973 59739 58039 59742
rect 58617 59666 58683 59669
rect 61856 59666 61916 60044
rect 58617 59664 61916 59666
rect 58617 59608 58622 59664
rect 58678 59608 61916 59664
rect 58617 59606 61916 59608
rect 62021 59666 62087 59669
rect 62868 59666 62928 60044
rect 62021 59664 62928 59666
rect 62021 59608 62026 59664
rect 62082 59608 62928 59664
rect 62021 59606 62928 59608
rect 58617 59603 58683 59606
rect 62021 59603 62087 59606
rect 61377 59530 61443 59533
rect 63788 59530 63848 60044
rect 61377 59528 63848 59530
rect 61377 59472 61382 59528
rect 61438 59472 63848 59528
rect 61377 59470 63848 59472
rect 63953 59530 64019 59533
rect 64800 59530 64860 60044
rect 63953 59528 64860 59530
rect 63953 59472 63958 59528
rect 64014 59472 64860 59528
rect 63953 59470 64860 59472
rect 61377 59467 61443 59470
rect 63953 59467 64019 59470
rect 59353 59394 59419 59397
rect 62021 59394 62087 59397
rect 59353 59392 62087 59394
rect 59353 59336 59358 59392
rect 59414 59336 62026 59392
rect 62082 59336 62087 59392
rect 59353 59334 62087 59336
rect 59353 59331 59419 59334
rect 62021 59331 62087 59334
rect 62757 59394 62823 59397
rect 65720 59394 65780 60044
rect 65885 59802 65951 59805
rect 66732 59802 66792 60044
rect 65885 59800 66792 59802
rect 65885 59744 65890 59800
rect 65946 59744 66792 59800
rect 65885 59742 66792 59744
rect 65885 59739 65951 59742
rect 65977 59666 66043 59669
rect 67744 59666 67804 60044
rect 67909 59802 67975 59805
rect 68664 59802 68724 60044
rect 67909 59800 68724 59802
rect 67909 59744 67914 59800
rect 67970 59744 68724 59800
rect 67909 59742 68724 59744
rect 68829 59802 68895 59805
rect 69676 59802 69736 60044
rect 70596 59938 70656 60044
rect 71608 59938 71668 60044
rect 70350 59878 70656 59938
rect 70718 59878 71668 59938
rect 68829 59800 69736 59802
rect 68829 59744 68834 59800
rect 68890 59744 69736 59800
rect 68829 59742 69736 59744
rect 69841 59802 69907 59805
rect 70350 59802 70410 59878
rect 69841 59800 70410 59802
rect 69841 59744 69846 59800
rect 69902 59744 70410 59800
rect 69841 59742 70410 59744
rect 67909 59739 67975 59742
rect 68829 59739 68895 59742
rect 69841 59739 69907 59742
rect 65977 59664 67804 59666
rect 65977 59608 65982 59664
rect 66038 59608 67804 59664
rect 65977 59606 67804 59608
rect 68461 59666 68527 59669
rect 70718 59666 70778 59878
rect 72620 59802 72680 60044
rect 68461 59664 70778 59666
rect 68461 59608 68466 59664
rect 68522 59608 70778 59664
rect 68461 59606 70778 59608
rect 70902 59742 72680 59802
rect 65977 59603 66043 59606
rect 68461 59603 68527 59606
rect 66897 59530 66963 59533
rect 68829 59530 68895 59533
rect 69841 59530 69907 59533
rect 66897 59528 68895 59530
rect 66897 59472 66902 59528
rect 66958 59472 68834 59528
rect 68890 59472 68895 59528
rect 66897 59470 68895 59472
rect 66897 59467 66963 59470
rect 68829 59467 68895 59470
rect 69246 59528 69907 59530
rect 69246 59472 69846 59528
rect 69902 59472 69907 59528
rect 69246 59470 69907 59472
rect 62757 59392 65780 59394
rect 62757 59336 62762 59392
rect 62818 59336 65780 59392
rect 62757 59334 65780 59336
rect 65885 59394 65951 59397
rect 67909 59394 67975 59397
rect 65885 59392 67975 59394
rect 65885 59336 65890 59392
rect 65946 59336 67914 59392
rect 67970 59336 67975 59392
rect 65885 59334 67975 59336
rect 62757 59331 62823 59334
rect 65885 59331 65951 59334
rect 67909 59331 67975 59334
rect 68277 59394 68343 59397
rect 69246 59394 69306 59470
rect 69841 59467 69907 59470
rect 68277 59392 69306 59394
rect 68277 59336 68282 59392
rect 68338 59336 69306 59392
rect 68277 59334 69306 59336
rect 69657 59394 69723 59397
rect 70902 59394 70962 59742
rect 71037 59666 71103 59669
rect 73540 59666 73600 60044
rect 71037 59664 73600 59666
rect 71037 59608 71042 59664
rect 71098 59608 73600 59664
rect 71037 59606 73600 59608
rect 71037 59603 71103 59606
rect 71773 59530 71839 59533
rect 74552 59530 74612 60044
rect 74993 59666 75059 59669
rect 75472 59666 75532 60044
rect 75637 59802 75703 59805
rect 76484 59802 76544 60044
rect 75637 59800 76544 59802
rect 75637 59744 75642 59800
rect 75698 59744 76544 59800
rect 75637 59742 76544 59744
rect 75637 59739 75703 59742
rect 74993 59664 75532 59666
rect 74993 59608 74998 59664
rect 75054 59608 75532 59664
rect 74993 59606 75532 59608
rect 75637 59666 75703 59669
rect 77404 59666 77464 60044
rect 75637 59664 77464 59666
rect 75637 59608 75642 59664
rect 75698 59608 77464 59664
rect 75637 59606 77464 59608
rect 77569 59666 77635 59669
rect 78416 59666 78476 60044
rect 79428 59938 79488 60044
rect 80348 59938 80408 60044
rect 77569 59664 78476 59666
rect 77569 59608 77574 59664
rect 77630 59608 78476 59664
rect 77569 59606 78476 59608
rect 78630 59878 79488 59938
rect 79550 59878 80408 59938
rect 74993 59603 75059 59606
rect 75637 59603 75703 59606
rect 77569 59603 77635 59606
rect 75453 59530 75519 59533
rect 71773 59528 74612 59530
rect 71773 59472 71778 59528
rect 71834 59472 74612 59528
rect 71773 59470 74612 59472
rect 74766 59528 75519 59530
rect 74766 59472 75458 59528
rect 75514 59472 75519 59528
rect 74766 59470 75519 59472
rect 71773 59467 71839 59470
rect 69657 59392 70962 59394
rect 69657 59336 69662 59392
rect 69718 59336 70962 59392
rect 69657 59334 70962 59336
rect 72417 59394 72483 59397
rect 73797 59394 73863 59397
rect 74766 59394 74826 59470
rect 75453 59467 75519 59470
rect 76557 59530 76623 59533
rect 78630 59530 78690 59878
rect 78765 59666 78831 59669
rect 79550 59666 79610 59878
rect 81360 59802 81420 60044
rect 78765 59664 79610 59666
rect 78765 59608 78770 59664
rect 78826 59608 79610 59664
rect 78765 59606 79610 59608
rect 79734 59742 81420 59802
rect 78765 59603 78831 59606
rect 76557 59528 78690 59530
rect 76557 59472 76562 59528
rect 76618 59472 78690 59528
rect 76557 59470 78690 59472
rect 76557 59467 76623 59470
rect 74993 59394 75059 59397
rect 77569 59394 77635 59397
rect 72417 59392 73722 59394
rect 72417 59336 72422 59392
rect 72478 59336 73722 59392
rect 72417 59334 73722 59336
rect 68277 59331 68343 59334
rect 69657 59331 69723 59334
rect 72417 59331 72483 59334
rect 73662 59258 73722 59334
rect 73797 59392 74826 59394
rect 73797 59336 73802 59392
rect 73858 59336 74826 59392
rect 73797 59334 74826 59336
rect 74950 59392 75059 59394
rect 74950 59336 74998 59392
rect 75054 59336 75059 59392
rect 73797 59331 73863 59334
rect 74950 59331 75059 59336
rect 75686 59392 77635 59394
rect 75686 59336 77574 59392
rect 77630 59336 77635 59392
rect 75686 59334 77635 59336
rect 74950 59258 75010 59331
rect 73662 59198 75010 59258
rect 75177 59258 75243 59261
rect 75686 59258 75746 59334
rect 77569 59331 77635 59334
rect 78581 59394 78647 59397
rect 79734 59394 79794 59742
rect 79961 59666 80027 59669
rect 82280 59666 82340 60044
rect 79961 59664 82340 59666
rect 79961 59608 79966 59664
rect 80022 59608 82340 59664
rect 79961 59606 82340 59608
rect 79961 59603 80027 59606
rect 81341 59530 81407 59533
rect 83292 59530 83352 60044
rect 84304 59802 84364 60044
rect 85224 59805 85284 60044
rect 85021 59802 85087 59805
rect 84304 59800 85087 59802
rect 84304 59744 85026 59800
rect 85082 59744 85087 59800
rect 84304 59742 85087 59744
rect 85021 59739 85087 59742
rect 85205 59800 85284 59805
rect 85205 59744 85210 59800
rect 85266 59744 85284 59800
rect 85205 59742 85284 59744
rect 85205 59739 85271 59742
rect 84101 59666 84167 59669
rect 86236 59666 86296 60044
rect 87156 59802 87216 60044
rect 87965 59802 88031 59805
rect 87156 59800 88031 59802
rect 87156 59744 87970 59800
rect 88026 59744 88031 59800
rect 87156 59742 88031 59744
rect 87965 59739 88031 59742
rect 88168 59666 88228 60044
rect 84101 59664 86296 59666
rect 84101 59608 84106 59664
rect 84162 59608 86296 59664
rect 84101 59606 86296 59608
rect 86358 59606 88228 59666
rect 84101 59603 84167 59606
rect 81341 59528 83352 59530
rect 81341 59472 81346 59528
rect 81402 59472 83352 59528
rect 81341 59470 83352 59472
rect 85389 59530 85455 59533
rect 86358 59530 86418 59606
rect 85389 59528 86418 59530
rect 85389 59472 85394 59528
rect 85450 59472 86418 59528
rect 85389 59470 86418 59472
rect 86861 59530 86927 59533
rect 89088 59530 89148 60044
rect 90100 59666 90160 60044
rect 86861 59528 89148 59530
rect 86861 59472 86866 59528
rect 86922 59472 89148 59528
rect 86861 59470 89148 59472
rect 89302 59606 90160 59666
rect 81341 59467 81407 59470
rect 85389 59467 85455 59470
rect 86861 59467 86927 59470
rect 78581 59392 79794 59394
rect 78581 59336 78586 59392
rect 78642 59336 79794 59392
rect 78581 59334 79794 59336
rect 82537 59394 82603 59397
rect 85205 59394 85271 59397
rect 82537 59392 85271 59394
rect 82537 59336 82542 59392
rect 82598 59336 85210 59392
rect 85266 59336 85271 59392
rect 82537 59334 85271 59336
rect 78581 59331 78647 59334
rect 82537 59331 82603 59334
rect 85205 59331 85271 59334
rect 88241 59394 88307 59397
rect 89302 59394 89362 59606
rect 89621 59530 89687 59533
rect 91112 59530 91172 60044
rect 89621 59528 91172 59530
rect 89621 59472 89626 59528
rect 89682 59472 91172 59528
rect 89621 59470 91172 59472
rect 91277 59530 91343 59533
rect 92032 59530 92092 60044
rect 93044 59938 93104 60044
rect 92430 59878 93104 59938
rect 92289 59802 92355 59805
rect 92430 59802 92490 59878
rect 92289 59800 92490 59802
rect 92289 59744 92294 59800
rect 92350 59744 92490 59800
rect 92289 59742 92490 59744
rect 92289 59739 92355 59742
rect 91277 59528 92092 59530
rect 91277 59472 91282 59528
rect 91338 59472 92092 59528
rect 91277 59470 92092 59472
rect 92381 59530 92447 59533
rect 93964 59530 94024 60044
rect 94129 59802 94195 59805
rect 94976 59802 95036 60044
rect 94129 59800 95036 59802
rect 94129 59744 94134 59800
rect 94190 59744 95036 59800
rect 94129 59742 95036 59744
rect 94129 59739 94195 59742
rect 95896 59666 95956 60044
rect 92381 59528 94024 59530
rect 92381 59472 92386 59528
rect 92442 59472 94024 59528
rect 92381 59470 94024 59472
rect 94086 59606 95956 59666
rect 89621 59467 89687 59470
rect 91277 59467 91343 59470
rect 92381 59467 92447 59470
rect 88241 59392 89362 59394
rect 88241 59336 88246 59392
rect 88302 59336 89362 59392
rect 88241 59334 89362 59336
rect 89437 59394 89503 59397
rect 90817 59394 90883 59397
rect 89437 59392 90883 59394
rect 89437 59336 89442 59392
rect 89498 59336 90822 59392
rect 90878 59336 90883 59392
rect 89437 59334 90883 59336
rect 88241 59331 88307 59334
rect 89437 59331 89503 59334
rect 90817 59331 90883 59334
rect 93209 59394 93275 59397
rect 94086 59394 94146 59606
rect 95141 59530 95207 59533
rect 96908 59530 96968 60044
rect 97073 59802 97139 59805
rect 97920 59802 97980 60044
rect 97073 59800 97980 59802
rect 97073 59744 97078 59800
rect 97134 59744 97980 59800
rect 97073 59742 97980 59744
rect 98085 59802 98151 59805
rect 98840 59802 98900 60044
rect 98085 59800 98900 59802
rect 98085 59744 98090 59800
rect 98146 59744 98900 59800
rect 98085 59742 98900 59744
rect 97073 59739 97139 59742
rect 98085 59739 98151 59742
rect 97257 59666 97323 59669
rect 97257 59664 99390 59666
rect 97257 59608 97262 59664
rect 97318 59608 99390 59664
rect 97257 59606 99390 59608
rect 97257 59603 97323 59606
rect 95141 59528 96968 59530
rect 95141 59472 95146 59528
rect 95202 59472 96968 59528
rect 95141 59470 96968 59472
rect 99330 59530 99390 59606
rect 99852 59530 99912 60044
rect 99330 59470 99912 59530
rect 95141 59467 95207 59470
rect 93209 59392 94146 59394
rect 93209 59336 93214 59392
rect 93270 59336 94146 59392
rect 93209 59334 94146 59336
rect 96061 59394 96127 59397
rect 98085 59394 98151 59397
rect 96061 59392 98151 59394
rect 96061 59336 96066 59392
rect 96122 59336 98090 59392
rect 98146 59336 98151 59392
rect 96061 59334 98151 59336
rect 93209 59331 93275 59334
rect 96061 59331 96127 59334
rect 98085 59331 98151 59334
rect 98637 59394 98703 59397
rect 100772 59394 100832 60044
rect 100937 59802 101003 59805
rect 101784 59802 101844 60044
rect 100937 59800 101844 59802
rect 100937 59744 100942 59800
rect 100998 59744 101844 59800
rect 100937 59742 101844 59744
rect 100937 59739 101003 59742
rect 102796 59666 102856 60044
rect 98637 59392 100832 59394
rect 98637 59336 98642 59392
rect 98698 59336 100832 59392
rect 98637 59334 100832 59336
rect 100894 59606 102856 59666
rect 98637 59331 98703 59334
rect 75177 59256 75746 59258
rect 75177 59200 75182 59256
rect 75238 59200 75746 59256
rect 75177 59198 75746 59200
rect 100017 59258 100083 59261
rect 100894 59258 100954 59606
rect 101581 59530 101647 59533
rect 103716 59530 103776 60044
rect 101581 59528 103776 59530
rect 101581 59472 101586 59528
rect 101642 59472 103776 59528
rect 101581 59470 103776 59472
rect 101581 59467 101647 59470
rect 101397 59394 101463 59397
rect 102777 59394 102843 59397
rect 103513 59394 103579 59397
rect 104728 59394 104788 60044
rect 104893 59530 104959 59533
rect 105648 59530 105708 60044
rect 104893 59528 105708 59530
rect 104893 59472 104898 59528
rect 104954 59472 105708 59528
rect 104893 59470 105708 59472
rect 104893 59467 104959 59470
rect 106660 59394 106720 60044
rect 107580 59938 107640 60044
rect 101397 59392 102610 59394
rect 101397 59336 101402 59392
rect 101458 59336 102610 59392
rect 101397 59334 102610 59336
rect 101397 59331 101463 59334
rect 100017 59256 100954 59258
rect 100017 59200 100022 59256
rect 100078 59200 100954 59256
rect 100017 59198 100954 59200
rect 102550 59258 102610 59334
rect 102777 59392 103579 59394
rect 102777 59336 102782 59392
rect 102838 59336 103518 59392
rect 103574 59336 103579 59392
rect 102777 59334 103579 59336
rect 102777 59331 102843 59334
rect 103513 59331 103579 59334
rect 103654 59334 104788 59394
rect 104942 59334 106720 59394
rect 106782 59878 107640 59938
rect 103654 59258 103714 59334
rect 102550 59198 103714 59258
rect 104341 59258 104407 59261
rect 104942 59258 105002 59334
rect 104341 59256 105002 59258
rect 104341 59200 104346 59256
rect 104402 59200 105002 59256
rect 104341 59198 105002 59200
rect 75177 59195 75243 59198
rect 100017 59195 100083 59198
rect 104341 59195 104407 59198
rect 104157 59122 104223 59125
rect 106782 59122 106842 59878
rect 107745 59802 107811 59805
rect 108592 59802 108652 60044
rect 107745 59800 108652 59802
rect 107745 59744 107750 59800
rect 107806 59744 108652 59800
rect 107745 59742 108652 59744
rect 107745 59739 107811 59742
rect 109604 59666 109664 60044
rect 107702 59606 109664 59666
rect 107101 59258 107167 59261
rect 107702 59258 107762 59606
rect 108297 59530 108363 59533
rect 110524 59530 110584 60044
rect 110689 59802 110755 59805
rect 111536 59802 111596 60044
rect 110689 59800 111596 59802
rect 110689 59744 110694 59800
rect 110750 59744 111596 59800
rect 110689 59742 111596 59744
rect 110689 59739 110755 59742
rect 112456 59666 112516 60044
rect 108297 59528 110584 59530
rect 108297 59472 108302 59528
rect 108358 59472 110584 59528
rect 108297 59470 110584 59472
rect 110646 59606 112516 59666
rect 108297 59467 108363 59470
rect 109677 59394 109743 59397
rect 110646 59394 110706 59606
rect 111241 59530 111307 59533
rect 113468 59530 113528 60044
rect 111241 59528 113528 59530
rect 111241 59472 111246 59528
rect 111302 59472 113528 59528
rect 111241 59470 113528 59472
rect 111241 59467 111307 59470
rect 109677 59392 110706 59394
rect 109677 59336 109682 59392
rect 109738 59336 110706 59392
rect 109677 59334 110706 59336
rect 111057 59394 111123 59397
rect 112437 59394 112503 59397
rect 113265 59394 113331 59397
rect 114480 59394 114540 60044
rect 114645 59530 114711 59533
rect 115400 59530 115460 60044
rect 115565 59802 115631 59805
rect 116412 59802 116472 60044
rect 115565 59800 116472 59802
rect 115565 59744 115570 59800
rect 115626 59744 116472 59800
rect 115565 59742 116472 59744
rect 115565 59739 115631 59742
rect 117332 59666 117392 60044
rect 114645 59528 115460 59530
rect 114645 59472 114650 59528
rect 114706 59472 115460 59528
rect 114645 59470 115460 59472
rect 115614 59606 117392 59666
rect 117497 59666 117563 59669
rect 118344 59666 118404 60044
rect 119264 59938 119324 60044
rect 120276 59938 120336 60044
rect 117497 59664 118404 59666
rect 117497 59608 117502 59664
rect 117558 59608 118404 59664
rect 117497 59606 118404 59608
rect 118558 59878 119324 59938
rect 119478 59878 120336 59938
rect 114645 59467 114711 59470
rect 111057 59392 112362 59394
rect 111057 59336 111062 59392
rect 111118 59336 112362 59392
rect 111057 59334 112362 59336
rect 109677 59331 109743 59334
rect 111057 59331 111123 59334
rect 107101 59256 107762 59258
rect 107101 59200 107106 59256
rect 107162 59200 107762 59256
rect 107101 59198 107762 59200
rect 112302 59258 112362 59334
rect 112437 59392 113331 59394
rect 112437 59336 112442 59392
rect 112498 59336 113270 59392
rect 113326 59336 113331 59392
rect 112437 59334 113331 59336
rect 112437 59331 112503 59334
rect 113265 59331 113331 59334
rect 113406 59334 114540 59394
rect 115197 59394 115263 59397
rect 115614 59394 115674 59606
rect 117497 59603 117563 59606
rect 116577 59530 116643 59533
rect 118558 59530 118618 59878
rect 119478 59802 119538 59878
rect 119294 59742 119538 59802
rect 119705 59802 119771 59805
rect 121288 59802 121348 60044
rect 119705 59800 121348 59802
rect 119705 59744 119710 59800
rect 119766 59744 121348 59800
rect 119705 59742 121348 59744
rect 118693 59666 118759 59669
rect 119294 59666 119354 59742
rect 119705 59739 119771 59742
rect 118693 59664 119354 59666
rect 118693 59608 118698 59664
rect 118754 59608 119354 59664
rect 118693 59606 119354 59608
rect 119429 59666 119495 59669
rect 122208 59666 122268 60044
rect 119429 59664 122268 59666
rect 119429 59608 119434 59664
rect 119490 59608 122268 59664
rect 119429 59606 122268 59608
rect 118693 59603 118759 59606
rect 119429 59603 119495 59606
rect 116577 59528 118618 59530
rect 116577 59472 116582 59528
rect 116638 59472 118618 59528
rect 116577 59470 118618 59472
rect 120901 59530 120967 59533
rect 123220 59530 123280 60044
rect 120901 59528 123280 59530
rect 120901 59472 120906 59528
rect 120962 59472 123280 59528
rect 120901 59470 123280 59472
rect 116577 59467 116643 59470
rect 120901 59467 120967 59470
rect 115197 59392 115674 59394
rect 115197 59336 115202 59392
rect 115258 59336 115674 59392
rect 115197 59334 115674 59336
rect 115749 59394 115815 59397
rect 117497 59394 117563 59397
rect 115749 59392 117563 59394
rect 115749 59336 115754 59392
rect 115810 59336 117502 59392
rect 117558 59336 117563 59392
rect 115749 59334 117563 59336
rect 113406 59258 113466 59334
rect 115197 59331 115263 59334
rect 115749 59331 115815 59334
rect 117497 59331 117563 59334
rect 117957 59394 118023 59397
rect 119705 59394 119771 59397
rect 117957 59392 119771 59394
rect 117957 59336 117962 59392
rect 118018 59336 119710 59392
rect 119766 59336 119771 59392
rect 117957 59334 119771 59336
rect 117957 59331 118023 59334
rect 119705 59331 119771 59334
rect 120717 59394 120783 59397
rect 122741 59394 122807 59397
rect 123017 59394 123083 59397
rect 124140 59394 124200 60044
rect 125152 59394 125212 60044
rect 125317 59666 125383 59669
rect 126072 59666 126132 60044
rect 125317 59664 126132 59666
rect 125317 59608 125322 59664
rect 125378 59608 126132 59664
rect 125317 59606 126132 59608
rect 125317 59603 125383 59606
rect 125317 59530 125383 59533
rect 127084 59530 127144 60044
rect 127249 59802 127315 59805
rect 128096 59802 128156 60044
rect 127249 59800 128156 59802
rect 127249 59744 127254 59800
rect 127310 59744 128156 59800
rect 127249 59742 128156 59744
rect 127249 59739 127315 59742
rect 129016 59666 129076 60044
rect 125317 59528 127144 59530
rect 125317 59472 125322 59528
rect 125378 59472 127144 59528
rect 125317 59470 127144 59472
rect 127206 59606 129076 59666
rect 125317 59467 125383 59470
rect 120717 59392 122666 59394
rect 120717 59336 120722 59392
rect 120778 59336 122666 59392
rect 120717 59334 122666 59336
rect 120717 59331 120783 59334
rect 112302 59198 113466 59258
rect 122606 59258 122666 59334
rect 122741 59392 123083 59394
rect 122741 59336 122746 59392
rect 122802 59336 123022 59392
rect 123078 59336 123083 59392
rect 122741 59334 123083 59336
rect 122741 59331 122807 59334
rect 123017 59331 123083 59334
rect 123158 59334 124200 59394
rect 124262 59334 125212 59394
rect 126237 59394 126303 59397
rect 127206 59394 127266 59606
rect 127801 59530 127867 59533
rect 130028 59530 130088 60044
rect 130948 59938 131008 60044
rect 130886 59878 131008 59938
rect 130886 59802 130946 59878
rect 127801 59528 130088 59530
rect 127801 59472 127806 59528
rect 127862 59472 130088 59528
rect 127801 59470 130088 59472
rect 130334 59742 130946 59802
rect 131113 59802 131179 59805
rect 131960 59802 132020 60044
rect 131113 59800 132020 59802
rect 131113 59744 131118 59800
rect 131174 59744 132020 59800
rect 131113 59742 132020 59744
rect 127801 59467 127867 59470
rect 126237 59392 127266 59394
rect 126237 59336 126242 59392
rect 126298 59336 127266 59392
rect 126237 59334 127266 59336
rect 127617 59394 127683 59397
rect 127617 59392 128922 59394
rect 127617 59336 127622 59392
rect 127678 59336 128922 59392
rect 127617 59334 128922 59336
rect 123158 59258 123218 59334
rect 122606 59198 123218 59258
rect 123293 59258 123359 59261
rect 124262 59258 124322 59334
rect 126237 59331 126303 59334
rect 127617 59331 127683 59334
rect 123293 59256 124322 59258
rect 123293 59200 123298 59256
rect 123354 59200 124322 59256
rect 123293 59198 124322 59200
rect 128862 59258 128922 59334
rect 130334 59258 130394 59742
rect 131113 59739 131179 59742
rect 132972 59666 133032 60044
rect 131070 59606 133032 59666
rect 128862 59198 130394 59258
rect 130469 59258 130535 59261
rect 131070 59258 131130 59606
rect 131941 59530 132007 59533
rect 133892 59530 133952 60044
rect 134057 59802 134123 59805
rect 134904 59802 134964 60044
rect 134057 59800 134964 59802
rect 134057 59744 134062 59800
rect 134118 59744 134964 59800
rect 134057 59742 134964 59744
rect 134057 59739 134123 59742
rect 135824 59666 135884 60044
rect 131941 59528 133952 59530
rect 131941 59472 131946 59528
rect 132002 59472 133952 59528
rect 131941 59470 133952 59472
rect 134014 59606 135884 59666
rect 131941 59467 132007 59470
rect 133137 59394 133203 59397
rect 134014 59394 134074 59606
rect 134517 59530 134583 59533
rect 136836 59530 136896 60044
rect 137001 59802 137067 59805
rect 137756 59802 137816 60044
rect 137001 59800 137816 59802
rect 137001 59744 137006 59800
rect 137062 59744 137816 59800
rect 137001 59742 137816 59744
rect 137001 59739 137067 59742
rect 138768 59666 138828 60044
rect 134517 59528 136896 59530
rect 134517 59472 134522 59528
rect 134578 59472 136896 59528
rect 134517 59470 136896 59472
rect 136958 59606 138828 59666
rect 134517 59467 134583 59470
rect 133137 59392 134074 59394
rect 133137 59336 133142 59392
rect 133198 59336 134074 59392
rect 133137 59334 134074 59336
rect 135897 59394 135963 59397
rect 136958 59394 137018 59606
rect 137277 59530 137343 59533
rect 139780 59530 139840 60044
rect 140700 59802 140760 60044
rect 137277 59528 139840 59530
rect 137277 59472 137282 59528
rect 137338 59472 139840 59528
rect 137277 59470 139840 59472
rect 139902 59742 140760 59802
rect 140865 59802 140931 59805
rect 141712 59802 141772 60044
rect 140865 59800 141772 59802
rect 140865 59744 140870 59800
rect 140926 59744 141772 59800
rect 140865 59742 141772 59744
rect 137277 59467 137343 59470
rect 135897 59392 137018 59394
rect 135897 59336 135902 59392
rect 135958 59336 137018 59392
rect 135897 59334 137018 59336
rect 137461 59394 137527 59397
rect 139902 59394 139962 59742
rect 140865 59739 140931 59742
rect 140037 59666 140103 59669
rect 142632 59666 142692 60044
rect 140037 59664 142692 59666
rect 140037 59608 140042 59664
rect 140098 59608 142692 59664
rect 140037 59606 142692 59608
rect 140037 59603 140103 59606
rect 141601 59530 141667 59533
rect 143644 59530 143704 60044
rect 143809 59802 143875 59805
rect 144656 59802 144716 60044
rect 143809 59800 144716 59802
rect 143809 59744 143814 59800
rect 143870 59744 144716 59800
rect 143809 59742 144716 59744
rect 143809 59739 143875 59742
rect 145576 59666 145636 60044
rect 141601 59528 143704 59530
rect 141601 59472 141606 59528
rect 141662 59472 143704 59528
rect 141601 59470 143704 59472
rect 143766 59606 145636 59666
rect 141601 59467 141667 59470
rect 140865 59394 140931 59397
rect 137461 59392 139962 59394
rect 137461 59336 137466 59392
rect 137522 59336 139962 59392
rect 137461 59334 139962 59336
rect 140086 59392 140931 59394
rect 140086 59336 140870 59392
rect 140926 59336 140931 59392
rect 140086 59334 140931 59336
rect 133137 59331 133203 59334
rect 135897 59331 135963 59334
rect 137461 59331 137527 59334
rect 130469 59256 131130 59258
rect 130469 59200 130474 59256
rect 130530 59200 131130 59256
rect 130469 59198 131130 59200
rect 138657 59258 138723 59261
rect 140086 59258 140146 59334
rect 140865 59331 140931 59334
rect 142797 59394 142863 59397
rect 143766 59394 143826 59606
rect 144361 59530 144427 59533
rect 146588 59530 146648 60044
rect 147508 59938 147568 60044
rect 147446 59878 147568 59938
rect 147446 59802 147506 59878
rect 144361 59528 146648 59530
rect 144361 59472 144366 59528
rect 144422 59472 146648 59528
rect 144361 59470 146648 59472
rect 146894 59742 147506 59802
rect 147673 59802 147739 59805
rect 148520 59802 148580 60044
rect 147673 59800 148580 59802
rect 147673 59744 147678 59800
rect 147734 59744 148580 59800
rect 147673 59742 148580 59744
rect 144361 59467 144427 59470
rect 142797 59392 143826 59394
rect 142797 59336 142802 59392
rect 142858 59336 143826 59392
rect 142797 59334 143826 59336
rect 144177 59394 144243 59397
rect 144177 59392 145482 59394
rect 144177 59336 144182 59392
rect 144238 59336 145482 59392
rect 144177 59334 145482 59336
rect 142797 59331 142863 59334
rect 144177 59331 144243 59334
rect 138657 59256 140146 59258
rect 138657 59200 138662 59256
rect 138718 59200 140146 59256
rect 138657 59198 140146 59200
rect 145422 59258 145482 59334
rect 146894 59258 146954 59742
rect 147673 59739 147739 59742
rect 149440 59666 149500 60044
rect 147630 59606 149500 59666
rect 145422 59198 146954 59258
rect 147029 59258 147095 59261
rect 147630 59258 147690 59606
rect 148501 59530 148567 59533
rect 150452 59530 150512 60044
rect 150617 59802 150683 59805
rect 151464 59802 151524 60044
rect 150617 59800 151524 59802
rect 150617 59744 150622 59800
rect 150678 59744 151524 59800
rect 150617 59742 151524 59744
rect 150617 59739 150683 59742
rect 152384 59666 152444 60044
rect 148501 59528 150512 59530
rect 148501 59472 148506 59528
rect 148562 59472 150512 59528
rect 148501 59470 150512 59472
rect 150574 59606 152444 59666
rect 148501 59467 148567 59470
rect 149697 59394 149763 59397
rect 150574 59394 150634 59606
rect 151261 59530 151327 59533
rect 153396 59530 153456 60044
rect 151261 59528 153456 59530
rect 151261 59472 151266 59528
rect 151322 59472 153456 59528
rect 151261 59470 153456 59472
rect 151261 59467 151327 59470
rect 149697 59392 150634 59394
rect 149697 59336 149702 59392
rect 149758 59336 150634 59392
rect 149697 59334 150634 59336
rect 151077 59394 151143 59397
rect 154316 59394 154376 60044
rect 154481 59530 154547 59533
rect 155328 59530 155388 60044
rect 154481 59528 155388 59530
rect 154481 59472 154486 59528
rect 154542 59472 155388 59528
rect 154481 59470 155388 59472
rect 154481 59467 154547 59470
rect 156248 59394 156308 60044
rect 157260 59802 157320 60044
rect 151077 59392 154376 59394
rect 151077 59336 151082 59392
rect 151138 59336 154376 59392
rect 151077 59334 154376 59336
rect 154438 59334 156308 59394
rect 156462 59742 157320 59802
rect 157425 59802 157491 59805
rect 158272 59802 158332 60044
rect 157425 59800 158332 59802
rect 157425 59744 157430 59800
rect 157486 59744 158332 59800
rect 157425 59742 158332 59744
rect 149697 59331 149763 59334
rect 151077 59331 151143 59334
rect 147029 59256 147690 59258
rect 147029 59200 147034 59256
rect 147090 59200 147690 59256
rect 147029 59198 147690 59200
rect 153837 59258 153903 59261
rect 154438 59258 154498 59334
rect 153837 59256 154498 59258
rect 153837 59200 153842 59256
rect 153898 59200 154498 59256
rect 153837 59198 154498 59200
rect 107101 59195 107167 59198
rect 123293 59195 123359 59198
rect 130469 59195 130535 59198
rect 138657 59195 138723 59198
rect 147029 59195 147095 59198
rect 153837 59195 153903 59198
rect 104157 59120 106842 59122
rect 104157 59064 104162 59120
rect 104218 59064 106842 59120
rect 104157 59062 106842 59064
rect 154021 59122 154087 59125
rect 156462 59122 156522 59742
rect 157425 59739 157491 59742
rect 156597 59666 156663 59669
rect 159192 59666 159252 60044
rect 156597 59664 159252 59666
rect 156597 59608 156602 59664
rect 156658 59608 159252 59664
rect 156597 59606 159252 59608
rect 156597 59603 156663 59606
rect 157977 59530 158043 59533
rect 160204 59530 160264 60044
rect 157977 59528 160264 59530
rect 157977 59472 157982 59528
rect 158038 59472 160264 59528
rect 157977 59470 160264 59472
rect 157977 59467 158043 59470
rect 158161 59394 158227 59397
rect 161124 59394 161184 60044
rect 161289 59666 161355 59669
rect 162136 59666 162196 60044
rect 161289 59664 162196 59666
rect 161289 59608 161294 59664
rect 161350 59608 162196 59664
rect 161289 59606 162196 59608
rect 161289 59603 161355 59606
rect 161289 59530 161355 59533
rect 163148 59530 163208 60044
rect 163313 59802 163379 59805
rect 164068 59802 164128 60044
rect 163313 59800 164128 59802
rect 163313 59744 163318 59800
rect 163374 59744 164128 59800
rect 163313 59742 164128 59744
rect 163313 59739 163379 59742
rect 165080 59666 165140 60044
rect 161289 59528 163208 59530
rect 161289 59472 161294 59528
rect 161350 59472 163208 59528
rect 161289 59470 163208 59472
rect 163270 59606 165140 59666
rect 161289 59467 161355 59470
rect 158161 59392 161184 59394
rect 158161 59336 158166 59392
rect 158222 59336 161184 59392
rect 158161 59334 161184 59336
rect 162117 59394 162183 59397
rect 163270 59394 163330 59606
rect 163497 59530 163563 59533
rect 166000 59530 166060 60044
rect 167012 59530 167072 60044
rect 163497 59528 166060 59530
rect 163497 59472 163502 59528
rect 163558 59472 166060 59528
rect 163497 59470 166060 59472
rect 166214 59470 167072 59530
rect 167177 59530 167243 59533
rect 167932 59530 167992 60044
rect 168944 59938 169004 60044
rect 167177 59528 167992 59530
rect 167177 59472 167182 59528
rect 167238 59472 167992 59528
rect 167177 59470 167992 59472
rect 168054 59878 169004 59938
rect 163497 59467 163563 59470
rect 162117 59392 163330 59394
rect 162117 59336 162122 59392
rect 162178 59336 163330 59392
rect 162117 59334 163330 59336
rect 164877 59394 164943 59397
rect 166214 59394 166274 59470
rect 167177 59467 167243 59470
rect 164877 59392 166274 59394
rect 164877 59336 164882 59392
rect 164938 59336 166274 59392
rect 164877 59334 166274 59336
rect 166441 59394 166507 59397
rect 168054 59394 168114 59878
rect 168281 59802 168347 59805
rect 169956 59802 170016 60044
rect 168281 59800 170016 59802
rect 168281 59744 168286 59800
rect 168342 59744 170016 59800
rect 168281 59742 170016 59744
rect 170121 59802 170187 59805
rect 170876 59802 170936 60044
rect 170121 59800 170936 59802
rect 170121 59744 170126 59800
rect 170182 59744 170936 59800
rect 170121 59742 170936 59744
rect 168281 59739 168347 59742
rect 170121 59739 170187 59742
rect 169109 59666 169175 59669
rect 171888 59666 171948 60044
rect 169109 59664 171948 59666
rect 169109 59608 169114 59664
rect 169170 59608 171948 59664
rect 169109 59606 171948 59608
rect 169109 59603 169175 59606
rect 170581 59530 170647 59533
rect 172808 59530 172868 60044
rect 173820 59802 173880 60044
rect 170581 59528 172868 59530
rect 170581 59472 170586 59528
rect 170642 59472 172868 59528
rect 170581 59470 172868 59472
rect 173022 59742 173880 59802
rect 173985 59802 174051 59805
rect 174740 59802 174800 60044
rect 173985 59800 174800 59802
rect 173985 59744 173990 59800
rect 174046 59744 174800 59800
rect 173985 59742 174800 59744
rect 170581 59467 170647 59470
rect 170121 59394 170187 59397
rect 166441 59392 168114 59394
rect 166441 59336 166446 59392
rect 166502 59336 168114 59392
rect 166441 59334 168114 59336
rect 169158 59392 170187 59394
rect 169158 59336 170126 59392
rect 170182 59336 170187 59392
rect 169158 59334 170187 59336
rect 158161 59331 158227 59334
rect 162117 59331 162183 59334
rect 164877 59331 164943 59334
rect 166441 59331 166507 59334
rect 167637 59258 167703 59261
rect 169158 59258 169218 59334
rect 170121 59331 170187 59334
rect 170397 59394 170463 59397
rect 173022 59394 173082 59742
rect 173985 59739 174051 59742
rect 173157 59666 173223 59669
rect 175752 59666 175812 60044
rect 173157 59664 175812 59666
rect 173157 59608 173162 59664
rect 173218 59608 175812 59664
rect 173157 59606 175812 59608
rect 173157 59603 173223 59606
rect 175089 59530 175155 59533
rect 176764 59530 176824 60044
rect 176929 59802 176995 59805
rect 177684 59802 177744 60044
rect 176929 59800 177744 59802
rect 176929 59744 176934 59800
rect 176990 59744 177744 59800
rect 176929 59742 177744 59744
rect 176929 59739 176995 59742
rect 178696 59666 178756 60044
rect 175089 59528 176824 59530
rect 175089 59472 175094 59528
rect 175150 59472 176824 59528
rect 175089 59470 176824 59472
rect 177622 59606 178756 59666
rect 175089 59467 175155 59470
rect 170397 59392 173082 59394
rect 170397 59336 170402 59392
rect 170458 59336 173082 59392
rect 170397 59334 173082 59336
rect 174905 59394 174971 59397
rect 176377 59394 176443 59397
rect 174905 59392 176443 59394
rect 174905 59336 174910 59392
rect 174966 59336 176382 59392
rect 176438 59336 176443 59392
rect 174905 59334 176443 59336
rect 170397 59331 170463 59334
rect 174905 59331 174971 59334
rect 176377 59331 176443 59334
rect 176561 59394 176627 59397
rect 177622 59394 177682 59606
rect 177757 59530 177823 59533
rect 179616 59530 179676 60044
rect 180628 59768 180688 60044
rect 177757 59528 179676 59530
rect 177757 59472 177762 59528
rect 177818 59472 179676 59528
rect 177757 59470 179676 59472
rect 180566 59708 180688 59768
rect 180793 59802 180859 59805
rect 181640 59802 181700 60044
rect 180793 59800 181700 59802
rect 180793 59744 180798 59800
rect 180854 59744 181700 59800
rect 180793 59742 181700 59744
rect 180793 59739 180859 59742
rect 177757 59467 177823 59470
rect 176561 59392 177682 59394
rect 176561 59336 176566 59392
rect 176622 59336 177682 59392
rect 176561 59334 177682 59336
rect 177941 59394 178007 59397
rect 180566 59394 180626 59708
rect 182560 59666 182620 60044
rect 180750 59606 182620 59666
rect 180750 59533 180810 59606
rect 180701 59528 180810 59533
rect 180701 59472 180706 59528
rect 180762 59472 180810 59528
rect 180701 59470 180810 59472
rect 181805 59530 181871 59533
rect 183572 59530 183632 60044
rect 181805 59528 183632 59530
rect 181805 59472 181810 59528
rect 181866 59472 183632 59528
rect 181805 59470 183632 59472
rect 180701 59467 180767 59470
rect 181805 59467 181871 59470
rect 177941 59392 179154 59394
rect 177941 59336 177946 59392
rect 178002 59336 179154 59392
rect 177941 59334 179154 59336
rect 176561 59331 176627 59334
rect 177941 59331 178007 59334
rect 167637 59256 169218 59258
rect 167637 59200 167642 59256
rect 167698 59200 169218 59256
rect 167637 59198 169218 59200
rect 179094 59258 179154 59334
rect 180014 59334 180626 59394
rect 181989 59394 182055 59397
rect 184492 59394 184552 60044
rect 185504 59394 185564 60044
rect 186424 59530 186484 60044
rect 186589 59802 186655 59805
rect 187436 59802 187496 60044
rect 188448 59938 188508 60044
rect 188448 59878 188538 59938
rect 188337 59802 188403 59805
rect 186589 59800 187496 59802
rect 186589 59744 186594 59800
rect 186650 59744 187496 59800
rect 186589 59742 187496 59744
rect 187558 59800 188403 59802
rect 187558 59744 188342 59800
rect 188398 59744 188403 59800
rect 187558 59742 188403 59744
rect 186589 59739 186655 59742
rect 187325 59666 187391 59669
rect 187558 59666 187618 59742
rect 188337 59739 188403 59742
rect 188478 59666 188538 59878
rect 188613 59802 188679 59805
rect 189368 59802 189428 60044
rect 188613 59800 189428 59802
rect 188613 59744 188618 59800
rect 188674 59744 189428 59800
rect 188613 59742 189428 59744
rect 188613 59739 188679 59742
rect 190380 59666 190440 60044
rect 187325 59664 187618 59666
rect 187325 59608 187330 59664
rect 187386 59608 187618 59664
rect 187325 59606 187618 59608
rect 188448 59606 188538 59666
rect 188662 59606 190440 59666
rect 187325 59603 187391 59606
rect 181989 59392 184552 59394
rect 181989 59336 181994 59392
rect 182050 59336 184552 59392
rect 181989 59334 184552 59336
rect 184614 59334 185564 59394
rect 185718 59470 186484 59530
rect 180014 59258 180074 59334
rect 181989 59331 182055 59334
rect 179094 59198 180074 59258
rect 183461 59258 183527 59261
rect 184614 59258 184674 59334
rect 183461 59256 184674 59258
rect 183461 59200 183466 59256
rect 183522 59200 184674 59256
rect 183461 59198 184674 59200
rect 167637 59195 167703 59198
rect 183461 59195 183527 59198
rect 154021 59120 156522 59122
rect 154021 59064 154026 59120
rect 154082 59064 156522 59120
rect 154021 59062 156522 59064
rect 184565 59122 184631 59125
rect 185718 59122 185778 59470
rect 186221 59394 186287 59397
rect 188448 59394 188508 59606
rect 186221 59392 188508 59394
rect 186221 59336 186226 59392
rect 186282 59336 188508 59392
rect 186221 59334 188508 59336
rect 186221 59331 186287 59334
rect 187509 59258 187575 59261
rect 188662 59258 188722 59606
rect 188981 59530 189047 59533
rect 191300 59530 191360 60044
rect 192312 59666 192372 60044
rect 193029 59666 193095 59669
rect 192312 59664 193095 59666
rect 192312 59608 193034 59664
rect 193090 59608 193095 59664
rect 192312 59606 193095 59608
rect 193029 59603 193095 59606
rect 188981 59528 191360 59530
rect 188981 59472 188986 59528
rect 189042 59472 191360 59528
rect 188981 59470 191360 59472
rect 191465 59530 191531 59533
rect 193324 59530 193384 60044
rect 194244 59938 194304 60044
rect 195256 59938 195316 60044
rect 196176 59938 196236 60044
rect 191465 59528 193384 59530
rect 191465 59472 191470 59528
rect 191526 59472 193384 59528
rect 191465 59470 193384 59472
rect 193492 59878 194304 59938
rect 194412 59878 195316 59938
rect 195470 59878 196236 59938
rect 188981 59467 189047 59470
rect 191465 59467 191531 59470
rect 191649 59394 191715 59397
rect 193492 59394 193552 59878
rect 194412 59768 194472 59878
rect 194366 59708 194472 59768
rect 194593 59802 194659 59805
rect 195470 59802 195530 59878
rect 197188 59802 197248 60044
rect 194593 59800 195530 59802
rect 194593 59744 194598 59800
rect 194654 59744 195530 59800
rect 194593 59742 195530 59744
rect 195654 59742 197248 59802
rect 194593 59739 194659 59742
rect 193765 59666 193831 59669
rect 194366 59666 194426 59708
rect 193765 59664 194426 59666
rect 193765 59608 193770 59664
rect 193826 59608 194426 59664
rect 193765 59606 194426 59608
rect 194593 59666 194659 59669
rect 195654 59666 195714 59742
rect 194593 59664 195714 59666
rect 194593 59608 194598 59664
rect 194654 59608 195714 59664
rect 194593 59606 195714 59608
rect 195881 59666 195947 59669
rect 198108 59666 198168 60044
rect 195881 59664 198168 59666
rect 195881 59608 195886 59664
rect 195942 59608 198168 59664
rect 195881 59606 198168 59608
rect 193765 59603 193831 59606
rect 194593 59603 194659 59606
rect 195881 59603 195947 59606
rect 197261 59530 197327 59533
rect 199120 59530 199180 60044
rect 200132 59530 200192 60044
rect 200297 59666 200363 59669
rect 201052 59666 201112 60044
rect 202064 59666 202124 60044
rect 200297 59664 201112 59666
rect 200297 59608 200302 59664
rect 200358 59608 201112 59664
rect 200297 59606 201112 59608
rect 201174 59606 202124 59666
rect 200297 59603 200363 59606
rect 197261 59528 199180 59530
rect 197261 59472 197266 59528
rect 197322 59472 199180 59528
rect 197261 59470 199180 59472
rect 199334 59470 200192 59530
rect 197261 59467 197327 59470
rect 191649 59392 193552 59394
rect 191649 59336 191654 59392
rect 191710 59336 193552 59392
rect 191649 59334 193552 59336
rect 198549 59394 198615 59397
rect 199334 59394 199394 59470
rect 198549 59392 199394 59394
rect 198549 59336 198554 59392
rect 198610 59336 199394 59392
rect 198549 59334 199394 59336
rect 200021 59394 200087 59397
rect 201174 59394 201234 59606
rect 201309 59530 201375 59533
rect 202984 59530 203044 60044
rect 201309 59528 203044 59530
rect 201309 59472 201314 59528
rect 201370 59472 203044 59528
rect 201309 59470 203044 59472
rect 201309 59467 201375 59470
rect 200021 59392 201234 59394
rect 200021 59336 200026 59392
rect 200082 59336 201234 59392
rect 200021 59334 201234 59336
rect 201309 59394 201375 59397
rect 203996 59394 204056 60044
rect 204161 59802 204227 59805
rect 204916 59802 204976 60044
rect 204161 59800 204976 59802
rect 204161 59744 204166 59800
rect 204222 59744 204976 59800
rect 204161 59742 204976 59744
rect 205928 59802 205988 60044
rect 206737 59802 206803 59805
rect 205928 59800 206803 59802
rect 205928 59744 206742 59800
rect 206798 59744 206803 59800
rect 205928 59742 206803 59744
rect 204161 59739 204227 59742
rect 206737 59739 206803 59742
rect 204161 59666 204227 59669
rect 206940 59666 207000 60044
rect 204161 59664 207000 59666
rect 204161 59608 204166 59664
rect 204222 59608 207000 59664
rect 204161 59606 207000 59608
rect 204161 59603 204227 59606
rect 205541 59530 205607 59533
rect 207860 59530 207920 60044
rect 205541 59528 207920 59530
rect 205541 59472 205546 59528
rect 205602 59472 207920 59528
rect 205541 59470 207920 59472
rect 205541 59467 205607 59470
rect 201309 59392 204056 59394
rect 201309 59336 201314 59392
rect 201370 59336 204056 59392
rect 201309 59334 204056 59336
rect 206921 59394 206987 59397
rect 208872 59394 208932 60044
rect 209792 59530 209852 60044
rect 209957 59802 210023 59805
rect 210804 59802 210864 60044
rect 209957 59800 210864 59802
rect 209957 59744 209962 59800
rect 210018 59744 210864 59800
rect 209957 59742 210864 59744
rect 209957 59739 210023 59742
rect 206921 59392 208932 59394
rect 206921 59336 206926 59392
rect 206982 59336 208932 59392
rect 206921 59334 208932 59336
rect 209086 59470 209852 59530
rect 191649 59331 191715 59334
rect 198549 59331 198615 59334
rect 200021 59331 200087 59334
rect 201309 59331 201375 59334
rect 206921 59331 206987 59334
rect 187509 59256 188722 59258
rect 187509 59200 187514 59256
rect 187570 59200 188722 59256
rect 187509 59198 188722 59200
rect 208209 59258 208275 59261
rect 209086 59258 209146 59470
rect 209681 59394 209747 59397
rect 211816 59394 211876 60044
rect 212736 59394 212796 60044
rect 213748 59938 213808 60044
rect 214668 59938 214728 60044
rect 212950 59878 213808 59938
rect 213870 59878 214728 59938
rect 212950 59805 213010 59878
rect 212901 59800 213010 59805
rect 212901 59744 212906 59800
rect 212962 59744 213010 59800
rect 212901 59742 213010 59744
rect 212901 59739 212967 59742
rect 213870 59666 213930 59878
rect 215680 59802 215740 60044
rect 214974 59742 215740 59802
rect 215845 59802 215911 59805
rect 216600 59802 216660 60044
rect 215845 59800 216660 59802
rect 215845 59744 215850 59800
rect 215906 59744 216660 59800
rect 215845 59742 216660 59744
rect 214974 59666 215034 59742
rect 215845 59739 215911 59742
rect 209681 59392 211876 59394
rect 209681 59336 209686 59392
rect 209742 59336 211876 59392
rect 209681 59334 211876 59336
rect 212030 59334 212796 59394
rect 212950 59606 213930 59666
rect 214054 59606 215034 59666
rect 215201 59666 215267 59669
rect 217612 59666 217672 60044
rect 215201 59664 217672 59666
rect 215201 59608 215206 59664
rect 215262 59608 217672 59664
rect 215201 59606 217672 59608
rect 209681 59331 209747 59334
rect 208209 59256 209146 59258
rect 208209 59200 208214 59256
rect 208270 59200 209146 59256
rect 208209 59198 209146 59200
rect 210785 59258 210851 59261
rect 212030 59258 212090 59334
rect 210785 59256 212090 59258
rect 210785 59200 210790 59256
rect 210846 59200 212090 59256
rect 210785 59198 212090 59200
rect 212441 59258 212507 59261
rect 212950 59258 213010 59606
rect 213545 59530 213611 59533
rect 214054 59530 214114 59606
rect 215201 59603 215267 59606
rect 213545 59528 214114 59530
rect 213545 59472 213550 59528
rect 213606 59472 214114 59528
rect 213545 59470 214114 59472
rect 216581 59530 216647 59533
rect 218624 59530 218684 60044
rect 219544 59805 219604 60044
rect 219525 59800 219604 59805
rect 219525 59744 219530 59800
rect 219586 59744 219604 59800
rect 219525 59742 219604 59744
rect 219525 59739 219591 59742
rect 220556 59666 220616 60044
rect 216581 59528 218684 59530
rect 216581 59472 216586 59528
rect 216642 59472 218684 59528
rect 216581 59470 218684 59472
rect 218838 59606 220616 59666
rect 220813 59666 220879 59669
rect 221476 59666 221536 60044
rect 220813 59664 221536 59666
rect 220813 59608 220818 59664
rect 220874 59608 221536 59664
rect 220813 59606 221536 59608
rect 213545 59467 213611 59470
rect 216581 59467 216647 59470
rect 215845 59394 215911 59397
rect 214790 59392 215911 59394
rect 214790 59336 215850 59392
rect 215906 59336 215911 59392
rect 214790 59334 215911 59336
rect 212441 59256 213010 59258
rect 212441 59200 212446 59256
rect 212502 59200 213010 59256
rect 212441 59198 213010 59200
rect 213729 59258 213795 59261
rect 214790 59258 214850 59334
rect 215845 59331 215911 59334
rect 217869 59394 217935 59397
rect 218838 59394 218898 59606
rect 220813 59603 220879 59606
rect 219525 59530 219591 59533
rect 217869 59392 218898 59394
rect 217869 59336 217874 59392
rect 217930 59336 218898 59392
rect 217869 59334 218898 59336
rect 219022 59528 219591 59530
rect 219022 59472 219530 59528
rect 219586 59472 219591 59528
rect 219022 59470 219591 59472
rect 217869 59331 217935 59334
rect 213729 59256 214850 59258
rect 213729 59200 213734 59256
rect 213790 59200 214850 59256
rect 213729 59198 214850 59200
rect 217685 59258 217751 59261
rect 219022 59258 219082 59470
rect 219525 59467 219591 59470
rect 220721 59530 220787 59533
rect 222488 59530 222548 60044
rect 222653 59802 222719 59805
rect 223500 59802 223560 60044
rect 222653 59800 223560 59802
rect 222653 59744 222658 59800
rect 222714 59744 223560 59800
rect 222653 59742 223560 59744
rect 223665 59802 223731 59805
rect 224420 59802 224480 60044
rect 223665 59800 224480 59802
rect 223665 59744 223670 59800
rect 223726 59744 224480 59800
rect 223665 59742 224480 59744
rect 222653 59739 222719 59742
rect 223665 59739 223731 59742
rect 223481 59666 223547 59669
rect 225432 59666 225492 60044
rect 223481 59664 225492 59666
rect 223481 59608 223486 59664
rect 223542 59608 225492 59664
rect 223481 59606 225492 59608
rect 223481 59603 223547 59606
rect 220721 59528 222548 59530
rect 220721 59472 220726 59528
rect 220782 59472 222548 59528
rect 220721 59470 222548 59472
rect 224769 59530 224835 59533
rect 226352 59530 226412 60044
rect 224769 59528 226412 59530
rect 224769 59472 224774 59528
rect 224830 59472 226412 59528
rect 224769 59470 226412 59472
rect 226517 59530 226583 59533
rect 227364 59530 227424 60044
rect 226517 59528 227424 59530
rect 226517 59472 226522 59528
rect 226578 59472 227424 59528
rect 226517 59470 227424 59472
rect 220721 59467 220787 59470
rect 224769 59467 224835 59470
rect 226517 59467 226583 59470
rect 219341 59394 219407 59397
rect 220813 59394 220879 59397
rect 219341 59392 220879 59394
rect 219341 59336 219346 59392
rect 219402 59336 220818 59392
rect 220874 59336 220879 59392
rect 219341 59334 220879 59336
rect 219341 59331 219407 59334
rect 220813 59331 220879 59334
rect 222101 59394 222167 59397
rect 223665 59394 223731 59397
rect 222101 59392 223731 59394
rect 222101 59336 222106 59392
rect 222162 59336 223670 59392
rect 223726 59336 223731 59392
rect 222101 59334 223731 59336
rect 222101 59331 222167 59334
rect 223665 59331 223731 59334
rect 224585 59394 224651 59397
rect 226057 59394 226123 59397
rect 224585 59392 226123 59394
rect 224585 59336 224590 59392
rect 224646 59336 226062 59392
rect 226118 59336 226123 59392
rect 224585 59334 226123 59336
rect 224585 59331 224651 59334
rect 226057 59331 226123 59334
rect 226241 59394 226307 59397
rect 228284 59394 228344 60044
rect 229296 59530 229356 60044
rect 229461 59802 229527 59805
rect 230308 59802 230368 60044
rect 229461 59800 230368 59802
rect 229461 59744 229466 59800
rect 229522 59744 230368 59800
rect 229461 59742 230368 59744
rect 229461 59739 229527 59742
rect 226241 59392 228344 59394
rect 226241 59336 226246 59392
rect 226302 59336 228344 59392
rect 226241 59334 228344 59336
rect 228406 59470 229356 59530
rect 226241 59331 226307 59334
rect 217685 59256 219082 59258
rect 217685 59200 217690 59256
rect 217746 59200 219082 59256
rect 217685 59198 219082 59200
rect 227345 59258 227411 59261
rect 228406 59258 228466 59470
rect 229001 59394 229067 59397
rect 231228 59394 231288 60044
rect 232240 59938 232300 60044
rect 233160 59938 233220 60044
rect 232086 59878 232300 59938
rect 232454 59878 233220 59938
rect 232086 59666 232146 59878
rect 232454 59805 232514 59878
rect 232405 59800 232514 59805
rect 234172 59802 234232 60044
rect 232405 59744 232410 59800
rect 232466 59744 232514 59800
rect 232405 59742 232514 59744
rect 232638 59742 234232 59802
rect 232405 59739 232471 59742
rect 232086 59606 232300 59666
rect 232240 59394 232300 59606
rect 232638 59394 232698 59742
rect 233141 59666 233207 59669
rect 235092 59666 235152 60044
rect 233141 59664 235152 59666
rect 233141 59608 233146 59664
rect 233202 59608 235152 59664
rect 233141 59606 235152 59608
rect 233141 59603 233207 59606
rect 234245 59530 234311 59533
rect 236104 59530 236164 60044
rect 234245 59528 236164 59530
rect 234245 59472 234250 59528
rect 234306 59472 236164 59528
rect 234245 59470 236164 59472
rect 234245 59467 234311 59470
rect 229001 59392 231288 59394
rect 229001 59336 229006 59392
rect 229062 59336 231288 59392
rect 229001 59334 231288 59336
rect 231350 59334 232300 59394
rect 232454 59334 232698 59394
rect 234429 59394 234495 59397
rect 237116 59394 237176 60044
rect 237373 59530 237439 59533
rect 238036 59530 238096 60044
rect 237373 59528 238096 59530
rect 237373 59472 237378 59528
rect 237434 59472 238096 59528
rect 237373 59470 238096 59472
rect 237373 59467 237439 59470
rect 239048 59394 239108 60044
rect 239968 59666 240028 60044
rect 240133 59802 240199 59805
rect 240980 59802 241040 60044
rect 240133 59800 241040 59802
rect 240133 59744 240138 59800
rect 240194 59744 241040 59800
rect 240133 59742 241040 59744
rect 240133 59739 240199 59742
rect 241992 59666 242052 60044
rect 234429 59392 237176 59394
rect 234429 59336 234434 59392
rect 234490 59336 237176 59392
rect 234429 59334 237176 59336
rect 237238 59334 239108 59394
rect 239262 59606 240028 59666
rect 240182 59606 242052 59666
rect 229001 59331 229067 59334
rect 227345 59256 228466 59258
rect 227345 59200 227350 59256
rect 227406 59200 228466 59256
rect 227345 59198 228466 59200
rect 230289 59258 230355 59261
rect 231350 59258 231410 59334
rect 230289 59256 231410 59258
rect 230289 59200 230294 59256
rect 230350 59200 231410 59256
rect 230289 59198 231410 59200
rect 231761 59258 231827 59261
rect 232454 59258 232514 59334
rect 234429 59331 234495 59334
rect 231761 59256 232514 59258
rect 231761 59200 231766 59256
rect 231822 59200 232514 59256
rect 231761 59198 232514 59200
rect 237005 59258 237071 59261
rect 237238 59258 237298 59334
rect 237005 59256 237298 59258
rect 237005 59200 237010 59256
rect 237066 59200 237298 59256
rect 237005 59198 237298 59200
rect 187509 59195 187575 59198
rect 208209 59195 208275 59198
rect 210785 59195 210851 59198
rect 212441 59195 212507 59198
rect 213729 59195 213795 59198
rect 217685 59195 217751 59198
rect 227345 59195 227411 59198
rect 230289 59195 230355 59198
rect 231761 59195 231827 59198
rect 237005 59195 237071 59198
rect 184565 59120 185778 59122
rect 184565 59064 184570 59120
rect 184626 59064 185778 59120
rect 184565 59062 185778 59064
rect 237281 59122 237347 59125
rect 239262 59122 239322 59606
rect 240041 59530 240107 59533
rect 240182 59530 240242 59606
rect 240041 59528 240242 59530
rect 240041 59472 240046 59528
rect 240102 59472 240242 59528
rect 240041 59470 240242 59472
rect 241421 59530 241487 59533
rect 242912 59530 242972 60044
rect 241421 59528 242972 59530
rect 241421 59472 241426 59528
rect 241482 59472 242972 59528
rect 241421 59470 242972 59472
rect 240041 59467 240107 59470
rect 241421 59467 241487 59470
rect 241237 59394 241303 59397
rect 243924 59394 243984 60044
rect 244089 59666 244155 59669
rect 244844 59666 244904 60044
rect 244089 59664 244904 59666
rect 244089 59608 244094 59664
rect 244150 59608 244904 59664
rect 244089 59606 244904 59608
rect 244089 59603 244155 59606
rect 244089 59530 244155 59533
rect 245856 59530 245916 60044
rect 244089 59528 245916 59530
rect 244089 59472 244094 59528
rect 244150 59472 245916 59528
rect 244089 59470 245916 59472
rect 246021 59530 246087 59533
rect 246776 59530 246836 60044
rect 246021 59528 246836 59530
rect 246021 59472 246026 59528
rect 246082 59472 246836 59528
rect 246021 59470 246836 59472
rect 244089 59467 244155 59470
rect 246021 59467 246087 59470
rect 241237 59392 243984 59394
rect 241237 59336 241242 59392
rect 241298 59336 243984 59392
rect 241237 59334 243984 59336
rect 245561 59394 245627 59397
rect 247788 59394 247848 60044
rect 248800 59530 248860 60044
rect 248965 59802 249031 59805
rect 249720 59802 249780 60044
rect 248965 59800 249780 59802
rect 248965 59744 248970 59800
rect 249026 59744 249780 59800
rect 248965 59742 249780 59744
rect 248965 59739 249031 59742
rect 250732 59666 250792 60044
rect 245561 59392 247848 59394
rect 245561 59336 245566 59392
rect 245622 59336 247848 59392
rect 245561 59334 247848 59336
rect 247910 59470 248860 59530
rect 249566 59606 250792 59666
rect 250897 59666 250963 59669
rect 251652 59666 251712 60044
rect 250897 59664 251712 59666
rect 250897 59608 250902 59664
rect 250958 59608 251712 59664
rect 250897 59606 251712 59608
rect 241237 59331 241303 59334
rect 245561 59331 245627 59334
rect 246849 59258 246915 59261
rect 247910 59258 247970 59470
rect 248321 59394 248387 59397
rect 249566 59394 249626 59606
rect 250897 59603 250963 59606
rect 250805 59530 250871 59533
rect 252664 59530 252724 60044
rect 253676 59938 253736 60044
rect 254596 59938 254656 60044
rect 255608 59938 255668 60044
rect 252878 59878 253736 59938
rect 253982 59878 254656 59938
rect 254718 59878 255668 59938
rect 252878 59805 252938 59878
rect 252829 59800 252938 59805
rect 252829 59744 252834 59800
rect 252890 59744 252938 59800
rect 252829 59742 252938 59744
rect 252829 59739 252895 59742
rect 253982 59530 254042 59878
rect 254301 59802 254367 59805
rect 254718 59802 254778 59878
rect 256528 59802 256588 60044
rect 254301 59800 254778 59802
rect 254301 59744 254306 59800
rect 254362 59744 254778 59800
rect 254301 59742 254778 59744
rect 255086 59742 256588 59802
rect 254301 59739 254367 59742
rect 250805 59528 252724 59530
rect 250805 59472 250810 59528
rect 250866 59472 252724 59528
rect 250805 59470 252724 59472
rect 252832 59470 254042 59530
rect 250805 59467 250871 59470
rect 248321 59392 249626 59394
rect 248321 59336 248326 59392
rect 248382 59336 249626 59392
rect 248321 59334 249626 59336
rect 249701 59394 249767 59397
rect 250897 59394 250963 59397
rect 249701 59392 250963 59394
rect 249701 59336 249706 59392
rect 249762 59336 250902 59392
rect 250958 59336 250963 59392
rect 249701 59334 250963 59336
rect 248321 59331 248387 59334
rect 249701 59331 249767 59334
rect 250897 59331 250963 59334
rect 252461 59394 252527 59397
rect 252832 59394 252892 59470
rect 252461 59392 252892 59394
rect 252461 59336 252466 59392
rect 252522 59336 252892 59392
rect 252461 59334 252892 59336
rect 253749 59394 253815 59397
rect 255086 59394 255146 59742
rect 255221 59666 255287 59669
rect 257540 59666 257600 60044
rect 258460 59938 258520 60044
rect 255221 59664 257600 59666
rect 255221 59608 255226 59664
rect 255282 59608 257600 59664
rect 255221 59606 257600 59608
rect 257662 59878 258520 59938
rect 255221 59603 255287 59606
rect 256601 59530 256667 59533
rect 257662 59530 257722 59878
rect 257981 59802 258047 59805
rect 259472 59802 259532 60044
rect 257981 59800 259532 59802
rect 257981 59744 257986 59800
rect 258042 59744 259532 59800
rect 257981 59742 259532 59744
rect 259637 59802 259703 59805
rect 260484 59802 260544 60044
rect 259637 59800 260544 59802
rect 259637 59744 259642 59800
rect 259698 59744 260544 59800
rect 259637 59742 260544 59744
rect 257981 59739 258047 59742
rect 259637 59739 259703 59742
rect 259361 59666 259427 59669
rect 261404 59666 261464 60044
rect 259361 59664 261464 59666
rect 259361 59608 259366 59664
rect 259422 59608 261464 59664
rect 259361 59606 261464 59608
rect 259361 59603 259427 59606
rect 256601 59528 257722 59530
rect 256601 59472 256606 59528
rect 256662 59472 257722 59528
rect 256601 59470 257722 59472
rect 260741 59530 260807 59533
rect 262416 59530 262476 60044
rect 260741 59528 262476 59530
rect 260741 59472 260746 59528
rect 260802 59472 262476 59528
rect 260741 59470 262476 59472
rect 256601 59467 256667 59470
rect 260741 59467 260807 59470
rect 253749 59392 255146 59394
rect 253749 59336 253754 59392
rect 253810 59336 255146 59392
rect 253749 59334 255146 59336
rect 257705 59394 257771 59397
rect 259637 59394 259703 59397
rect 257705 59392 259703 59394
rect 257705 59336 257710 59392
rect 257766 59336 259642 59392
rect 259698 59336 259703 59392
rect 257705 59334 259703 59336
rect 252461 59331 252527 59334
rect 253749 59331 253815 59334
rect 257705 59331 257771 59334
rect 259637 59331 259703 59334
rect 260649 59394 260715 59397
rect 263336 59394 263396 60044
rect 264348 59802 264408 60044
rect 264789 59802 264855 59805
rect 264348 59800 264855 59802
rect 264348 59744 264794 59800
rect 264850 59744 264855 59800
rect 264348 59742 264855 59744
rect 264789 59739 264855 59742
rect 264973 59802 265039 59805
rect 265268 59802 265328 60044
rect 264973 59800 265328 59802
rect 264973 59744 264978 59800
rect 265034 59744 265328 59800
rect 264973 59742 265328 59744
rect 264973 59739 265039 59742
rect 263501 59666 263567 59669
rect 266280 59666 266340 60044
rect 263501 59664 266340 59666
rect 263501 59608 263506 59664
rect 263562 59608 266340 59664
rect 263501 59606 266340 59608
rect 263501 59603 263567 59606
rect 263501 59530 263567 59533
rect 264973 59530 265039 59533
rect 263501 59528 265039 59530
rect 263501 59472 263506 59528
rect 263562 59472 264978 59528
rect 265034 59472 265039 59528
rect 263501 59470 265039 59472
rect 263501 59467 263567 59470
rect 264973 59467 265039 59470
rect 260649 59392 263396 59394
rect 260649 59336 260654 59392
rect 260710 59336 263396 59392
rect 260649 59334 263396 59336
rect 264881 59394 264947 59397
rect 267292 59394 267352 60044
rect 267641 59666 267707 59669
rect 268212 59666 268272 60044
rect 267641 59664 268272 59666
rect 267641 59608 267646 59664
rect 267702 59608 268272 59664
rect 267641 59606 268272 59608
rect 267641 59603 267707 59606
rect 267457 59530 267523 59533
rect 269224 59530 269284 60044
rect 267457 59528 269284 59530
rect 267457 59472 267462 59528
rect 267518 59472 269284 59528
rect 267457 59470 269284 59472
rect 267457 59467 267523 59470
rect 264881 59392 267352 59394
rect 264881 59336 264886 59392
rect 264942 59336 267352 59392
rect 264881 59334 267352 59336
rect 267549 59394 267615 59397
rect 270144 59394 270204 60044
rect 270309 59666 270375 59669
rect 271156 59666 271216 60044
rect 270309 59664 271216 59666
rect 270309 59608 270314 59664
rect 270370 59608 271216 59664
rect 270309 59606 271216 59608
rect 270309 59603 270375 59606
rect 270309 59530 270375 59533
rect 272168 59530 272228 60044
rect 273088 59666 273148 60044
rect 273253 59802 273319 59805
rect 274100 59802 274160 60044
rect 273253 59800 274160 59802
rect 273253 59744 273258 59800
rect 273314 59744 274160 59800
rect 273253 59742 274160 59744
rect 273253 59739 273319 59742
rect 275020 59666 275080 60044
rect 270309 59528 272228 59530
rect 270309 59472 270314 59528
rect 270370 59472 272228 59528
rect 270309 59470 272228 59472
rect 272566 59606 273148 59666
rect 273302 59606 275080 59666
rect 270309 59467 270375 59470
rect 267549 59392 270204 59394
rect 267549 59336 267554 59392
rect 267610 59336 270204 59392
rect 267549 59334 270204 59336
rect 270358 59334 271706 59394
rect 260649 59331 260715 59334
rect 264881 59331 264947 59334
rect 267549 59331 267615 59334
rect 246849 59256 247970 59258
rect 246849 59200 246854 59256
rect 246910 59200 247970 59256
rect 246849 59198 247970 59200
rect 270125 59258 270191 59261
rect 270358 59258 270418 59334
rect 270125 59256 270418 59258
rect 270125 59200 270130 59256
rect 270186 59200 270418 59256
rect 270125 59198 270418 59200
rect 271646 59258 271706 59334
rect 272566 59258 272626 59606
rect 273161 59530 273227 59533
rect 273302 59530 273362 59606
rect 273161 59528 273362 59530
rect 273161 59472 273166 59528
rect 273222 59472 273362 59528
rect 273161 59470 273362 59472
rect 274449 59530 274515 59533
rect 276032 59530 276092 60044
rect 274449 59528 276092 59530
rect 274449 59472 274454 59528
rect 274510 59472 276092 59528
rect 274449 59470 276092 59472
rect 273161 59467 273227 59470
rect 274449 59467 274515 59470
rect 274265 59394 274331 59397
rect 276952 59394 277012 60044
rect 277117 59666 277183 59669
rect 277964 59666 278024 60044
rect 277117 59664 278024 59666
rect 277117 59608 277122 59664
rect 277178 59608 278024 59664
rect 277117 59606 278024 59608
rect 277117 59603 277183 59606
rect 277301 59530 277367 59533
rect 278976 59530 279036 60044
rect 277301 59528 279036 59530
rect 277301 59472 277306 59528
rect 277362 59472 279036 59528
rect 277301 59470 279036 59472
rect 277301 59467 277367 59470
rect 274265 59392 277012 59394
rect 274265 59336 274270 59392
rect 274326 59336 277012 59392
rect 274265 59334 277012 59336
rect 277117 59394 277183 59397
rect 279896 59394 279956 60044
rect 280061 59802 280127 59805
rect 280908 59802 280968 60044
rect 280061 59800 280968 59802
rect 280061 59744 280066 59800
rect 280122 59744 280968 59800
rect 280061 59742 280968 59744
rect 281073 59802 281139 59805
rect 281828 59802 281888 60044
rect 282840 59938 282900 60044
rect 281073 59800 281888 59802
rect 281073 59744 281078 59800
rect 281134 59744 281888 59800
rect 281073 59742 281888 59744
rect 281950 59878 282900 59938
rect 280061 59739 280127 59742
rect 281073 59739 281139 59742
rect 280061 59666 280127 59669
rect 281950 59666 282010 59878
rect 283852 59802 283912 60044
rect 280061 59664 282010 59666
rect 280061 59608 280066 59664
rect 280122 59608 282010 59664
rect 280061 59606 282010 59608
rect 282134 59742 283912 59802
rect 280061 59603 280127 59606
rect 281441 59530 281507 59533
rect 282134 59530 282194 59742
rect 282821 59666 282887 59669
rect 284772 59666 284832 60044
rect 282821 59664 284832 59666
rect 282821 59608 282826 59664
rect 282882 59608 284832 59664
rect 282821 59606 284832 59608
rect 282821 59603 282887 59606
rect 281441 59528 282194 59530
rect 281441 59472 281446 59528
rect 281502 59472 282194 59528
rect 281441 59470 282194 59472
rect 284109 59530 284175 59533
rect 285784 59530 285844 60044
rect 284109 59528 285844 59530
rect 284109 59472 284114 59528
rect 284170 59472 285844 59528
rect 284109 59470 285844 59472
rect 281441 59467 281507 59470
rect 284109 59467 284175 59470
rect 281073 59394 281139 59397
rect 277117 59392 279956 59394
rect 277117 59336 277122 59392
rect 277178 59336 279956 59392
rect 277117 59334 279956 59336
rect 280110 59392 281139 59394
rect 280110 59336 281078 59392
rect 281134 59336 281139 59392
rect 280110 59334 281139 59336
rect 274265 59331 274331 59334
rect 277117 59331 277183 59334
rect 271646 59198 272626 59258
rect 279877 59258 279943 59261
rect 280110 59258 280170 59334
rect 281073 59331 281139 59334
rect 283925 59394 283991 59397
rect 286704 59394 286764 60044
rect 286869 59666 286935 59669
rect 287716 59666 287776 60044
rect 286869 59664 287776 59666
rect 286869 59608 286874 59664
rect 286930 59608 287776 59664
rect 286869 59606 287776 59608
rect 286869 59603 286935 59606
rect 286869 59530 286935 59533
rect 288636 59530 288696 60044
rect 286869 59528 288696 59530
rect 286869 59472 286874 59528
rect 286930 59472 288696 59528
rect 286869 59470 288696 59472
rect 286869 59467 286935 59470
rect 283925 59392 286764 59394
rect 283925 59336 283930 59392
rect 283986 59336 286764 59392
rect 283925 59334 286764 59336
rect 286869 59394 286935 59397
rect 289648 59394 289708 60044
rect 289813 59802 289879 59805
rect 290660 59802 290720 60044
rect 289813 59800 290720 59802
rect 289813 59744 289818 59800
rect 289874 59744 290720 59800
rect 289813 59742 290720 59744
rect 289813 59739 289879 59742
rect 291580 59666 291640 60044
rect 286869 59392 289708 59394
rect 286869 59336 286874 59392
rect 286930 59336 289708 59392
rect 286869 59334 289708 59336
rect 289862 59606 291640 59666
rect 283925 59331 283991 59334
rect 286869 59331 286935 59334
rect 279877 59256 280170 59258
rect 279877 59200 279882 59256
rect 279938 59200 280170 59256
rect 279877 59198 280170 59200
rect 289077 59258 289143 59261
rect 289862 59258 289922 59606
rect 290641 59530 290707 59533
rect 292592 59530 292652 60044
rect 292757 59802 292823 59805
rect 293512 59802 293572 60044
rect 292757 59800 293572 59802
rect 292757 59744 292762 59800
rect 292818 59744 293572 59800
rect 292757 59742 293572 59744
rect 292757 59739 292823 59742
rect 294524 59666 294584 60044
rect 290641 59528 292652 59530
rect 290641 59472 290646 59528
rect 290702 59472 292652 59528
rect 290641 59470 292652 59472
rect 292806 59606 294584 59666
rect 290641 59467 290707 59470
rect 291837 59394 291903 59397
rect 292806 59394 292866 59606
rect 293217 59530 293283 59533
rect 295444 59530 295504 60044
rect 293217 59528 295504 59530
rect 293217 59472 293222 59528
rect 293278 59472 295504 59528
rect 293217 59470 295504 59472
rect 293217 59467 293283 59470
rect 291837 59392 292866 59394
rect 291837 59336 291842 59392
rect 291898 59336 292866 59392
rect 291837 59334 292866 59336
rect 293401 59394 293467 59397
rect 296456 59394 296516 60044
rect 296621 59666 296687 59669
rect 297468 59666 297528 60044
rect 296621 59664 297528 59666
rect 296621 59608 296626 59664
rect 296682 59608 297528 59664
rect 296621 59606 297528 59608
rect 296621 59603 296687 59606
rect 296621 59530 296687 59533
rect 298388 59530 298448 60044
rect 296621 59528 298448 59530
rect 296621 59472 296626 59528
rect 296682 59472 298448 59528
rect 296621 59470 298448 59472
rect 296621 59467 296687 59470
rect 299400 59394 299460 60044
rect 300320 59530 300380 60044
rect 301332 59666 301392 60044
rect 302344 59802 302404 60044
rect 303264 59938 303324 60044
rect 303264 59878 304090 59938
rect 302344 59742 303906 59802
rect 303613 59666 303679 59669
rect 301332 59664 303679 59666
rect 301332 59608 303618 59664
rect 303674 59608 303679 59664
rect 301332 59606 303679 59608
rect 303613 59603 303679 59606
rect 302233 59530 302299 59533
rect 300320 59528 302299 59530
rect 300320 59472 302238 59528
rect 302294 59472 302299 59528
rect 300320 59470 302299 59472
rect 302233 59467 302299 59470
rect 293401 59392 296516 59394
rect 293401 59336 293406 59392
rect 293462 59336 296516 59392
rect 293401 59334 296516 59336
rect 296670 59334 299460 59394
rect 291837 59331 291903 59334
rect 293401 59331 293467 59334
rect 289077 59256 289922 59258
rect 289077 59200 289082 59256
rect 289138 59200 289922 59256
rect 289077 59198 289922 59200
rect 296161 59258 296227 59261
rect 296670 59258 296730 59334
rect 296161 59256 296730 59258
rect 296161 59200 296166 59256
rect 296222 59200 296730 59256
rect 296161 59198 296730 59200
rect 246849 59195 246915 59198
rect 270125 59195 270191 59198
rect 279877 59195 279943 59198
rect 289077 59195 289143 59198
rect 296161 59195 296227 59198
rect 237281 59120 239322 59122
rect 237281 59064 237286 59120
rect 237342 59064 239322 59120
rect 237281 59062 239322 59064
rect 303846 59122 303906 59742
rect 304030 59258 304090 59878
rect 304276 59394 304336 60044
rect 305196 59938 305256 60044
rect 305134 59878 305256 59938
rect 304993 59802 305059 59805
rect 305134 59802 305194 59878
rect 304993 59800 305194 59802
rect 304993 59744 304998 59800
rect 305054 59744 305194 59800
rect 304993 59742 305194 59744
rect 304993 59739 305059 59742
rect 306208 59530 306268 60044
rect 307128 59530 307188 60044
rect 308140 59666 308200 60044
rect 308949 59802 309015 59805
rect 309152 59802 309212 60044
rect 308949 59800 309212 59802
rect 308949 59744 308954 59800
rect 309010 59744 309212 59800
rect 308949 59742 309212 59744
rect 308949 59739 309015 59742
rect 308140 59606 309978 59666
rect 309133 59530 309199 59533
rect 306208 59470 307034 59530
rect 307128 59528 309199 59530
rect 307128 59472 309138 59528
rect 309194 59472 309199 59528
rect 307128 59470 309199 59472
rect 306373 59394 306439 59397
rect 304276 59392 306439 59394
rect 304276 59336 306378 59392
rect 306434 59336 306439 59392
rect 304276 59334 306439 59336
rect 306974 59394 307034 59470
rect 309133 59467 309199 59470
rect 307937 59394 308003 59397
rect 306974 59392 308003 59394
rect 306974 59336 307942 59392
rect 307998 59336 308003 59392
rect 306974 59334 308003 59336
rect 309918 59394 309978 59606
rect 310072 59530 310132 60044
rect 311084 59666 311144 60044
rect 312004 59805 312064 60044
rect 311985 59800 312064 59805
rect 311985 59744 311990 59800
rect 312046 59744 312064 59800
rect 311985 59742 312064 59744
rect 311985 59739 312051 59742
rect 311084 59606 312186 59666
rect 310072 59470 311910 59530
rect 311850 59397 311910 59470
rect 310513 59394 310579 59397
rect 309918 59392 310579 59394
rect 309918 59336 310518 59392
rect 310574 59336 310579 59392
rect 309918 59334 310579 59336
rect 311850 59392 311959 59397
rect 311850 59336 311898 59392
rect 311954 59336 311959 59392
rect 311850 59334 311959 59336
rect 312126 59394 312186 59606
rect 313016 59530 313076 60044
rect 313936 59666 313996 60044
rect 314948 59802 315008 60044
rect 315757 59802 315823 59805
rect 314948 59800 315823 59802
rect 314948 59744 315762 59800
rect 315818 59744 315823 59800
rect 314948 59742 315823 59744
rect 315757 59739 315823 59742
rect 313936 59606 315866 59666
rect 314837 59530 314903 59533
rect 313016 59528 314903 59530
rect 313016 59472 314842 59528
rect 314898 59472 314903 59528
rect 313016 59470 314903 59472
rect 314837 59467 314903 59470
rect 313273 59394 313339 59397
rect 312126 59392 313339 59394
rect 312126 59336 313278 59392
rect 313334 59336 313339 59392
rect 312126 59334 313339 59336
rect 315806 59394 315866 59606
rect 315960 59530 316020 60044
rect 316880 59666 316940 60044
rect 317892 59802 317952 60044
rect 318812 59938 318872 60044
rect 318812 59878 319546 59938
rect 319486 59802 319546 59878
rect 319621 59802 319687 59805
rect 317892 59742 319362 59802
rect 319486 59800 319687 59802
rect 319486 59744 319626 59800
rect 319682 59744 319687 59800
rect 319486 59742 319687 59744
rect 318793 59666 318859 59669
rect 316880 59664 318859 59666
rect 316880 59608 318798 59664
rect 318854 59608 318859 59664
rect 316880 59606 318859 59608
rect 318793 59603 318859 59606
rect 317413 59530 317479 59533
rect 315960 59528 317479 59530
rect 315960 59472 317418 59528
rect 317474 59472 317479 59528
rect 315960 59470 317479 59472
rect 319302 59530 319362 59742
rect 319621 59739 319687 59742
rect 319824 59666 319884 60044
rect 320449 59666 320515 59669
rect 319824 59664 320515 59666
rect 319824 59608 320454 59664
rect 320510 59608 320515 59664
rect 319824 59606 320515 59608
rect 320449 59603 320515 59606
rect 320265 59530 320331 59533
rect 319302 59528 320331 59530
rect 319302 59472 320270 59528
rect 320326 59472 320331 59528
rect 319302 59470 320331 59472
rect 317413 59467 317479 59470
rect 320265 59467 320331 59470
rect 316125 59394 316191 59397
rect 315806 59392 316191 59394
rect 315806 59336 316130 59392
rect 316186 59336 316191 59392
rect 315806 59334 316191 59336
rect 320836 59394 320896 60044
rect 321756 59938 321816 60044
rect 321756 59878 322490 59938
rect 322430 59802 322490 59878
rect 322565 59802 322631 59805
rect 322430 59800 322631 59802
rect 322430 59744 322570 59800
rect 322626 59744 322631 59800
rect 322430 59742 322631 59744
rect 322565 59739 322631 59742
rect 322768 59530 322828 60044
rect 323688 59666 323748 60044
rect 324497 59666 324563 59669
rect 323688 59664 324563 59666
rect 323688 59608 324502 59664
rect 324558 59608 324563 59664
rect 323688 59606 324563 59608
rect 324497 59603 324563 59606
rect 324497 59530 324563 59533
rect 322768 59528 324563 59530
rect 322768 59472 324502 59528
rect 324558 59472 324563 59528
rect 322768 59470 324563 59472
rect 324497 59467 324563 59470
rect 322933 59394 322999 59397
rect 320836 59392 322999 59394
rect 320836 59336 322938 59392
rect 322994 59336 322999 59392
rect 320836 59334 322999 59336
rect 324700 59394 324760 60044
rect 325620 59666 325680 60044
rect 326153 59802 326219 59805
rect 326632 59802 326692 60044
rect 326153 59800 326692 59802
rect 326153 59744 326158 59800
rect 326214 59744 326692 59800
rect 326153 59742 326692 59744
rect 326153 59739 326219 59742
rect 327257 59666 327323 59669
rect 325620 59664 327323 59666
rect 325620 59608 327262 59664
rect 327318 59608 327323 59664
rect 325620 59606 327323 59608
rect 327257 59603 327323 59606
rect 327073 59394 327139 59397
rect 324700 59392 327139 59394
rect 324700 59336 327078 59392
rect 327134 59336 327139 59392
rect 324700 59334 327139 59336
rect 327644 59394 327704 60044
rect 328564 59533 328624 60044
rect 328545 59528 328624 59533
rect 328545 59472 328550 59528
rect 328606 59472 328624 59528
rect 328545 59470 328624 59472
rect 329576 59530 329636 60044
rect 330496 59666 330556 60044
rect 331508 59802 331568 60044
rect 332520 59938 332580 60044
rect 332520 59878 333346 59938
rect 331508 59742 332978 59802
rect 330496 59606 332426 59666
rect 331397 59530 331463 59533
rect 329576 59528 331463 59530
rect 329576 59472 331402 59528
rect 331458 59472 331463 59528
rect 329576 59470 331463 59472
rect 328545 59467 328611 59470
rect 331397 59467 331463 59470
rect 329925 59394 329991 59397
rect 327644 59392 329991 59394
rect 327644 59336 329930 59392
rect 329986 59336 329991 59392
rect 327644 59334 329991 59336
rect 332366 59394 332426 59606
rect 332593 59394 332659 59397
rect 332366 59392 332659 59394
rect 332366 59336 332598 59392
rect 332654 59336 332659 59392
rect 332366 59334 332659 59336
rect 332918 59394 332978 59742
rect 333286 59666 333346 59878
rect 333440 59802 333500 60044
rect 334452 59938 334512 60044
rect 334452 59878 335002 59938
rect 334341 59802 334407 59805
rect 333440 59800 334407 59802
rect 333440 59744 334346 59800
rect 334402 59744 334407 59800
rect 333440 59742 334407 59744
rect 334341 59739 334407 59742
rect 334157 59666 334223 59669
rect 333286 59664 334223 59666
rect 333286 59608 334162 59664
rect 334218 59608 334223 59664
rect 333286 59606 334223 59608
rect 334157 59603 334223 59606
rect 334249 59394 334315 59397
rect 332918 59392 334315 59394
rect 332918 59336 334254 59392
rect 334310 59336 334315 59392
rect 332918 59334 334315 59336
rect 334942 59394 335002 59878
rect 335372 59530 335432 60044
rect 336384 59530 336444 60044
rect 337304 59666 337364 60044
rect 338316 59802 338376 60044
rect 339125 59802 339191 59805
rect 338316 59800 339191 59802
rect 338316 59744 339130 59800
rect 339186 59744 339191 59800
rect 338316 59742 339191 59744
rect 339125 59739 339191 59742
rect 337304 59606 339234 59666
rect 338297 59530 338363 59533
rect 335372 59470 336290 59530
rect 336384 59528 338363 59530
rect 336384 59472 338302 59528
rect 338358 59472 338363 59528
rect 336384 59470 338363 59472
rect 336230 59394 336290 59470
rect 338297 59467 338363 59470
rect 338481 59394 338547 59397
rect 334942 59334 336106 59394
rect 336230 59392 338547 59394
rect 336230 59336 338486 59392
rect 338542 59336 338547 59392
rect 336230 59334 338547 59336
rect 339174 59394 339234 59606
rect 339328 59530 339388 60044
rect 340248 59666 340308 60044
rect 340873 59802 340939 59805
rect 341260 59802 341320 60044
rect 340873 59800 341320 59802
rect 340873 59744 340878 59800
rect 340934 59744 341320 59800
rect 340873 59742 341320 59744
rect 340873 59739 340939 59742
rect 340248 59606 341994 59666
rect 341149 59530 341215 59533
rect 339328 59528 341215 59530
rect 339328 59472 341154 59528
rect 341210 59472 341215 59528
rect 339328 59470 341215 59472
rect 341149 59467 341215 59470
rect 339493 59394 339559 59397
rect 339174 59392 339559 59394
rect 339174 59336 339498 59392
rect 339554 59336 339559 59392
rect 339174 59334 339559 59336
rect 306373 59331 306439 59334
rect 307937 59331 308003 59334
rect 310513 59331 310579 59334
rect 311893 59331 311959 59334
rect 313273 59331 313339 59334
rect 316125 59331 316191 59334
rect 322933 59331 322999 59334
rect 327073 59331 327139 59334
rect 329925 59331 329991 59334
rect 332593 59331 332659 59334
rect 334249 59331 334315 59334
rect 305269 59258 305335 59261
rect 304030 59256 305335 59258
rect 304030 59200 305274 59256
rect 305330 59200 305335 59256
rect 304030 59198 305335 59200
rect 336046 59258 336106 59334
rect 338481 59331 338547 59334
rect 339493 59331 339559 59334
rect 336733 59258 336799 59261
rect 336046 59256 336799 59258
rect 336046 59200 336738 59256
rect 336794 59200 336799 59256
rect 336046 59198 336799 59200
rect 341934 59258 341994 59606
rect 342180 59394 342240 60044
rect 343192 59394 343252 60044
rect 344112 59802 344172 60044
rect 345124 59938 345184 60044
rect 345124 59878 345490 59938
rect 345430 59805 345490 59878
rect 344112 59742 345306 59802
rect 345246 59530 345306 59742
rect 345381 59800 345490 59805
rect 345381 59744 345386 59800
rect 345442 59744 345490 59800
rect 345381 59742 345490 59744
rect 345381 59739 345447 59742
rect 346136 59666 346196 60044
rect 347056 59802 347116 60044
rect 347681 59802 347747 59805
rect 347056 59800 347747 59802
rect 347056 59744 347686 59800
rect 347742 59744 347747 59800
rect 347056 59742 347747 59744
rect 347681 59739 347747 59742
rect 347865 59666 347931 59669
rect 346136 59664 347931 59666
rect 346136 59608 347870 59664
rect 347926 59608 347931 59664
rect 346136 59606 347931 59608
rect 347865 59603 347931 59606
rect 346485 59530 346551 59533
rect 345246 59528 346551 59530
rect 345246 59472 346490 59528
rect 346546 59472 346551 59528
rect 345246 59470 346551 59472
rect 346485 59467 346551 59470
rect 347773 59530 347839 59533
rect 348068 59530 348128 60044
rect 347773 59528 348128 59530
rect 347773 59472 347778 59528
rect 347834 59472 348128 59528
rect 347773 59470 348128 59472
rect 348988 59530 349048 60044
rect 349153 59530 349219 59533
rect 348988 59528 349219 59530
rect 348988 59472 349158 59528
rect 349214 59472 349219 59528
rect 348988 59470 349219 59472
rect 350000 59530 350060 60044
rect 350000 59470 350826 59530
rect 347773 59467 347839 59470
rect 349153 59467 349219 59470
rect 345013 59394 345079 59397
rect 342180 59334 343098 59394
rect 343192 59392 345079 59394
rect 343192 59336 345018 59392
rect 345074 59336 345079 59392
rect 343192 59334 345079 59336
rect 342253 59258 342319 59261
rect 341934 59256 342319 59258
rect 341934 59200 342258 59256
rect 342314 59200 342319 59256
rect 341934 59198 342319 59200
rect 343038 59258 343098 59334
rect 345013 59331 345079 59334
rect 347681 59394 347747 59397
rect 349337 59394 349403 59397
rect 347681 59392 349403 59394
rect 347681 59336 347686 59392
rect 347742 59336 349342 59392
rect 349398 59336 349403 59392
rect 347681 59334 349403 59336
rect 347681 59331 347747 59334
rect 349337 59331 349403 59334
rect 343817 59258 343883 59261
rect 343038 59256 343883 59258
rect 343038 59200 343822 59256
rect 343878 59200 343883 59256
rect 343038 59198 343883 59200
rect 350766 59258 350826 59470
rect 351012 59394 351072 60044
rect 351932 59530 351992 60044
rect 352741 59530 352807 59533
rect 351932 59528 352807 59530
rect 351932 59472 352746 59528
rect 352802 59472 352807 59528
rect 351932 59470 352807 59472
rect 352944 59530 353004 60044
rect 353864 59666 353924 60044
rect 354876 59802 354936 60044
rect 355593 59802 355659 59805
rect 354876 59800 355659 59802
rect 354876 59744 355598 59800
rect 355654 59744 355659 59800
rect 354876 59742 355659 59744
rect 355593 59739 355659 59742
rect 353864 59606 355610 59666
rect 355317 59530 355383 59533
rect 352944 59528 355383 59530
rect 352944 59472 355322 59528
rect 355378 59472 355383 59528
rect 352944 59470 355383 59472
rect 352741 59467 352807 59470
rect 355317 59467 355383 59470
rect 353937 59394 354003 59397
rect 351012 59392 354003 59394
rect 351012 59336 353942 59392
rect 353998 59336 354003 59392
rect 351012 59334 354003 59336
rect 355550 59394 355610 59606
rect 355796 59530 355856 60044
rect 356808 59666 356868 60044
rect 357617 59666 357683 59669
rect 356808 59664 357683 59666
rect 356808 59608 357622 59664
rect 357678 59608 357683 59664
rect 356808 59606 357683 59608
rect 357820 59666 357880 60044
rect 358740 59666 358800 60044
rect 359752 59938 359812 60044
rect 360672 59938 360732 60044
rect 359752 59878 360394 59938
rect 360672 59878 361498 59938
rect 360334 59805 360394 59878
rect 361438 59805 361498 59878
rect 360334 59800 360443 59805
rect 360334 59744 360382 59800
rect 360438 59744 360443 59800
rect 360334 59742 360443 59744
rect 361438 59800 361547 59805
rect 361438 59744 361486 59800
rect 361542 59744 361547 59800
rect 361438 59742 361547 59744
rect 361684 59802 361744 60044
rect 362696 59938 362756 60044
rect 362696 59878 363522 59938
rect 361684 59742 362602 59802
rect 360377 59739 360443 59742
rect 361481 59739 361547 59742
rect 362542 59666 362602 59742
rect 363321 59666 363387 59669
rect 357820 59606 358554 59666
rect 358740 59606 360732 59666
rect 362542 59664 363387 59666
rect 362542 59608 363326 59664
rect 363382 59608 363387 59664
rect 362542 59606 363387 59608
rect 357617 59603 357683 59606
rect 358077 59530 358143 59533
rect 355796 59528 358143 59530
rect 355796 59472 358082 59528
rect 358138 59472 358143 59528
rect 355796 59470 358143 59472
rect 358494 59530 358554 59606
rect 360469 59530 360535 59533
rect 358494 59528 360535 59530
rect 358494 59472 360474 59528
rect 360530 59472 360535 59528
rect 358494 59470 360535 59472
rect 360672 59530 360732 59606
rect 363321 59603 363387 59606
rect 361021 59530 361087 59533
rect 362217 59530 362283 59533
rect 360672 59528 361087 59530
rect 360672 59472 361026 59528
rect 361082 59472 361087 59528
rect 360672 59470 361087 59472
rect 358077 59467 358143 59470
rect 360469 59467 360535 59470
rect 361021 59467 361087 59470
rect 361254 59528 362283 59530
rect 361254 59472 362222 59528
rect 362278 59472 362283 59528
rect 361254 59470 362283 59472
rect 363462 59530 363522 59878
rect 363616 59666 363676 60044
rect 364628 59938 364688 60044
rect 364628 59878 365362 59938
rect 365302 59805 365362 59878
rect 365302 59800 365411 59805
rect 365302 59744 365350 59800
rect 365406 59744 365411 59800
rect 365302 59742 365411 59744
rect 365345 59739 365411 59742
rect 363616 59606 365362 59666
rect 365161 59530 365227 59533
rect 363462 59528 365227 59530
rect 363462 59472 365166 59528
rect 365222 59472 365227 59528
rect 363462 59470 365227 59472
rect 356697 59394 356763 59397
rect 355550 59392 356763 59394
rect 355550 59336 356702 59392
rect 356758 59336 356763 59392
rect 355550 59334 356763 59336
rect 353937 59331 354003 59334
rect 356697 59331 356763 59334
rect 357617 59394 357683 59397
rect 359457 59394 359523 59397
rect 357617 59392 359523 59394
rect 357617 59336 357622 59392
rect 357678 59336 359462 59392
rect 359518 59336 359523 59392
rect 357617 59334 359523 59336
rect 357617 59331 357683 59334
rect 359457 59331 359523 59334
rect 360377 59394 360443 59397
rect 361254 59394 361314 59470
rect 362217 59467 362283 59470
rect 365161 59467 365227 59470
rect 360377 59392 361314 59394
rect 360377 59336 360382 59392
rect 360438 59336 361314 59392
rect 360377 59334 361314 59336
rect 361481 59394 361547 59397
rect 363597 59394 363663 59397
rect 361481 59392 363663 59394
rect 361481 59336 361486 59392
rect 361542 59336 363602 59392
rect 363658 59336 363663 59392
rect 361481 59334 363663 59336
rect 360377 59331 360443 59334
rect 361481 59331 361547 59334
rect 363597 59331 363663 59334
rect 363781 59394 363847 59397
rect 364977 59394 365043 59397
rect 363781 59392 365043 59394
rect 363781 59336 363786 59392
rect 363842 59336 364982 59392
rect 365038 59336 365043 59392
rect 363781 59334 365043 59336
rect 363781 59331 363847 59334
rect 364977 59331 365043 59334
rect 352557 59258 352623 59261
rect 350766 59256 352623 59258
rect 350766 59200 352562 59256
rect 352618 59200 352623 59256
rect 350766 59198 352623 59200
rect 365302 59258 365362 59606
rect 365548 59394 365608 60044
rect 366560 59530 366620 60044
rect 367480 59666 367540 60044
rect 368492 59802 368552 60044
rect 369301 59802 369367 59805
rect 368492 59800 369367 59802
rect 368492 59744 369306 59800
rect 369362 59744 369367 59800
rect 368492 59742 369367 59744
rect 369301 59739 369367 59742
rect 367480 59606 369410 59666
rect 369117 59530 369183 59533
rect 366560 59528 369183 59530
rect 366560 59472 369122 59528
rect 369178 59472 369183 59528
rect 366560 59470 369183 59472
rect 369117 59467 369183 59470
rect 365548 59334 367386 59394
rect 366357 59258 366423 59261
rect 365302 59256 366423 59258
rect 365302 59200 366362 59256
rect 366418 59200 366423 59256
rect 365302 59198 366423 59200
rect 367326 59258 367386 59334
rect 367921 59258 367987 59261
rect 367326 59256 367987 59258
rect 367326 59200 367926 59256
rect 367982 59200 367987 59256
rect 367326 59198 367987 59200
rect 369350 59258 369410 59606
rect 369504 59394 369564 60044
rect 370424 59530 370484 60044
rect 371141 59530 371207 59533
rect 370424 59528 371207 59530
rect 370424 59472 371146 59528
rect 371202 59472 371207 59528
rect 370424 59470 371207 59472
rect 371141 59467 371207 59470
rect 371436 59394 371496 60044
rect 372356 59530 372416 60044
rect 373368 59666 373428 60044
rect 374085 59666 374151 59669
rect 373368 59664 374151 59666
rect 373368 59608 374090 59664
rect 374146 59608 374151 59664
rect 373368 59606 374151 59608
rect 374085 59603 374151 59606
rect 374085 59530 374151 59533
rect 372356 59528 374151 59530
rect 372356 59472 374090 59528
rect 374146 59472 374151 59528
rect 372356 59470 374151 59472
rect 374085 59467 374151 59470
rect 374085 59394 374151 59397
rect 369504 59334 371250 59394
rect 371436 59392 374151 59394
rect 371436 59336 374090 59392
rect 374146 59336 374151 59392
rect 371436 59334 374151 59336
rect 374288 59394 374348 60044
rect 375300 59530 375360 60044
rect 376312 59666 376372 60044
rect 377232 59802 377292 60044
rect 378041 59802 378107 59805
rect 377232 59800 378107 59802
rect 377232 59744 378046 59800
rect 378102 59744 378107 59800
rect 377232 59742 378107 59744
rect 378041 59739 378107 59742
rect 376312 59606 378058 59666
rect 377581 59530 377647 59533
rect 375300 59528 377647 59530
rect 375300 59472 377586 59528
rect 377642 59472 377647 59528
rect 375300 59470 377647 59472
rect 377581 59467 377647 59470
rect 377397 59394 377463 59397
rect 374288 59392 377463 59394
rect 374288 59336 377402 59392
rect 377458 59336 377463 59392
rect 374288 59334 377463 59336
rect 370497 59258 370563 59261
rect 369350 59256 370563 59258
rect 369350 59200 370502 59256
rect 370558 59200 370563 59256
rect 369350 59198 370563 59200
rect 371190 59258 371250 59334
rect 374085 59331 374151 59334
rect 377397 59331 377463 59334
rect 372153 59258 372219 59261
rect 371190 59256 372219 59258
rect 371190 59200 372158 59256
rect 372214 59200 372219 59256
rect 371190 59198 372219 59200
rect 377998 59258 378058 59606
rect 378244 59394 378304 60044
rect 378409 59530 378475 59533
rect 379164 59530 379224 60044
rect 380176 59666 380236 60044
rect 381188 59802 381248 60044
rect 381905 59802 381971 59805
rect 381188 59800 381971 59802
rect 381188 59744 381910 59800
rect 381966 59744 381971 59800
rect 381188 59742 381971 59744
rect 381905 59739 381971 59742
rect 380176 59606 381922 59666
rect 381537 59530 381603 59533
rect 378409 59528 378978 59530
rect 378409 59472 378414 59528
rect 378470 59472 378978 59528
rect 378409 59470 378978 59472
rect 379164 59528 381603 59530
rect 379164 59472 381542 59528
rect 381598 59472 381603 59528
rect 379164 59470 381603 59472
rect 378409 59467 378475 59470
rect 378918 59394 378978 59470
rect 381537 59467 381603 59470
rect 380157 59394 380223 59397
rect 381721 59394 381787 59397
rect 378244 59334 378794 59394
rect 378918 59392 380223 59394
rect 378918 59336 380162 59392
rect 380218 59336 380223 59392
rect 378918 59334 380223 59336
rect 378593 59258 378659 59261
rect 377998 59256 378659 59258
rect 377998 59200 378598 59256
rect 378654 59200 378659 59256
rect 377998 59198 378659 59200
rect 378734 59258 378794 59334
rect 380157 59331 380223 59334
rect 380390 59392 381787 59394
rect 380390 59336 381726 59392
rect 381782 59336 381787 59392
rect 380390 59334 381787 59336
rect 381862 59394 381922 59606
rect 382108 59530 382168 60044
rect 383120 59938 383180 60044
rect 383120 59878 383210 59938
rect 383150 59666 383210 59878
rect 383285 59802 383351 59805
rect 383837 59802 383903 59805
rect 383285 59800 383903 59802
rect 383285 59744 383290 59800
rect 383346 59744 383842 59800
rect 383898 59744 383903 59800
rect 383285 59742 383903 59744
rect 384040 59802 384100 60044
rect 384849 59802 384915 59805
rect 384040 59800 384915 59802
rect 384040 59744 384854 59800
rect 384910 59744 384915 59800
rect 384040 59742 384915 59744
rect 385052 59802 385112 60044
rect 385972 59938 386032 60044
rect 385972 59878 386890 59938
rect 385953 59802 386019 59805
rect 385052 59800 386019 59802
rect 385052 59744 385958 59800
rect 386014 59744 386019 59800
rect 385052 59742 386019 59744
rect 383285 59739 383351 59742
rect 383837 59739 383903 59742
rect 384849 59739 384915 59742
rect 385953 59739 386019 59742
rect 385677 59666 385743 59669
rect 383150 59664 385743 59666
rect 383150 59608 385682 59664
rect 385738 59608 385743 59664
rect 383150 59606 385743 59608
rect 385677 59603 385743 59606
rect 383837 59530 383903 59533
rect 382108 59528 383903 59530
rect 382108 59472 383842 59528
rect 383898 59472 383903 59528
rect 382108 59470 383903 59472
rect 386830 59530 386890 59878
rect 386984 59666 387044 60044
rect 387996 59802 388056 60044
rect 388713 59802 388779 59805
rect 387996 59800 388779 59802
rect 387996 59744 388718 59800
rect 388774 59744 388779 59800
rect 387996 59742 388779 59744
rect 388713 59739 388779 59742
rect 386984 59606 388730 59666
rect 388437 59530 388503 59533
rect 386830 59528 388503 59530
rect 386830 59472 388442 59528
rect 388498 59472 388503 59528
rect 386830 59470 388503 59472
rect 383837 59467 383903 59470
rect 388437 59467 388503 59470
rect 383009 59394 383075 59397
rect 381862 59392 383075 59394
rect 381862 59336 383014 59392
rect 383070 59336 383075 59392
rect 381862 59334 383075 59336
rect 380390 59258 380450 59334
rect 381721 59331 381787 59334
rect 383009 59331 383075 59334
rect 384849 59394 384915 59397
rect 387057 59394 387123 59397
rect 384849 59392 387123 59394
rect 384849 59336 384854 59392
rect 384910 59336 387062 59392
rect 387118 59336 387123 59392
rect 384849 59334 387123 59336
rect 388670 59394 388730 59606
rect 388916 59530 388976 60044
rect 389928 59666 389988 60044
rect 390848 59802 390908 60044
rect 391657 59802 391723 59805
rect 390848 59800 391723 59802
rect 390848 59744 391662 59800
rect 391718 59744 391723 59800
rect 390848 59742 391723 59744
rect 391657 59739 391723 59742
rect 389928 59606 391674 59666
rect 391197 59530 391263 59533
rect 388916 59528 391263 59530
rect 388916 59472 391202 59528
rect 391258 59472 391263 59528
rect 388916 59470 391263 59472
rect 391197 59467 391263 59470
rect 389817 59394 389883 59397
rect 388670 59392 389883 59394
rect 388670 59336 389822 59392
rect 389878 59336 389883 59392
rect 388670 59334 389883 59336
rect 391614 59394 391674 59606
rect 391860 59530 391920 60044
rect 392872 59666 392932 60044
rect 393792 59802 393852 60044
rect 394601 59802 394667 59805
rect 393792 59800 394667 59802
rect 393792 59744 394606 59800
rect 394662 59744 394667 59800
rect 393792 59742 394667 59744
rect 394804 59802 394864 60044
rect 395724 59938 395784 60044
rect 395724 59878 396642 59938
rect 395705 59802 395771 59805
rect 394804 59800 395771 59802
rect 394804 59744 395710 59800
rect 395766 59744 395771 59800
rect 394804 59742 395771 59744
rect 394601 59739 394667 59742
rect 395705 59739 395771 59742
rect 395337 59666 395403 59669
rect 392872 59664 395403 59666
rect 392872 59608 395342 59664
rect 395398 59608 395403 59664
rect 392872 59606 395403 59608
rect 395337 59603 395403 59606
rect 393589 59530 393655 59533
rect 391860 59528 393655 59530
rect 391860 59472 393594 59528
rect 393650 59472 393655 59528
rect 391860 59470 393655 59472
rect 396582 59530 396642 59878
rect 396736 59666 396796 60044
rect 397656 59938 397716 60044
rect 397656 59878 398482 59938
rect 398422 59805 398482 59878
rect 398422 59800 398531 59805
rect 398422 59744 398470 59800
rect 398526 59744 398531 59800
rect 398422 59742 398531 59744
rect 398465 59739 398531 59742
rect 396736 59606 398482 59666
rect 398281 59530 398347 59533
rect 396582 59528 398347 59530
rect 396582 59472 398286 59528
rect 398342 59472 398347 59528
rect 396582 59470 398347 59472
rect 393589 59467 393655 59470
rect 398281 59467 398347 59470
rect 392669 59394 392735 59397
rect 391614 59392 392735 59394
rect 391614 59336 392674 59392
rect 392730 59336 392735 59392
rect 391614 59334 392735 59336
rect 384849 59331 384915 59334
rect 387057 59331 387123 59334
rect 389817 59331 389883 59334
rect 392669 59331 392735 59334
rect 394601 59394 394667 59397
rect 396717 59394 396783 59397
rect 394601 59392 396783 59394
rect 394601 59336 394606 59392
rect 394662 59336 396722 59392
rect 396778 59336 396783 59392
rect 394601 59334 396783 59336
rect 398422 59394 398482 59606
rect 398668 59530 398728 60044
rect 399680 59530 399740 60044
rect 400600 59666 400660 60044
rect 401612 59802 401672 60044
rect 402532 59938 402592 60044
rect 403544 59938 403604 60044
rect 402532 59878 403450 59938
rect 403544 59878 404186 59938
rect 402421 59802 402487 59805
rect 401612 59800 402487 59802
rect 401612 59744 402426 59800
rect 402482 59744 402487 59800
rect 401612 59742 402487 59744
rect 402421 59739 402487 59742
rect 402329 59666 402395 59669
rect 400600 59664 402395 59666
rect 400600 59608 402334 59664
rect 402390 59608 402395 59664
rect 400600 59606 402395 59608
rect 402329 59603 402395 59606
rect 402237 59530 402303 59533
rect 398668 59470 399586 59530
rect 399680 59528 402303 59530
rect 399680 59472 402242 59528
rect 402298 59472 402303 59528
rect 399680 59470 402303 59472
rect 403390 59530 403450 59878
rect 404126 59666 404186 59878
rect 404464 59802 404524 60044
rect 405273 59802 405339 59805
rect 404464 59800 405339 59802
rect 404464 59744 405278 59800
rect 405334 59744 405339 59800
rect 404464 59742 405339 59744
rect 405273 59739 405339 59742
rect 404126 59606 405290 59666
rect 404997 59530 405063 59533
rect 403390 59528 405063 59530
rect 403390 59472 405002 59528
rect 405058 59472 405063 59528
rect 403390 59470 405063 59472
rect 399385 59394 399451 59397
rect 398422 59392 399451 59394
rect 398422 59336 399390 59392
rect 399446 59336 399451 59392
rect 398422 59334 399451 59336
rect 399526 59394 399586 59470
rect 402237 59467 402303 59470
rect 404997 59467 405063 59470
rect 400857 59394 400923 59397
rect 399526 59392 400923 59394
rect 399526 59336 400862 59392
rect 400918 59336 400923 59392
rect 399526 59334 400923 59336
rect 394601 59331 394667 59334
rect 396717 59331 396783 59334
rect 399385 59331 399451 59334
rect 400857 59331 400923 59334
rect 402329 59394 402395 59397
rect 403617 59394 403683 59397
rect 402329 59392 403683 59394
rect 402329 59336 402334 59392
rect 402390 59336 403622 59392
rect 403678 59336 403683 59392
rect 402329 59334 403683 59336
rect 405230 59394 405290 59606
rect 405476 59530 405536 60044
rect 406488 59666 406548 60044
rect 407408 59802 407468 60044
rect 408420 59938 408480 60044
rect 408420 59878 408602 59938
rect 408401 59802 408467 59805
rect 407408 59800 408467 59802
rect 407408 59744 408406 59800
rect 408462 59744 408467 59800
rect 407408 59742 408467 59744
rect 408401 59739 408467 59742
rect 408542 59666 408602 59878
rect 409340 59802 409400 60044
rect 410149 59802 410215 59805
rect 409340 59800 410215 59802
rect 409340 59744 410154 59800
rect 410210 59744 410215 59800
rect 409340 59742 410215 59744
rect 410149 59739 410215 59742
rect 406488 59606 408050 59666
rect 407757 59530 407823 59533
rect 405476 59528 407823 59530
rect 405476 59472 407762 59528
rect 407818 59472 407823 59528
rect 405476 59470 407823 59472
rect 407757 59467 407823 59470
rect 406377 59394 406443 59397
rect 405230 59392 406443 59394
rect 405230 59336 406382 59392
rect 406438 59336 406443 59392
rect 405230 59334 406443 59336
rect 407990 59394 408050 59606
rect 408420 59606 408602 59666
rect 408677 59666 408743 59669
rect 410149 59666 410215 59669
rect 408677 59664 410215 59666
rect 408677 59608 408682 59664
rect 408738 59608 410154 59664
rect 410210 59608 410215 59664
rect 408677 59606 410215 59608
rect 410352 59666 410412 60044
rect 411364 59802 411424 60044
rect 412081 59802 412147 59805
rect 411364 59800 412147 59802
rect 411364 59744 412086 59800
rect 412142 59744 412147 59800
rect 411364 59742 412147 59744
rect 412081 59739 412147 59742
rect 410352 59606 410810 59666
rect 408420 59530 408480 59606
rect 408677 59603 408743 59606
rect 410149 59603 410215 59606
rect 410517 59530 410583 59533
rect 408420 59528 410583 59530
rect 408420 59472 410522 59528
rect 410578 59472 410583 59528
rect 408420 59470 410583 59472
rect 410750 59530 410810 59606
rect 412284 59530 412344 60044
rect 412449 59802 412515 59805
rect 413093 59802 413159 59805
rect 412449 59800 413159 59802
rect 412449 59744 412454 59800
rect 412510 59744 413098 59800
rect 413154 59744 413159 59800
rect 412449 59742 413159 59744
rect 412449 59739 412515 59742
rect 413093 59739 413159 59742
rect 413296 59666 413356 60044
rect 413921 59666 413987 59669
rect 413296 59664 413987 59666
rect 413296 59608 413926 59664
rect 413982 59608 413987 59664
rect 413296 59606 413987 59608
rect 413921 59603 413987 59606
rect 414013 59530 414079 59533
rect 410750 59470 411546 59530
rect 412284 59528 414079 59530
rect 412284 59472 414018 59528
rect 414074 59472 414079 59528
rect 412284 59470 414079 59472
rect 414216 59530 414276 60044
rect 415025 59530 415091 59533
rect 414216 59528 415091 59530
rect 414216 59472 415030 59528
rect 415086 59472 415091 59528
rect 414216 59470 415091 59472
rect 415228 59530 415288 60044
rect 416148 59666 416208 60044
rect 417160 59802 417220 60044
rect 418172 59938 418232 60044
rect 419092 59938 419152 60044
rect 418172 59878 418906 59938
rect 419092 59878 420010 59938
rect 417160 59742 418722 59802
rect 418153 59666 418219 59669
rect 416148 59664 418219 59666
rect 416148 59608 418158 59664
rect 418214 59608 418219 59664
rect 416148 59606 418219 59608
rect 418153 59603 418219 59606
rect 417049 59530 417115 59533
rect 415228 59528 417115 59530
rect 415228 59472 417054 59528
rect 417110 59472 417115 59528
rect 415228 59470 417115 59472
rect 418662 59530 418722 59742
rect 418846 59666 418906 59878
rect 419809 59666 419875 59669
rect 418846 59664 419875 59666
rect 418846 59608 419814 59664
rect 419870 59608 419875 59664
rect 418846 59606 419875 59608
rect 419809 59603 419875 59606
rect 419533 59530 419599 59533
rect 418662 59528 419599 59530
rect 418662 59472 419538 59528
rect 419594 59472 419599 59528
rect 418662 59470 419599 59472
rect 410517 59467 410583 59470
rect 409137 59394 409203 59397
rect 407990 59392 409203 59394
rect 407990 59336 409142 59392
rect 409198 59336 409203 59392
rect 407990 59334 409203 59336
rect 402329 59331 402395 59334
rect 403617 59331 403683 59334
rect 406377 59331 406443 59334
rect 409137 59331 409203 59334
rect 410149 59394 410215 59397
rect 410701 59394 410767 59397
rect 410149 59392 410767 59394
rect 410149 59336 410154 59392
rect 410210 59336 410706 59392
rect 410762 59336 410767 59392
rect 410149 59334 410767 59336
rect 411486 59394 411546 59470
rect 414013 59467 414079 59470
rect 415025 59467 415091 59470
rect 417049 59467 417115 59470
rect 419533 59467 419599 59470
rect 413093 59394 413159 59397
rect 411486 59392 413159 59394
rect 411486 59336 413098 59392
rect 413154 59336 413159 59392
rect 411486 59334 413159 59336
rect 410149 59331 410215 59334
rect 410701 59331 410767 59334
rect 413093 59331 413159 59334
rect 413921 59394 413987 59397
rect 415393 59394 415459 59397
rect 413921 59392 415459 59394
rect 413921 59336 413926 59392
rect 413982 59336 415398 59392
rect 415454 59336 415459 59392
rect 413921 59334 415459 59336
rect 413921 59331 413987 59334
rect 415393 59331 415459 59334
rect 415577 59394 415643 59397
rect 416865 59394 416931 59397
rect 415577 59392 416931 59394
rect 415577 59336 415582 59392
rect 415638 59336 416870 59392
rect 416926 59336 416931 59392
rect 415577 59334 416931 59336
rect 415577 59331 415643 59334
rect 416865 59331 416931 59334
rect 378734 59198 380450 59258
rect 305269 59195 305335 59198
rect 336733 59195 336799 59198
rect 342253 59195 342319 59198
rect 343817 59195 343883 59198
rect 352557 59195 352623 59198
rect 366357 59195 366423 59198
rect 367921 59195 367987 59198
rect 370497 59195 370563 59198
rect 372153 59195 372219 59198
rect 378593 59195 378659 59198
rect 305085 59122 305151 59125
rect 303846 59120 305151 59122
rect 303846 59064 305090 59120
rect 305146 59064 305151 59120
rect 303846 59062 305151 59064
rect 419950 59122 420010 59878
rect 420104 59394 420164 60044
rect 421024 59530 421084 60044
rect 421833 59530 421899 59533
rect 421024 59528 421899 59530
rect 421024 59472 421838 59528
rect 421894 59472 421899 59528
rect 421024 59470 421899 59472
rect 421833 59467 421899 59470
rect 422036 59394 422096 60044
rect 423048 59394 423108 60044
rect 423968 59530 424028 60044
rect 424777 59530 424843 59533
rect 423968 59528 424843 59530
rect 423968 59472 424782 59528
rect 424838 59472 424843 59528
rect 423968 59470 424843 59472
rect 424980 59530 425040 60044
rect 425900 59666 425960 60044
rect 426912 59802 426972 60044
rect 427445 59802 427511 59805
rect 426912 59800 427511 59802
rect 426912 59744 427450 59800
rect 427506 59744 427511 59800
rect 426912 59742 427511 59744
rect 427445 59739 427511 59742
rect 427629 59802 427695 59805
rect 427832 59802 427892 60044
rect 427629 59800 427892 59802
rect 427629 59744 427634 59800
rect 427690 59744 427892 59800
rect 427629 59742 427892 59744
rect 427629 59739 427695 59742
rect 427905 59666 427971 59669
rect 425900 59664 427971 59666
rect 425900 59608 427910 59664
rect 427966 59608 427971 59664
rect 425900 59606 427971 59608
rect 427905 59603 427971 59606
rect 426525 59530 426591 59533
rect 424980 59528 426591 59530
rect 424980 59472 426530 59528
rect 426586 59472 426591 59528
rect 424980 59470 426591 59472
rect 424777 59467 424843 59470
rect 426525 59467 426591 59470
rect 425053 59394 425119 59397
rect 420104 59334 420930 59394
rect 422036 59334 422954 59394
rect 423048 59392 425119 59394
rect 423048 59336 425058 59392
rect 425114 59336 425119 59392
rect 423048 59334 425119 59336
rect 420870 59258 420930 59334
rect 422385 59258 422451 59261
rect 420870 59256 422451 59258
rect 420870 59200 422390 59256
rect 422446 59200 422451 59256
rect 420870 59198 422451 59200
rect 422894 59258 422954 59334
rect 425053 59331 425119 59334
rect 425237 59394 425303 59397
rect 426709 59394 426775 59397
rect 425237 59392 426775 59394
rect 425237 59336 425242 59392
rect 425298 59336 426714 59392
rect 426770 59336 426775 59392
rect 425237 59334 426775 59336
rect 425237 59331 425303 59334
rect 426709 59331 426775 59334
rect 427445 59394 427511 59397
rect 428844 59394 428904 60044
rect 429856 59394 429916 60044
rect 430573 59530 430639 59533
rect 430776 59530 430836 60044
rect 430573 59528 430836 59530
rect 430573 59472 430578 59528
rect 430634 59472 430836 59528
rect 430573 59470 430836 59472
rect 431788 59530 431848 60044
rect 432708 59666 432768 60044
rect 433720 59802 433780 60044
rect 434437 59802 434503 59805
rect 433720 59800 434503 59802
rect 433720 59744 434442 59800
rect 434498 59744 434503 59800
rect 433720 59742 434503 59744
rect 434437 59739 434503 59742
rect 432708 59606 434546 59666
rect 433517 59530 433583 59533
rect 431788 59528 433583 59530
rect 431788 59472 433522 59528
rect 433578 59472 433583 59528
rect 431788 59470 433583 59472
rect 430573 59467 430639 59470
rect 433517 59467 433583 59470
rect 432045 59394 432111 59397
rect 427445 59392 428658 59394
rect 427445 59336 427450 59392
rect 427506 59336 428658 59392
rect 427445 59334 428658 59336
rect 428844 59334 429762 59394
rect 429856 59392 432111 59394
rect 429856 59336 432050 59392
rect 432106 59336 432111 59392
rect 429856 59334 432111 59336
rect 434486 59394 434546 59606
rect 434640 59530 434700 60044
rect 435652 59666 435712 60044
rect 436664 59802 436724 60044
rect 437584 59938 437644 60044
rect 437584 59878 438226 59938
rect 438025 59802 438091 59805
rect 436664 59800 438091 59802
rect 436664 59744 438030 59800
rect 438086 59744 438091 59800
rect 436664 59742 438091 59744
rect 438025 59739 438091 59742
rect 437565 59666 437631 59669
rect 435652 59664 437631 59666
rect 435652 59608 437570 59664
rect 437626 59608 437631 59664
rect 435652 59606 437631 59608
rect 437565 59603 437631 59606
rect 436185 59530 436251 59533
rect 434640 59528 436251 59530
rect 434640 59472 436190 59528
rect 436246 59472 436251 59528
rect 434640 59470 436251 59472
rect 436185 59467 436251 59470
rect 434713 59394 434779 59397
rect 434486 59392 434779 59394
rect 434486 59336 434718 59392
rect 434774 59336 434779 59392
rect 434486 59334 434779 59336
rect 427445 59331 427511 59334
rect 423949 59258 424015 59261
rect 422894 59256 424015 59258
rect 422894 59200 423954 59256
rect 424010 59200 424015 59256
rect 422894 59198 424015 59200
rect 428598 59258 428658 59334
rect 429193 59258 429259 59261
rect 428598 59256 429259 59258
rect 428598 59200 429198 59256
rect 429254 59200 429259 59256
rect 428598 59198 429259 59200
rect 429702 59258 429762 59334
rect 432045 59331 432111 59334
rect 434713 59331 434779 59334
rect 434897 59394 434963 59397
rect 436369 59394 436435 59397
rect 434897 59392 436435 59394
rect 434897 59336 434902 59392
rect 434958 59336 436374 59392
rect 436430 59336 436435 59392
rect 434897 59334 436435 59336
rect 434897 59331 434963 59334
rect 436369 59331 436435 59334
rect 430665 59258 430731 59261
rect 429702 59256 430731 59258
rect 429702 59200 430670 59256
rect 430726 59200 430731 59256
rect 429702 59198 430731 59200
rect 422385 59195 422451 59198
rect 423949 59195 424015 59198
rect 429193 59195 429259 59198
rect 430665 59195 430731 59198
rect 421281 59122 421347 59125
rect 419950 59120 421347 59122
rect 419950 59064 421286 59120
rect 421342 59064 421347 59120
rect 419950 59062 421347 59064
rect 104157 59059 104223 59062
rect 154021 59059 154087 59062
rect 184565 59059 184631 59062
rect 237281 59059 237347 59062
rect 305085 59059 305151 59062
rect 421281 59059 421347 59062
rect 421833 59122 421899 59125
rect 424133 59122 424199 59125
rect 421833 59120 424199 59122
rect 421833 59064 421838 59120
rect 421894 59064 424138 59120
rect 424194 59064 424199 59120
rect 421833 59062 424199 59064
rect 438166 59122 438226 59878
rect 438596 59394 438656 60044
rect 439516 59530 439576 60044
rect 440528 59666 440588 60044
rect 441061 59666 441127 59669
rect 440528 59664 441127 59666
rect 440528 59608 441066 59664
rect 441122 59608 441127 59664
rect 440528 59606 441127 59608
rect 441540 59666 441600 60044
rect 441981 59802 442047 59805
rect 442460 59802 442520 60044
rect 441981 59800 442520 59802
rect 441981 59744 441986 59800
rect 442042 59744 442520 59800
rect 441981 59742 442520 59744
rect 441981 59739 442047 59742
rect 443085 59666 443151 59669
rect 441540 59664 443151 59666
rect 441540 59608 443090 59664
rect 443146 59608 443151 59664
rect 441540 59606 443151 59608
rect 441061 59603 441127 59606
rect 443085 59603 443151 59606
rect 443472 59530 443532 60044
rect 444392 59666 444452 60044
rect 445404 59802 445464 60044
rect 446324 59938 446384 60044
rect 446324 59878 447196 59938
rect 446397 59802 446463 59805
rect 445404 59800 446463 59802
rect 445404 59744 446402 59800
rect 446458 59744 446463 59800
rect 445404 59742 446463 59744
rect 446397 59739 446463 59742
rect 447136 59669 447196 59878
rect 447336 59802 447396 60044
rect 448145 59802 448211 59805
rect 447336 59800 448211 59802
rect 447336 59744 448150 59800
rect 448206 59744 448211 59800
rect 447336 59742 448211 59744
rect 448145 59739 448211 59742
rect 446949 59666 447015 59669
rect 444392 59664 447015 59666
rect 444392 59608 446954 59664
rect 447010 59608 447015 59664
rect 444392 59606 447015 59608
rect 446949 59603 447015 59606
rect 447133 59664 447199 59669
rect 447133 59608 447138 59664
rect 447194 59608 447199 59664
rect 447133 59603 447199 59608
rect 445753 59530 445819 59533
rect 439516 59470 441630 59530
rect 443472 59528 445819 59530
rect 443472 59472 445758 59528
rect 445814 59472 445819 59528
rect 443472 59470 445819 59472
rect 448348 59530 448408 60044
rect 449268 59666 449328 60044
rect 449268 59606 450186 59666
rect 449985 59530 450051 59533
rect 448348 59528 450051 59530
rect 448348 59472 449990 59528
rect 450046 59472 450051 59528
rect 448348 59470 450051 59472
rect 441570 59397 441630 59470
rect 445753 59467 445819 59470
rect 449985 59467 450051 59470
rect 440509 59394 440575 59397
rect 438596 59392 440575 59394
rect 438596 59336 440514 59392
rect 440570 59336 440575 59392
rect 438596 59334 440575 59336
rect 440509 59331 440575 59334
rect 441061 59394 441127 59397
rect 441061 59392 441354 59394
rect 441061 59336 441066 59392
rect 441122 59336 441354 59392
rect 441061 59334 441354 59336
rect 441570 59392 441679 59397
rect 443269 59394 443335 59397
rect 441570 59336 441618 59392
rect 441674 59336 441679 59392
rect 441570 59334 441679 59336
rect 441061 59331 441127 59334
rect 441294 59258 441354 59334
rect 441613 59331 441679 59334
rect 441846 59392 443335 59394
rect 441846 59336 443274 59392
rect 443330 59336 443335 59392
rect 441846 59334 443335 59336
rect 441846 59258 441906 59334
rect 443269 59331 443335 59334
rect 441294 59198 441906 59258
rect 450126 59258 450186 59606
rect 450280 59394 450340 60044
rect 451200 59530 451260 60044
rect 452212 59666 452272 60044
rect 453224 59802 453284 60044
rect 453941 59802 454007 59805
rect 453224 59800 454007 59802
rect 453224 59744 453946 59800
rect 454002 59744 454007 59800
rect 453224 59742 454007 59744
rect 453941 59739 454007 59742
rect 452212 59606 454050 59666
rect 453021 59530 453087 59533
rect 451200 59528 453087 59530
rect 451200 59472 453026 59528
rect 453082 59472 453087 59528
rect 451200 59470 453087 59472
rect 453021 59467 453087 59470
rect 453990 59397 454050 59606
rect 454144 59530 454204 60044
rect 455156 59666 455216 60044
rect 455873 59666 455939 59669
rect 455156 59664 455939 59666
rect 455156 59608 455878 59664
rect 455934 59608 455939 59664
rect 455156 59606 455939 59608
rect 456076 59666 456136 60044
rect 456885 59666 456951 59669
rect 456076 59664 456951 59666
rect 456076 59608 456890 59664
rect 456946 59608 456951 59664
rect 456076 59606 456951 59608
rect 455873 59603 455939 59606
rect 456885 59603 456951 59606
rect 456609 59530 456675 59533
rect 456885 59530 456951 59533
rect 454144 59528 456675 59530
rect 454144 59472 456614 59528
rect 456670 59472 456675 59528
rect 454144 59470 456675 59472
rect 456609 59467 456675 59470
rect 456750 59528 456951 59530
rect 456750 59472 456890 59528
rect 456946 59472 456951 59528
rect 456750 59470 456951 59472
rect 452837 59394 452903 59397
rect 450280 59392 452903 59394
rect 450280 59336 452842 59392
rect 452898 59336 452903 59392
rect 450280 59334 452903 59336
rect 453990 59392 454099 59397
rect 453990 59336 454038 59392
rect 454094 59336 454099 59392
rect 453990 59334 454099 59336
rect 452837 59331 452903 59334
rect 454033 59331 454099 59334
rect 454217 59394 454283 59397
rect 455505 59394 455571 59397
rect 454217 59392 455571 59394
rect 454217 59336 454222 59392
rect 454278 59336 455510 59392
rect 455566 59336 455571 59392
rect 454217 59334 455571 59336
rect 454217 59331 454283 59334
rect 455505 59331 455571 59334
rect 455873 59394 455939 59397
rect 456750 59394 456810 59470
rect 456885 59467 456951 59470
rect 455873 59392 456810 59394
rect 455873 59336 455878 59392
rect 455934 59336 456810 59392
rect 455873 59334 456810 59336
rect 457088 59394 457148 60044
rect 458008 59530 458068 60044
rect 459020 59666 459080 60044
rect 460032 59802 460092 60044
rect 460952 59938 461012 60044
rect 460952 59878 461778 59938
rect 461577 59802 461643 59805
rect 460032 59800 461643 59802
rect 460032 59744 461582 59800
rect 461638 59744 461643 59800
rect 460032 59742 461643 59744
rect 461577 59739 461643 59742
rect 460933 59666 460999 59669
rect 459020 59664 460999 59666
rect 459020 59608 460938 59664
rect 460994 59608 460999 59664
rect 459020 59606 460999 59608
rect 460933 59603 460999 59606
rect 459829 59530 459895 59533
rect 458008 59528 459895 59530
rect 458008 59472 459834 59528
rect 459890 59472 459895 59528
rect 458008 59470 459895 59472
rect 459829 59467 459895 59470
rect 459645 59394 459711 59397
rect 457088 59392 459711 59394
rect 457088 59336 459650 59392
rect 459706 59336 459711 59392
rect 457088 59334 459711 59336
rect 461718 59394 461778 59878
rect 461964 59530 462024 60044
rect 462884 59666 462944 60044
rect 463601 59802 463667 59805
rect 463896 59802 463956 60044
rect 463601 59800 463956 59802
rect 463601 59744 463606 59800
rect 463662 59744 463956 59800
rect 463601 59742 463956 59744
rect 463601 59739 463667 59742
rect 462884 59606 464722 59666
rect 463693 59530 463759 59533
rect 461964 59528 463759 59530
rect 461964 59472 463698 59528
rect 463754 59472 463759 59528
rect 461964 59470 463759 59472
rect 463693 59467 463759 59470
rect 463877 59394 463943 59397
rect 461718 59392 463943 59394
rect 461718 59336 463882 59392
rect 463938 59336 463943 59392
rect 461718 59334 463943 59336
rect 464662 59394 464722 59606
rect 464816 59530 464876 60044
rect 465828 59666 465888 60044
rect 466840 59802 466900 60044
rect 467557 59802 467623 59805
rect 466840 59800 467623 59802
rect 466840 59744 467562 59800
rect 467618 59744 467623 59800
rect 466840 59742 467623 59744
rect 467557 59739 467623 59742
rect 465828 59606 467666 59666
rect 466637 59530 466703 59533
rect 464816 59528 466703 59530
rect 464816 59472 466642 59528
rect 466698 59472 466703 59528
rect 464816 59470 466703 59472
rect 466637 59467 466703 59470
rect 465073 59394 465139 59397
rect 464662 59392 465139 59394
rect 464662 59336 465078 59392
rect 465134 59336 465139 59392
rect 464662 59334 465139 59336
rect 467606 59394 467666 59606
rect 467760 59530 467820 60044
rect 468772 59666 468832 60044
rect 469692 59802 469752 60044
rect 470704 59938 470764 60044
rect 470704 59878 471530 59938
rect 470593 59802 470659 59805
rect 469692 59800 470659 59802
rect 469692 59744 470598 59800
rect 470654 59744 470659 59800
rect 469692 59742 470659 59744
rect 470593 59739 470659 59742
rect 470547 59666 470613 59669
rect 468772 59664 470613 59666
rect 468772 59608 470552 59664
rect 470608 59608 470613 59664
rect 468772 59606 470613 59608
rect 470547 59603 470613 59606
rect 469305 59530 469371 59533
rect 467760 59528 469371 59530
rect 467760 59472 469310 59528
rect 469366 59472 469371 59528
rect 467760 59470 469371 59472
rect 469305 59467 469371 59470
rect 467833 59394 467899 59397
rect 467606 59392 467899 59394
rect 467606 59336 467838 59392
rect 467894 59336 467899 59392
rect 467606 59334 467899 59336
rect 455873 59331 455939 59334
rect 459645 59331 459711 59334
rect 463877 59331 463943 59334
rect 465073 59331 465139 59334
rect 467833 59331 467899 59334
rect 468017 59394 468083 59397
rect 469489 59394 469555 59397
rect 468017 59392 469555 59394
rect 468017 59336 468022 59392
rect 468078 59336 469494 59392
rect 469550 59336 469555 59392
rect 468017 59334 469555 59336
rect 471470 59394 471530 59878
rect 471716 59530 471776 60044
rect 472636 59666 472696 60044
rect 473648 59802 473708 60044
rect 474365 59802 474431 59805
rect 473648 59800 474431 59802
rect 473648 59744 474370 59800
rect 474426 59744 474431 59800
rect 473648 59742 474431 59744
rect 474365 59739 474431 59742
rect 472636 59606 474474 59666
rect 473629 59530 473695 59533
rect 471716 59528 473695 59530
rect 471716 59472 473634 59528
rect 473690 59472 473695 59528
rect 471716 59470 473695 59472
rect 473629 59467 473695 59470
rect 473445 59394 473511 59397
rect 471470 59392 473511 59394
rect 471470 59336 473450 59392
rect 473506 59336 473511 59392
rect 471470 59334 473511 59336
rect 474414 59394 474474 59606
rect 474568 59530 474628 60044
rect 475580 59666 475640 60044
rect 476297 59666 476363 59669
rect 475580 59664 476363 59666
rect 475580 59608 476302 59664
rect 476358 59608 476363 59664
rect 475580 59606 476363 59608
rect 476297 59603 476363 59606
rect 476205 59530 476271 59533
rect 474568 59528 476271 59530
rect 474568 59472 476210 59528
rect 476266 59472 476271 59528
rect 474568 59470 476271 59472
rect 476500 59530 476560 60044
rect 477512 59666 477572 60044
rect 478321 59666 478387 59669
rect 477512 59664 478387 59666
rect 477512 59608 478326 59664
rect 478382 59608 478387 59664
rect 477512 59606 478387 59608
rect 478524 59666 478584 60044
rect 479444 59802 479504 60044
rect 480253 59802 480319 59805
rect 479444 59800 480319 59802
rect 479444 59744 480258 59800
rect 480314 59744 480319 59800
rect 479444 59742 480319 59744
rect 480253 59739 480319 59742
rect 480253 59666 480319 59669
rect 478524 59664 480319 59666
rect 478524 59608 480258 59664
rect 480314 59608 480319 59664
rect 478524 59606 480319 59608
rect 478321 59603 478387 59606
rect 480253 59603 480319 59606
rect 478873 59530 478939 59533
rect 476500 59528 478939 59530
rect 476500 59472 478878 59528
rect 478934 59472 478939 59528
rect 476500 59470 478939 59472
rect 480456 59530 480516 60044
rect 481376 59530 481436 60044
rect 482388 59666 482448 60044
rect 483308 59805 483368 60044
rect 483289 59800 483368 59805
rect 483289 59744 483294 59800
rect 483350 59744 483368 59800
rect 483289 59742 483368 59744
rect 483473 59802 483539 59805
rect 484320 59802 484380 60044
rect 483473 59800 484380 59802
rect 483473 59744 483478 59800
rect 483534 59744 484380 59800
rect 483473 59742 484380 59744
rect 483289 59739 483355 59742
rect 483473 59739 483539 59742
rect 484393 59666 484459 59669
rect 482388 59664 484459 59666
rect 482388 59608 484398 59664
rect 484454 59608 484459 59664
rect 482388 59606 484459 59608
rect 484393 59603 484459 59606
rect 483105 59530 483171 59533
rect 480456 59470 481282 59530
rect 481376 59528 483171 59530
rect 481376 59472 483110 59528
rect 483166 59472 483171 59528
rect 481376 59470 483171 59472
rect 485332 59530 485392 60044
rect 486252 59666 486312 60044
rect 487061 59666 487127 59669
rect 486252 59664 487127 59666
rect 486252 59608 487066 59664
rect 487122 59608 487127 59664
rect 486252 59606 487127 59608
rect 487264 59666 487324 60044
rect 488184 59802 488244 60044
rect 488441 59802 488507 59805
rect 488184 59800 488507 59802
rect 488184 59744 488446 59800
rect 488502 59744 488507 59800
rect 488184 59742 488507 59744
rect 488441 59739 488507 59742
rect 488625 59802 488691 59805
rect 489196 59802 489256 60044
rect 488625 59800 489256 59802
rect 488625 59744 488630 59800
rect 488686 59744 489256 59800
rect 488625 59742 489256 59744
rect 488625 59739 488691 59742
rect 489913 59666 489979 59669
rect 487264 59664 489979 59666
rect 487264 59608 489918 59664
rect 489974 59608 489979 59664
rect 487264 59606 489979 59608
rect 487061 59603 487127 59606
rect 489913 59603 489979 59606
rect 487245 59530 487311 59533
rect 485332 59528 487311 59530
rect 485332 59472 487250 59528
rect 487306 59472 487311 59528
rect 485332 59470 487311 59472
rect 476205 59467 476271 59470
rect 478873 59467 478939 59470
rect 474733 59394 474799 59397
rect 474414 59392 474799 59394
rect 474414 59336 474738 59392
rect 474794 59336 474799 59392
rect 474414 59334 474799 59336
rect 468017 59331 468083 59334
rect 469489 59331 469555 59334
rect 473445 59331 473511 59334
rect 474733 59331 474799 59334
rect 476297 59394 476363 59397
rect 477585 59394 477651 59397
rect 476297 59392 477651 59394
rect 476297 59336 476302 59392
rect 476358 59336 477590 59392
rect 477646 59336 477651 59392
rect 476297 59334 477651 59336
rect 476297 59331 476363 59334
rect 477585 59331 477651 59334
rect 478321 59394 478387 59397
rect 481222 59394 481282 59470
rect 483105 59467 483171 59470
rect 487245 59467 487311 59470
rect 488441 59530 488507 59533
rect 490005 59530 490071 59533
rect 488441 59528 490071 59530
rect 488441 59472 488446 59528
rect 488502 59472 490010 59528
rect 490066 59472 490071 59528
rect 488441 59470 490071 59472
rect 488441 59467 488507 59470
rect 490005 59467 490071 59470
rect 483289 59394 483355 59397
rect 485957 59394 486023 59397
rect 478321 59392 480270 59394
rect 478321 59336 478326 59392
rect 478382 59336 480270 59392
rect 478321 59334 480270 59336
rect 481222 59334 483122 59394
rect 478321 59331 478387 59334
rect 451273 59258 451339 59261
rect 450126 59256 451339 59258
rect 450126 59200 451278 59256
rect 451334 59200 451339 59256
rect 450126 59198 451339 59200
rect 480210 59258 480270 59334
rect 480345 59258 480411 59261
rect 480210 59256 480411 59258
rect 480210 59200 480350 59256
rect 480406 59200 480411 59256
rect 480210 59198 480411 59200
rect 483062 59258 483122 59334
rect 483289 59392 486023 59394
rect 483289 59336 483294 59392
rect 483350 59336 485962 59392
rect 486018 59336 486023 59392
rect 483289 59334 486023 59336
rect 483289 59331 483355 59334
rect 485957 59331 486023 59334
rect 487061 59394 487127 59397
rect 488533 59394 488599 59397
rect 487061 59392 488599 59394
rect 487061 59336 487066 59392
rect 487122 59336 488538 59392
rect 488594 59336 488599 59392
rect 487061 59334 488599 59336
rect 490208 59394 490268 60044
rect 491128 59530 491188 60044
rect 492140 59666 492200 60044
rect 492857 59666 492923 59669
rect 492140 59664 492923 59666
rect 492140 59608 492862 59664
rect 492918 59608 492923 59664
rect 492140 59606 492923 59608
rect 493060 59666 493120 60044
rect 493060 59606 493978 59666
rect 492857 59603 492923 59606
rect 492949 59530 493015 59533
rect 491128 59528 493015 59530
rect 491128 59472 492954 59528
rect 493010 59472 493015 59528
rect 491128 59470 493015 59472
rect 492949 59467 493015 59470
rect 492765 59394 492831 59397
rect 490208 59392 492831 59394
rect 490208 59336 492770 59392
rect 492826 59336 492831 59392
rect 490208 59334 492831 59336
rect 493918 59394 493978 59606
rect 494072 59530 494132 60044
rect 494992 59802 495052 60044
rect 496004 59938 496064 60044
rect 496004 59878 496922 59938
rect 495893 59802 495959 59805
rect 494992 59800 495959 59802
rect 494992 59744 495898 59800
rect 495954 59744 495959 59800
rect 494992 59742 495959 59744
rect 495893 59739 495959 59742
rect 494072 59470 495818 59530
rect 495525 59394 495591 59397
rect 493918 59392 495591 59394
rect 493918 59336 495530 59392
rect 495586 59336 495591 59392
rect 493918 59334 495591 59336
rect 487061 59331 487127 59334
rect 488533 59331 488599 59334
rect 492765 59331 492831 59334
rect 495525 59331 495591 59334
rect 483289 59258 483355 59261
rect 483062 59256 483355 59258
rect 483062 59200 483294 59256
rect 483350 59200 483355 59256
rect 483062 59198 483355 59200
rect 495758 59258 495818 59470
rect 496862 59394 496922 59878
rect 497016 59530 497076 60044
rect 497733 59530 497799 59533
rect 497016 59528 497799 59530
rect 497016 59472 497738 59528
rect 497794 59472 497799 59528
rect 497016 59470 497799 59472
rect 497936 59530 497996 60044
rect 498948 59666 499008 60044
rect 499868 59802 499928 60044
rect 500677 59802 500743 59805
rect 499868 59800 500743 59802
rect 499868 59744 500682 59800
rect 500738 59744 500743 59800
rect 499868 59742 500743 59744
rect 500677 59739 500743 59742
rect 498948 59606 500786 59666
rect 499849 59530 499915 59533
rect 497936 59528 499915 59530
rect 497936 59472 499854 59528
rect 499910 59472 499915 59528
rect 497936 59470 499915 59472
rect 497733 59467 497799 59470
rect 499849 59467 499915 59470
rect 498377 59394 498443 59397
rect 496862 59392 498443 59394
rect 496862 59336 498382 59392
rect 498438 59336 498443 59392
rect 496862 59334 498443 59336
rect 500726 59394 500786 59606
rect 500880 59530 500940 60044
rect 501892 59666 501952 60044
rect 502812 59802 502872 60044
rect 503621 59802 503687 59805
rect 502812 59800 503687 59802
rect 502812 59744 503626 59800
rect 503682 59744 503687 59800
rect 502812 59742 503687 59744
rect 503621 59739 503687 59742
rect 503621 59666 503687 59669
rect 501892 59664 503687 59666
rect 501892 59608 503626 59664
rect 503682 59608 503687 59664
rect 501892 59606 503687 59608
rect 503621 59603 503687 59606
rect 502425 59530 502491 59533
rect 500880 59528 502491 59530
rect 500880 59472 502430 59528
rect 502486 59472 502491 59528
rect 500880 59470 502491 59472
rect 502425 59467 502491 59470
rect 501045 59394 501111 59397
rect 500726 59392 501111 59394
rect 500726 59336 501050 59392
rect 501106 59336 501111 59392
rect 500726 59334 501111 59336
rect 503824 59394 503884 60044
rect 504744 59394 504804 60044
rect 505756 59394 505816 60044
rect 506676 59530 506736 60044
rect 507485 59530 507551 59533
rect 506676 59528 507551 59530
rect 506676 59472 507490 59528
rect 507546 59472 507551 59528
rect 506676 59470 507551 59472
rect 507485 59467 507551 59470
rect 507688 59394 507748 60044
rect 508700 59530 508760 60044
rect 509620 59666 509680 60044
rect 510632 59802 510692 60044
rect 511552 59938 511612 60044
rect 511552 59878 512378 59938
rect 510632 59742 512194 59802
rect 511993 59666 512059 59669
rect 509620 59664 512059 59666
rect 509620 59608 511998 59664
rect 512054 59608 512059 59664
rect 509620 59606 512059 59608
rect 511993 59603 512059 59606
rect 510613 59530 510679 59533
rect 508700 59528 510679 59530
rect 508700 59472 510618 59528
rect 510674 59472 510679 59528
rect 508700 59470 510679 59472
rect 510613 59467 510679 59470
rect 509601 59394 509667 59397
rect 503824 59334 504650 59394
rect 504744 59334 505570 59394
rect 505756 59334 507594 59394
rect 507688 59392 509667 59394
rect 507688 59336 509606 59392
rect 509662 59336 509667 59392
rect 507688 59334 509667 59336
rect 498377 59331 498443 59334
rect 501045 59331 501111 59334
rect 497089 59258 497155 59261
rect 495758 59256 497155 59258
rect 495758 59200 497094 59256
rect 497150 59200 497155 59256
rect 495758 59198 497155 59200
rect 451273 59195 451339 59198
rect 480345 59195 480411 59198
rect 483289 59195 483355 59198
rect 497089 59195 497155 59198
rect 440325 59122 440391 59125
rect 438166 59120 440391 59122
rect 438166 59064 440330 59120
rect 440386 59064 440391 59120
rect 438166 59062 440391 59064
rect 504590 59122 504650 59334
rect 505510 59258 505570 59334
rect 506749 59258 506815 59261
rect 505510 59256 506815 59258
rect 505510 59200 506754 59256
rect 506810 59200 506815 59256
rect 505510 59198 506815 59200
rect 507534 59258 507594 59334
rect 509601 59331 509667 59334
rect 507945 59258 508011 59261
rect 507534 59256 508011 59258
rect 507534 59200 507950 59256
rect 508006 59200 508011 59256
rect 507534 59198 508011 59200
rect 506749 59195 506815 59198
rect 507945 59195 508011 59198
rect 506565 59122 506631 59125
rect 504590 59120 506631 59122
rect 504590 59064 506570 59120
rect 506626 59064 506631 59120
rect 504590 59062 506631 59064
rect 512134 59122 512194 59742
rect 512318 59258 512378 59878
rect 512564 59394 512624 60044
rect 513484 59802 513544 60044
rect 514293 59802 514359 59805
rect 513484 59800 514359 59802
rect 513484 59744 514298 59800
rect 514354 59744 514359 59800
rect 513484 59742 514359 59744
rect 514293 59739 514359 59742
rect 514496 59530 514556 60044
rect 515508 59666 515568 60044
rect 516428 59802 516488 60044
rect 517237 59802 517303 59805
rect 516428 59800 517303 59802
rect 516428 59744 517242 59800
rect 517298 59744 517303 59800
rect 516428 59742 517303 59744
rect 517237 59739 517303 59742
rect 515508 59606 517346 59666
rect 516317 59530 516383 59533
rect 514496 59528 516383 59530
rect 514496 59472 516322 59528
rect 516378 59472 516383 59528
rect 514496 59470 516383 59472
rect 516317 59467 516383 59470
rect 514753 59394 514819 59397
rect 512564 59392 514819 59394
rect 512564 59336 514758 59392
rect 514814 59336 514819 59392
rect 512564 59334 514819 59336
rect 514753 59331 514819 59334
rect 514937 59394 515003 59397
rect 516501 59394 516567 59397
rect 514937 59392 516567 59394
rect 514937 59336 514942 59392
rect 514998 59336 516506 59392
rect 516562 59336 516567 59392
rect 514937 59334 516567 59336
rect 517286 59394 517346 59606
rect 517440 59530 517500 60044
rect 518360 59666 518420 60044
rect 518360 59606 519186 59666
rect 518985 59530 519051 59533
rect 517440 59528 519051 59530
rect 517440 59472 518990 59528
rect 519046 59472 519051 59528
rect 517440 59470 519051 59472
rect 518985 59467 519051 59470
rect 517513 59394 517579 59397
rect 517286 59392 517579 59394
rect 517286 59336 517518 59392
rect 517574 59336 517579 59392
rect 517286 59334 517579 59336
rect 519126 59394 519186 59606
rect 519372 59530 519432 60044
rect 520384 59666 520444 60044
rect 521304 59802 521364 60044
rect 522316 59938 522376 60044
rect 523236 59938 523296 60044
rect 522316 59878 523050 59938
rect 523236 59878 523970 59938
rect 522113 59802 522179 59805
rect 521304 59800 522179 59802
rect 521304 59744 522118 59800
rect 522174 59744 522179 59800
rect 521304 59742 522179 59744
rect 522113 59739 522179 59742
rect 520384 59606 522130 59666
rect 521653 59530 521719 59533
rect 519372 59528 521719 59530
rect 519372 59472 521658 59528
rect 521714 59472 521719 59528
rect 519372 59470 521719 59472
rect 521653 59467 521719 59470
rect 520365 59394 520431 59397
rect 519126 59392 520431 59394
rect 519126 59336 520370 59392
rect 520426 59336 520431 59392
rect 519126 59334 520431 59336
rect 522070 59394 522130 59606
rect 522990 59530 523050 59878
rect 523910 59802 523970 59878
rect 524045 59802 524111 59805
rect 523910 59800 524111 59802
rect 523910 59744 524050 59800
rect 524106 59744 524111 59800
rect 523910 59742 524111 59744
rect 524045 59739 524111 59742
rect 524248 59530 524308 60044
rect 525168 59666 525228 60044
rect 526180 59802 526240 60044
rect 526989 59802 527055 59805
rect 526180 59800 527055 59802
rect 526180 59744 526994 59800
rect 527050 59744 527055 59800
rect 526180 59742 527055 59744
rect 526989 59739 527055 59742
rect 525168 59606 527098 59666
rect 526621 59530 526687 59533
rect 522990 59470 523786 59530
rect 524248 59528 526687 59530
rect 524248 59472 526626 59528
rect 526682 59472 526687 59528
rect 524248 59470 526687 59472
rect 523726 59394 523786 59470
rect 526621 59467 526687 59470
rect 525057 59394 525123 59397
rect 522070 59334 523050 59394
rect 523726 59392 525123 59394
rect 523726 59336 525062 59392
rect 525118 59336 525123 59392
rect 523726 59334 525123 59336
rect 514937 59331 515003 59334
rect 516501 59331 516567 59334
rect 517513 59331 517579 59334
rect 520365 59331 520431 59334
rect 513649 59258 513715 59261
rect 512318 59256 513715 59258
rect 512318 59200 513654 59256
rect 513710 59200 513715 59256
rect 512318 59198 513715 59200
rect 522990 59258 523050 59334
rect 525057 59331 525123 59334
rect 523125 59258 523191 59261
rect 522990 59256 523191 59258
rect 522990 59200 523130 59256
rect 523186 59200 523191 59256
rect 522990 59198 523191 59200
rect 527038 59258 527098 59606
rect 527192 59394 527252 60044
rect 528112 59530 528172 60044
rect 529124 59666 529184 60044
rect 530044 59802 530104 60044
rect 530853 59802 530919 59805
rect 530044 59800 530919 59802
rect 530044 59744 530858 59800
rect 530914 59744 530919 59800
rect 530044 59742 530919 59744
rect 530853 59739 530919 59742
rect 529124 59606 530962 59666
rect 530761 59530 530827 59533
rect 528112 59528 530827 59530
rect 528112 59472 530766 59528
rect 530822 59472 530827 59528
rect 528112 59470 530827 59472
rect 530761 59467 530827 59470
rect 530577 59394 530643 59397
rect 527192 59392 530643 59394
rect 527192 59336 530582 59392
rect 530638 59336 530643 59392
rect 527192 59334 530643 59336
rect 530902 59394 530962 59606
rect 531056 59530 531116 60044
rect 532068 59666 532128 60044
rect 532988 59802 533048 60044
rect 533797 59802 533863 59805
rect 532988 59800 533863 59802
rect 532988 59744 533802 59800
rect 533858 59744 533863 59800
rect 532988 59742 533863 59744
rect 533797 59739 533863 59742
rect 532068 59606 533906 59666
rect 533337 59530 533403 59533
rect 531056 59528 533403 59530
rect 531056 59472 533342 59528
rect 533398 59472 533403 59528
rect 531056 59470 533403 59472
rect 533337 59467 533403 59470
rect 531957 59394 532023 59397
rect 530902 59392 532023 59394
rect 530902 59336 531962 59392
rect 532018 59336 532023 59392
rect 530902 59334 532023 59336
rect 533846 59394 533906 59606
rect 534000 59530 534060 60044
rect 534920 59666 534980 60044
rect 535932 59802 535992 60044
rect 535932 59742 537770 59802
rect 537477 59666 537543 59669
rect 534920 59664 537543 59666
rect 534920 59608 537482 59664
rect 537538 59608 537543 59664
rect 534920 59606 537543 59608
rect 537477 59603 537543 59606
rect 535729 59530 535795 59533
rect 534000 59528 535795 59530
rect 534000 59472 535734 59528
rect 535790 59472 535795 59528
rect 534000 59470 535795 59472
rect 535729 59467 535795 59470
rect 534717 59394 534783 59397
rect 533846 59392 534783 59394
rect 533846 59336 534722 59392
rect 534778 59336 534783 59392
rect 533846 59334 534783 59336
rect 537710 59394 537770 59742
rect 537864 59530 537924 60044
rect 538673 59530 538739 59533
rect 537864 59528 538739 59530
rect 537864 59472 538678 59528
rect 538734 59472 538739 59528
rect 537864 59470 538739 59472
rect 538876 59530 538936 60044
rect 539520 59666 539580 60044
rect 541617 59666 541683 59669
rect 539520 59664 541683 59666
rect 539520 59608 541622 59664
rect 541678 59608 541683 59664
rect 539520 59606 541683 59608
rect 541617 59603 541683 59606
rect 542261 59530 542327 59533
rect 538876 59528 542327 59530
rect 538876 59472 542266 59528
rect 542322 59472 542327 59528
rect 583520 59516 584960 59756
rect 538876 59470 542327 59472
rect 538673 59467 538739 59470
rect 542261 59467 542327 59470
rect 538857 59394 538923 59397
rect 537710 59392 538923 59394
rect 537710 59336 538862 59392
rect 538918 59336 538923 59392
rect 537710 59334 538923 59336
rect 530577 59331 530643 59334
rect 531957 59331 532023 59334
rect 534717 59331 534783 59334
rect 538857 59331 538923 59334
rect 539041 59394 539107 59397
rect 540237 59394 540303 59397
rect 539041 59392 540303 59394
rect 539041 59336 539046 59392
rect 539102 59336 540242 59392
rect 540298 59336 540303 59392
rect 539041 59334 540303 59336
rect 539041 59331 539107 59334
rect 540237 59331 540303 59334
rect 527817 59258 527883 59261
rect 527038 59256 527883 59258
rect 527038 59200 527822 59256
rect 527878 59200 527883 59256
rect 527038 59198 527883 59200
rect 513649 59195 513715 59198
rect 523125 59195 523191 59198
rect 527817 59195 527883 59198
rect 513465 59122 513531 59125
rect 512134 59120 513531 59122
rect 512134 59064 513470 59120
rect 513526 59064 513531 59120
rect 512134 59062 513531 59064
rect 421833 59059 421899 59062
rect 424133 59059 424199 59062
rect 440325 59059 440391 59062
rect 506565 59059 506631 59062
rect 513465 59059 513531 59062
rect -960 58564 480 58804
rect 583520 46188 584960 46428
rect -960 35036 480 35276
rect 583520 32996 584960 33236
rect 583520 19668 584960 19908
rect -960 11644 480 11884
rect 583520 6476 584960 6716
rect 494145 3634 494211 3637
rect 489870 3632 494211 3634
rect 489870 3576 494150 3632
rect 494206 3576 494211 3632
rect 489870 3574 494211 3576
rect 6453 3362 6519 3365
rect 159357 3362 159423 3365
rect 6453 3360 159423 3362
rect 6453 3304 6458 3360
rect 6514 3304 159362 3360
rect 159418 3304 159423 3360
rect 6453 3302 159423 3304
rect 6453 3299 6519 3302
rect 159357 3299 159423 3302
rect 418981 3362 419047 3365
rect 489870 3362 489930 3574
rect 494145 3571 494211 3574
rect 418981 3360 489930 3362
rect 418981 3304 418986 3360
rect 419042 3304 489930 3360
rect 418981 3302 489930 3304
rect 418981 3299 419047 3302
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 562004 60134 564618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 562004 63854 568338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 562004 67574 572058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 562004 74414 578898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 562004 78134 582618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 562004 81854 586338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 562004 85574 590058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 562004 92414 596898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 562004 96134 564618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 562004 99854 568338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 562004 103574 572058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 562004 110414 578898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 562004 114134 582618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 562004 117854 586338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 562004 121574 590058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 562004 128414 596898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 562004 132134 564618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 562004 135854 568338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 562004 139574 572058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 562004 146414 578898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 562004 150134 582618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 562004 153854 586338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 562004 157574 590058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 562004 164414 596898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 562004 168134 564618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 562004 171854 568338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 562004 175574 572058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 562004 182414 578898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 562004 186134 582618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 562004 189854 586338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 562004 193574 590058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 562004 200414 596898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 562004 204134 564618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 562004 207854 568338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 562004 211574 572058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 562004 218414 578898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 562004 222134 582618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 562004 225854 586338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 562004 229574 590058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 562004 236414 596898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 562004 240134 564618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 562004 243854 568338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 562004 247574 572058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 562004 254414 578898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 562004 258134 582618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 562004 261854 586338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 562004 265574 590058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 562004 272414 596898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 562004 276134 564618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 562004 279854 568338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 562004 283574 572058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 562004 290414 578898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 562004 294134 582618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 562004 297854 586338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 562004 301574 590058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 562004 308414 596898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 562004 312134 564618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 562004 315854 568338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 562004 319574 572058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 562004 326414 578898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 562004 330134 582618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 562004 333854 586338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 562004 337574 590058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 562004 344414 596898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 562004 348134 564618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 562004 351854 568338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 562004 355574 572058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 562004 362414 578898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 562004 366134 582618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 562004 369854 586338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 562004 373574 590058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 562004 380414 596898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 562004 384134 564618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 562004 387854 568338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 562004 391574 572058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 562004 398414 578898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 562004 402134 582618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 562004 405854 586338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 562004 409574 590058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 562004 416414 596898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 562004 420134 564618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 562004 423854 568338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 562004 427574 572058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 562004 434414 578898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 562004 438134 582618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 562004 441854 586338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 562004 445574 590058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 562004 452414 596898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 562004 456134 564618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 562004 459854 568338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 562004 463574 572058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 562004 470414 578898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 562004 474134 582618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 562004 477854 586338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 562004 481574 590058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 562004 488414 596898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 562004 492134 564618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 562004 495854 568338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 562004 499574 572058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 562004 506414 578898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 562004 510134 582618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 562004 513854 586338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 562004 517574 590058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 562004 524414 596898
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 562004 528134 564618
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 562004 531854 568338
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 562004 535574 572058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 562004 542414 578898
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 58000
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 28894 63854 58000
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 32614 67574 58000
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 39454 74414 58000
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 43174 78134 58000
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 46894 81854 58000
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 50614 85574 58000
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 58000
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 58000
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 28894 99854 58000
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 32614 103574 58000
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 39454 110414 58000
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 43174 114134 58000
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 46894 117854 58000
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 50614 121574 58000
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 58000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 58000
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 28894 135854 58000
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 32614 139574 58000
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 39454 146414 58000
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 43174 150134 58000
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 46894 153854 58000
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 50614 157574 58000
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 57454 164414 58000
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 25174 168134 58000
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 28894 171854 58000
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 32614 175574 58000
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 39454 182414 58000
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 43174 186134 58000
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 46894 189854 58000
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 50614 193574 58000
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 57454 200414 58000
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 58000
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 28894 207854 58000
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 32614 211574 58000
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 39454 218414 58000
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 43174 222134 58000
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 46894 225854 58000
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 50614 229574 58000
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 57454 236414 58000
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 58000
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 28894 243854 58000
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 32614 247574 58000
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 39454 254414 58000
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 43174 258134 58000
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 46894 261854 58000
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 50614 265574 58000
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 57454 272414 58000
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 25174 276134 58000
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 28894 279854 58000
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 32614 283574 58000
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 39454 290414 58000
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 43174 294134 58000
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 46894 297854 58000
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 50614 301574 58000
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 57454 308414 58000
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 25174 312134 58000
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 28894 315854 58000
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 32614 319574 58000
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 39454 326414 58000
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 43174 330134 58000
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 46894 333854 58000
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 50614 337574 58000
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 57454 344414 58000
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 25174 348134 58000
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 28894 351854 58000
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 32614 355574 58000
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 39454 362414 58000
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 43174 366134 58000
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 46894 369854 58000
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 50614 373574 58000
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 57454 380414 58000
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 25174 384134 58000
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 28894 387854 58000
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 32614 391574 58000
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 39454 398414 58000
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 43174 402134 58000
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 46894 405854 58000
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 50614 409574 58000
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 57454 416414 58000
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 25174 420134 58000
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 28894 423854 58000
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 32614 427574 58000
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 39454 434414 58000
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 43174 438134 58000
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 46894 441854 58000
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 50614 445574 58000
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 57454 452414 58000
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 25174 456134 58000
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 28894 459854 58000
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 32614 463574 58000
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 39454 470414 58000
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 43174 474134 58000
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 46894 477854 58000
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 50614 481574 58000
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 57454 488414 58000
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 25174 492134 58000
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 28894 495854 58000
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 32614 499574 58000
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 39454 506414 58000
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 43174 510134 58000
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 46894 513854 58000
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 50614 517574 58000
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 57454 524414 58000
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 25174 528134 58000
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 28894 531854 58000
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 32614 535574 58000
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 39454 542414 58000
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 58000 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 58000 561454
rect -2966 561134 58000 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 58000 561134
rect -2966 560866 58000 560898
rect 541964 561454 586890 561486
rect 541964 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 541964 561134 586890 561218
rect 541964 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 541964 560866 586890 560898
rect -8726 554614 58000 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 58000 554614
rect -8726 554294 58000 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 58000 554294
rect -8726 554026 58000 554058
rect 541964 554614 592650 554646
rect 541964 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect 541964 554294 592650 554378
rect 541964 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect 541964 554026 592650 554058
rect -6806 550894 58000 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 58000 550894
rect -6806 550574 58000 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 58000 550574
rect -6806 550306 58000 550338
rect 541964 550894 590730 550926
rect 541964 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect 541964 550574 590730 550658
rect 541964 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect 541964 550306 590730 550338
rect -4886 547174 58000 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 58000 547174
rect -4886 546854 58000 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 58000 546854
rect -4886 546586 58000 546618
rect 541964 547174 588810 547206
rect 541964 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect 541964 546854 588810 546938
rect 541964 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect 541964 546586 588810 546618
rect -2966 543454 58000 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 58000 543454
rect -2966 543134 58000 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 58000 543134
rect -2966 542866 58000 542898
rect 541964 543454 586890 543486
rect 541964 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect 541964 543134 586890 543218
rect 541964 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect 541964 542866 586890 542898
rect -8726 536614 58000 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 58000 536614
rect -8726 536294 58000 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 58000 536294
rect -8726 536026 58000 536058
rect 541964 536614 592650 536646
rect 541964 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 541964 536294 592650 536378
rect 541964 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 541964 536026 592650 536058
rect -6806 532894 58000 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 58000 532894
rect -6806 532574 58000 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 58000 532574
rect -6806 532306 58000 532338
rect 541964 532894 590730 532926
rect 541964 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 541964 532574 590730 532658
rect 541964 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 541964 532306 590730 532338
rect -4886 529174 58000 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 58000 529174
rect -4886 528854 58000 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 58000 528854
rect -4886 528586 58000 528618
rect 541964 529174 588810 529206
rect 541964 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 541964 528854 588810 528938
rect 541964 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 541964 528586 588810 528618
rect -2966 525454 58000 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 58000 525454
rect -2966 525134 58000 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 58000 525134
rect -2966 524866 58000 524898
rect 541964 525454 586890 525486
rect 541964 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 541964 525134 586890 525218
rect 541964 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 541964 524866 586890 524898
rect -8726 518614 58000 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 58000 518614
rect -8726 518294 58000 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 58000 518294
rect -8726 518026 58000 518058
rect 541964 518614 592650 518646
rect 541964 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect 541964 518294 592650 518378
rect 541964 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect 541964 518026 592650 518058
rect -6806 514894 58000 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 58000 514894
rect -6806 514574 58000 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 58000 514574
rect -6806 514306 58000 514338
rect 541964 514894 590730 514926
rect 541964 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect 541964 514574 590730 514658
rect 541964 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect 541964 514306 590730 514338
rect -4886 511174 58000 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 58000 511174
rect -4886 510854 58000 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 58000 510854
rect -4886 510586 58000 510618
rect 541964 511174 588810 511206
rect 541964 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect 541964 510854 588810 510938
rect 541964 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect 541964 510586 588810 510618
rect -2966 507454 58000 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 58000 507454
rect -2966 507134 58000 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 58000 507134
rect -2966 506866 58000 506898
rect 541964 507454 586890 507486
rect 541964 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect 541964 507134 586890 507218
rect 541964 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect 541964 506866 586890 506898
rect -8726 500614 58000 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 58000 500614
rect -8726 500294 58000 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 58000 500294
rect -8726 500026 58000 500058
rect 541964 500614 592650 500646
rect 541964 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 541964 500294 592650 500378
rect 541964 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 541964 500026 592650 500058
rect -6806 496894 58000 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 58000 496894
rect -6806 496574 58000 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 58000 496574
rect -6806 496306 58000 496338
rect 541964 496894 590730 496926
rect 541964 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 541964 496574 590730 496658
rect 541964 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 541964 496306 590730 496338
rect -4886 493174 58000 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 58000 493174
rect -4886 492854 58000 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 58000 492854
rect -4886 492586 58000 492618
rect 541964 493174 588810 493206
rect 541964 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 541964 492854 588810 492938
rect 541964 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 541964 492586 588810 492618
rect -2966 489454 58000 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 58000 489454
rect -2966 489134 58000 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 58000 489134
rect -2966 488866 58000 488898
rect 541964 489454 586890 489486
rect 541964 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 541964 489134 586890 489218
rect 541964 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 541964 488866 586890 488898
rect -8726 482614 58000 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 58000 482614
rect -8726 482294 58000 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 58000 482294
rect -8726 482026 58000 482058
rect 541964 482614 592650 482646
rect 541964 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect 541964 482294 592650 482378
rect 541964 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect 541964 482026 592650 482058
rect -6806 478894 58000 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 58000 478894
rect -6806 478574 58000 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 58000 478574
rect -6806 478306 58000 478338
rect 541964 478894 590730 478926
rect 541964 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect 541964 478574 590730 478658
rect 541964 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect 541964 478306 590730 478338
rect -4886 475174 58000 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 58000 475174
rect -4886 474854 58000 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 58000 474854
rect -4886 474586 58000 474618
rect 541964 475174 588810 475206
rect 541964 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect 541964 474854 588810 474938
rect 541964 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect 541964 474586 588810 474618
rect -2966 471454 58000 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 58000 471454
rect -2966 471134 58000 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 58000 471134
rect -2966 470866 58000 470898
rect 541964 471454 586890 471486
rect 541964 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect 541964 471134 586890 471218
rect 541964 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect 541964 470866 586890 470898
rect -8726 464614 58000 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 58000 464614
rect -8726 464294 58000 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 58000 464294
rect -8726 464026 58000 464058
rect 541964 464614 592650 464646
rect 541964 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 541964 464294 592650 464378
rect 541964 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 541964 464026 592650 464058
rect -6806 460894 58000 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 58000 460894
rect -6806 460574 58000 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 58000 460574
rect -6806 460306 58000 460338
rect 541964 460894 590730 460926
rect 541964 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 541964 460574 590730 460658
rect 541964 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 541964 460306 590730 460338
rect -4886 457174 58000 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 58000 457174
rect -4886 456854 58000 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 58000 456854
rect -4886 456586 58000 456618
rect 541964 457174 588810 457206
rect 541964 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 541964 456854 588810 456938
rect 541964 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 541964 456586 588810 456618
rect -2966 453454 58000 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 58000 453454
rect -2966 453134 58000 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 58000 453134
rect -2966 452866 58000 452898
rect 541964 453454 586890 453486
rect 541964 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 541964 453134 586890 453218
rect 541964 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 541964 452866 586890 452898
rect -8726 446614 58000 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 58000 446614
rect -8726 446294 58000 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 58000 446294
rect -8726 446026 58000 446058
rect 541964 446614 592650 446646
rect 541964 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect 541964 446294 592650 446378
rect 541964 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect 541964 446026 592650 446058
rect -6806 442894 58000 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 58000 442894
rect -6806 442574 58000 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 58000 442574
rect -6806 442306 58000 442338
rect 541964 442894 590730 442926
rect 541964 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect 541964 442574 590730 442658
rect 541964 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect 541964 442306 590730 442338
rect -4886 439174 58000 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 58000 439174
rect -4886 438854 58000 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 58000 438854
rect -4886 438586 58000 438618
rect 541964 439174 588810 439206
rect 541964 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect 541964 438854 588810 438938
rect 541964 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect 541964 438586 588810 438618
rect -2966 435454 58000 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 58000 435454
rect -2966 435134 58000 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 58000 435134
rect -2966 434866 58000 434898
rect 541964 435454 586890 435486
rect 541964 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect 541964 435134 586890 435218
rect 541964 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect 541964 434866 586890 434898
rect -8726 428614 58000 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 58000 428614
rect -8726 428294 58000 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 58000 428294
rect -8726 428026 58000 428058
rect 541964 428614 592650 428646
rect 541964 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 541964 428294 592650 428378
rect 541964 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 541964 428026 592650 428058
rect -6806 424894 58000 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 58000 424894
rect -6806 424574 58000 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 58000 424574
rect -6806 424306 58000 424338
rect 541964 424894 590730 424926
rect 541964 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 541964 424574 590730 424658
rect 541964 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 541964 424306 590730 424338
rect -4886 421174 58000 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 58000 421174
rect -4886 420854 58000 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 58000 420854
rect -4886 420586 58000 420618
rect 541964 421174 588810 421206
rect 541964 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 541964 420854 588810 420938
rect 541964 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 541964 420586 588810 420618
rect -2966 417454 58000 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 58000 417454
rect -2966 417134 58000 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 58000 417134
rect -2966 416866 58000 416898
rect 541964 417454 586890 417486
rect 541964 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 541964 417134 586890 417218
rect 541964 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 541964 416866 586890 416898
rect -8726 410614 58000 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 58000 410614
rect -8726 410294 58000 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 58000 410294
rect -8726 410026 58000 410058
rect 541964 410614 592650 410646
rect 541964 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect 541964 410294 592650 410378
rect 541964 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect 541964 410026 592650 410058
rect -6806 406894 58000 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 58000 406894
rect -6806 406574 58000 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 58000 406574
rect -6806 406306 58000 406338
rect 541964 406894 590730 406926
rect 541964 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect 541964 406574 590730 406658
rect 541964 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect 541964 406306 590730 406338
rect -4886 403174 58000 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 58000 403174
rect -4886 402854 58000 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 58000 402854
rect -4886 402586 58000 402618
rect 541964 403174 588810 403206
rect 541964 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect 541964 402854 588810 402938
rect 541964 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect 541964 402586 588810 402618
rect -2966 399454 58000 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 58000 399454
rect -2966 399134 58000 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 58000 399134
rect -2966 398866 58000 398898
rect 541964 399454 586890 399486
rect 541964 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect 541964 399134 586890 399218
rect 541964 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect 541964 398866 586890 398898
rect -8726 392614 58000 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 58000 392614
rect -8726 392294 58000 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 58000 392294
rect -8726 392026 58000 392058
rect 541964 392614 592650 392646
rect 541964 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 541964 392294 592650 392378
rect 541964 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 541964 392026 592650 392058
rect -6806 388894 58000 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 58000 388894
rect -6806 388574 58000 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 58000 388574
rect -6806 388306 58000 388338
rect 541964 388894 590730 388926
rect 541964 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 541964 388574 590730 388658
rect 541964 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 541964 388306 590730 388338
rect -4886 385174 58000 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 58000 385174
rect -4886 384854 58000 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 58000 384854
rect -4886 384586 58000 384618
rect 541964 385174 588810 385206
rect 541964 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 541964 384854 588810 384938
rect 541964 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 541964 384586 588810 384618
rect -2966 381454 58000 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 58000 381454
rect -2966 381134 58000 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 58000 381134
rect -2966 380866 58000 380898
rect 541964 381454 586890 381486
rect 541964 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 541964 381134 586890 381218
rect 541964 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 541964 380866 586890 380898
rect -8726 374614 58000 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 58000 374614
rect -8726 374294 58000 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 58000 374294
rect -8726 374026 58000 374058
rect 541964 374614 592650 374646
rect 541964 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect 541964 374294 592650 374378
rect 541964 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect 541964 374026 592650 374058
rect -6806 370894 58000 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 58000 370894
rect -6806 370574 58000 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 58000 370574
rect -6806 370306 58000 370338
rect 541964 370894 590730 370926
rect 541964 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect 541964 370574 590730 370658
rect 541964 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect 541964 370306 590730 370338
rect -4886 367174 58000 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 58000 367174
rect -4886 366854 58000 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 58000 366854
rect -4886 366586 58000 366618
rect 541964 367174 588810 367206
rect 541964 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect 541964 366854 588810 366938
rect 541964 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect 541964 366586 588810 366618
rect -2966 363454 58000 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 58000 363454
rect -2966 363134 58000 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 58000 363134
rect -2966 362866 58000 362898
rect 541964 363454 586890 363486
rect 541964 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect 541964 363134 586890 363218
rect 541964 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect 541964 362866 586890 362898
rect -8726 356614 58000 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 58000 356614
rect -8726 356294 58000 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 58000 356294
rect -8726 356026 58000 356058
rect 541964 356614 592650 356646
rect 541964 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 541964 356294 592650 356378
rect 541964 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 541964 356026 592650 356058
rect -6806 352894 58000 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 58000 352894
rect -6806 352574 58000 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 58000 352574
rect -6806 352306 58000 352338
rect 541964 352894 590730 352926
rect 541964 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 541964 352574 590730 352658
rect 541964 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 541964 352306 590730 352338
rect -4886 349174 58000 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 58000 349174
rect -4886 348854 58000 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 58000 348854
rect -4886 348586 58000 348618
rect 541964 349174 588810 349206
rect 541964 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 541964 348854 588810 348938
rect 541964 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 541964 348586 588810 348618
rect -2966 345454 58000 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 58000 345454
rect -2966 345134 58000 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 58000 345134
rect -2966 344866 58000 344898
rect 541964 345454 586890 345486
rect 541964 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 541964 345134 586890 345218
rect 541964 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 541964 344866 586890 344898
rect -8726 338614 58000 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 58000 338614
rect -8726 338294 58000 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 58000 338294
rect -8726 338026 58000 338058
rect 541964 338614 592650 338646
rect 541964 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect 541964 338294 592650 338378
rect 541964 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect 541964 338026 592650 338058
rect -6806 334894 58000 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 58000 334894
rect -6806 334574 58000 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 58000 334574
rect -6806 334306 58000 334338
rect 541964 334894 590730 334926
rect 541964 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect 541964 334574 590730 334658
rect 541964 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect 541964 334306 590730 334338
rect -4886 331174 58000 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 58000 331174
rect -4886 330854 58000 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 58000 330854
rect -4886 330586 58000 330618
rect 541964 331174 588810 331206
rect 541964 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect 541964 330854 588810 330938
rect 541964 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect 541964 330586 588810 330618
rect -2966 327454 58000 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 58000 327454
rect -2966 327134 58000 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 58000 327134
rect -2966 326866 58000 326898
rect 541964 327454 586890 327486
rect 541964 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect 541964 327134 586890 327218
rect 541964 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect 541964 326866 586890 326898
rect -8726 320614 58000 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 58000 320614
rect -8726 320294 58000 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 58000 320294
rect -8726 320026 58000 320058
rect 541964 320614 592650 320646
rect 541964 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 541964 320294 592650 320378
rect 541964 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 541964 320026 592650 320058
rect -6806 316894 58000 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 58000 316894
rect -6806 316574 58000 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 58000 316574
rect -6806 316306 58000 316338
rect 541964 316894 590730 316926
rect 541964 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 541964 316574 590730 316658
rect 541964 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 541964 316306 590730 316338
rect -4886 313174 58000 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 58000 313174
rect -4886 312854 58000 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 58000 312854
rect -4886 312586 58000 312618
rect 541964 313174 588810 313206
rect 541964 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 541964 312854 588810 312938
rect 541964 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 541964 312586 588810 312618
rect -2966 309454 58000 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 58000 309454
rect -2966 309134 58000 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 58000 309134
rect -2966 308866 58000 308898
rect 541964 309454 586890 309486
rect 541964 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 541964 309134 586890 309218
rect 541964 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 541964 308866 586890 308898
rect -8726 302614 58000 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 58000 302614
rect -8726 302294 58000 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 58000 302294
rect -8726 302026 58000 302058
rect 541964 302614 592650 302646
rect 541964 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect 541964 302294 592650 302378
rect 541964 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect 541964 302026 592650 302058
rect -6806 298894 58000 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 58000 298894
rect -6806 298574 58000 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 58000 298574
rect -6806 298306 58000 298338
rect 541964 298894 590730 298926
rect 541964 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect 541964 298574 590730 298658
rect 541964 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect 541964 298306 590730 298338
rect -4886 295174 58000 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 58000 295174
rect -4886 294854 58000 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 58000 294854
rect -4886 294586 58000 294618
rect 541964 295174 588810 295206
rect 541964 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect 541964 294854 588810 294938
rect 541964 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect 541964 294586 588810 294618
rect -2966 291454 58000 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 58000 291454
rect -2966 291134 58000 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 58000 291134
rect -2966 290866 58000 290898
rect 541964 291454 586890 291486
rect 541964 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect 541964 291134 586890 291218
rect 541964 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect 541964 290866 586890 290898
rect -8726 284614 58000 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 58000 284614
rect -8726 284294 58000 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 58000 284294
rect -8726 284026 58000 284058
rect 541964 284614 592650 284646
rect 541964 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 541964 284294 592650 284378
rect 541964 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 541964 284026 592650 284058
rect -6806 280894 58000 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 58000 280894
rect -6806 280574 58000 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 58000 280574
rect -6806 280306 58000 280338
rect 541964 280894 590730 280926
rect 541964 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 541964 280574 590730 280658
rect 541964 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 541964 280306 590730 280338
rect -4886 277174 58000 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 58000 277174
rect -4886 276854 58000 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 58000 276854
rect -4886 276586 58000 276618
rect 541964 277174 588810 277206
rect 541964 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 541964 276854 588810 276938
rect 541964 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 541964 276586 588810 276618
rect -2966 273454 58000 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 58000 273454
rect -2966 273134 58000 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 58000 273134
rect -2966 272866 58000 272898
rect 541964 273454 586890 273486
rect 541964 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 541964 273134 586890 273218
rect 541964 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 541964 272866 586890 272898
rect -8726 266614 58000 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 58000 266614
rect -8726 266294 58000 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 58000 266294
rect -8726 266026 58000 266058
rect 541964 266614 592650 266646
rect 541964 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect 541964 266294 592650 266378
rect 541964 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect 541964 266026 592650 266058
rect -6806 262894 58000 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 58000 262894
rect -6806 262574 58000 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 58000 262574
rect -6806 262306 58000 262338
rect 541964 262894 590730 262926
rect 541964 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect 541964 262574 590730 262658
rect 541964 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect 541964 262306 590730 262338
rect -4886 259174 58000 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 58000 259174
rect -4886 258854 58000 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 58000 258854
rect -4886 258586 58000 258618
rect 541964 259174 588810 259206
rect 541964 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect 541964 258854 588810 258938
rect 541964 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect 541964 258586 588810 258618
rect -2966 255454 58000 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 58000 255454
rect -2966 255134 58000 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 58000 255134
rect -2966 254866 58000 254898
rect 541964 255454 586890 255486
rect 541964 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect 541964 255134 586890 255218
rect 541964 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect 541964 254866 586890 254898
rect -8726 248614 58000 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 58000 248614
rect -8726 248294 58000 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 58000 248294
rect -8726 248026 58000 248058
rect 541964 248614 592650 248646
rect 541964 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 541964 248294 592650 248378
rect 541964 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 541964 248026 592650 248058
rect -6806 244894 58000 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 58000 244894
rect -6806 244574 58000 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 58000 244574
rect -6806 244306 58000 244338
rect 541964 244894 590730 244926
rect 541964 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 541964 244574 590730 244658
rect 541964 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 541964 244306 590730 244338
rect -4886 241174 58000 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 58000 241174
rect -4886 240854 58000 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 58000 240854
rect -4886 240586 58000 240618
rect 541964 241174 588810 241206
rect 541964 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 541964 240854 588810 240938
rect 541964 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 541964 240586 588810 240618
rect -2966 237454 58000 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 58000 237454
rect -2966 237134 58000 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 58000 237134
rect -2966 236866 58000 236898
rect 541964 237454 586890 237486
rect 541964 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 541964 237134 586890 237218
rect 541964 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 541964 236866 586890 236898
rect -8726 230614 58000 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 58000 230614
rect -8726 230294 58000 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 58000 230294
rect -8726 230026 58000 230058
rect 541964 230614 592650 230646
rect 541964 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect 541964 230294 592650 230378
rect 541964 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect 541964 230026 592650 230058
rect -6806 226894 58000 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 58000 226894
rect -6806 226574 58000 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 58000 226574
rect -6806 226306 58000 226338
rect 541964 226894 590730 226926
rect 541964 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect 541964 226574 590730 226658
rect 541964 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect 541964 226306 590730 226338
rect -4886 223174 58000 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 58000 223174
rect -4886 222854 58000 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 58000 222854
rect -4886 222586 58000 222618
rect 541964 223174 588810 223206
rect 541964 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect 541964 222854 588810 222938
rect 541964 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect 541964 222586 588810 222618
rect -2966 219454 58000 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 58000 219454
rect -2966 219134 58000 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 58000 219134
rect -2966 218866 58000 218898
rect 541964 219454 586890 219486
rect 541964 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect 541964 219134 586890 219218
rect 541964 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect 541964 218866 586890 218898
rect -8726 212614 58000 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 58000 212614
rect -8726 212294 58000 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 58000 212294
rect -8726 212026 58000 212058
rect 541964 212614 592650 212646
rect 541964 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 541964 212294 592650 212378
rect 541964 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 541964 212026 592650 212058
rect -6806 208894 58000 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 58000 208894
rect -6806 208574 58000 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 58000 208574
rect -6806 208306 58000 208338
rect 541964 208894 590730 208926
rect 541964 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 541964 208574 590730 208658
rect 541964 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 541964 208306 590730 208338
rect -4886 205174 58000 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 58000 205174
rect -4886 204854 58000 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 58000 204854
rect -4886 204586 58000 204618
rect 541964 205174 588810 205206
rect 541964 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 541964 204854 588810 204938
rect 541964 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 541964 204586 588810 204618
rect -2966 201454 58000 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 58000 201454
rect -2966 201134 58000 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 58000 201134
rect -2966 200866 58000 200898
rect 541964 201454 586890 201486
rect 541964 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 541964 201134 586890 201218
rect 541964 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 541964 200866 586890 200898
rect -8726 194614 58000 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 58000 194614
rect -8726 194294 58000 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 58000 194294
rect -8726 194026 58000 194058
rect 541964 194614 592650 194646
rect 541964 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect 541964 194294 592650 194378
rect 541964 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect 541964 194026 592650 194058
rect -6806 190894 58000 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 58000 190894
rect -6806 190574 58000 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 58000 190574
rect -6806 190306 58000 190338
rect 541964 190894 590730 190926
rect 541964 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect 541964 190574 590730 190658
rect 541964 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect 541964 190306 590730 190338
rect -4886 187174 58000 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 58000 187174
rect -4886 186854 58000 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 58000 186854
rect -4886 186586 58000 186618
rect 541964 187174 588810 187206
rect 541964 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect 541964 186854 588810 186938
rect 541964 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect 541964 186586 588810 186618
rect -2966 183454 58000 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 58000 183454
rect -2966 183134 58000 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 58000 183134
rect -2966 182866 58000 182898
rect 541964 183454 586890 183486
rect 541964 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect 541964 183134 586890 183218
rect 541964 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect 541964 182866 586890 182898
rect -8726 176614 58000 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 58000 176614
rect -8726 176294 58000 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 58000 176294
rect -8726 176026 58000 176058
rect 541964 176614 592650 176646
rect 541964 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 541964 176294 592650 176378
rect 541964 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 541964 176026 592650 176058
rect -6806 172894 58000 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 58000 172894
rect -6806 172574 58000 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 58000 172574
rect -6806 172306 58000 172338
rect 541964 172894 590730 172926
rect 541964 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 541964 172574 590730 172658
rect 541964 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 541964 172306 590730 172338
rect -4886 169174 58000 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 58000 169174
rect -4886 168854 58000 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 58000 168854
rect -4886 168586 58000 168618
rect 541964 169174 588810 169206
rect 541964 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 541964 168854 588810 168938
rect 541964 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 541964 168586 588810 168618
rect -2966 165454 58000 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 58000 165454
rect -2966 165134 58000 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 58000 165134
rect -2966 164866 58000 164898
rect 541964 165454 586890 165486
rect 541964 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 541964 165134 586890 165218
rect 541964 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 541964 164866 586890 164898
rect -8726 158614 58000 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 58000 158614
rect -8726 158294 58000 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 58000 158294
rect -8726 158026 58000 158058
rect 541964 158614 592650 158646
rect 541964 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect 541964 158294 592650 158378
rect 541964 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect 541964 158026 592650 158058
rect -6806 154894 58000 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 58000 154894
rect -6806 154574 58000 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 58000 154574
rect -6806 154306 58000 154338
rect 541964 154894 590730 154926
rect 541964 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect 541964 154574 590730 154658
rect 541964 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect 541964 154306 590730 154338
rect -4886 151174 58000 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 58000 151174
rect -4886 150854 58000 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 58000 150854
rect -4886 150586 58000 150618
rect 541964 151174 588810 151206
rect 541964 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect 541964 150854 588810 150938
rect 541964 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect 541964 150586 588810 150618
rect -2966 147454 58000 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 58000 147454
rect -2966 147134 58000 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 58000 147134
rect -2966 146866 58000 146898
rect 541964 147454 586890 147486
rect 541964 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect 541964 147134 586890 147218
rect 541964 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect 541964 146866 586890 146898
rect -8726 140614 58000 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 58000 140614
rect -8726 140294 58000 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 58000 140294
rect -8726 140026 58000 140058
rect 541964 140614 592650 140646
rect 541964 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 541964 140294 592650 140378
rect 541964 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 541964 140026 592650 140058
rect -6806 136894 58000 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 58000 136894
rect -6806 136574 58000 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 58000 136574
rect -6806 136306 58000 136338
rect 541964 136894 590730 136926
rect 541964 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 541964 136574 590730 136658
rect 541964 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 541964 136306 590730 136338
rect -4886 133174 58000 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 58000 133174
rect -4886 132854 58000 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 58000 132854
rect -4886 132586 58000 132618
rect 541964 133174 588810 133206
rect 541964 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 541964 132854 588810 132938
rect 541964 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 541964 132586 588810 132618
rect -2966 129454 58000 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 58000 129454
rect -2966 129134 58000 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 58000 129134
rect -2966 128866 58000 128898
rect 541964 129454 586890 129486
rect 541964 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 541964 129134 586890 129218
rect 541964 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 541964 128866 586890 128898
rect -8726 122614 58000 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 58000 122614
rect -8726 122294 58000 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 58000 122294
rect -8726 122026 58000 122058
rect 541964 122614 592650 122646
rect 541964 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect 541964 122294 592650 122378
rect 541964 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect 541964 122026 592650 122058
rect -6806 118894 58000 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 58000 118894
rect -6806 118574 58000 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 58000 118574
rect -6806 118306 58000 118338
rect 541964 118894 590730 118926
rect 541964 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect 541964 118574 590730 118658
rect 541964 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect 541964 118306 590730 118338
rect -4886 115174 58000 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 58000 115174
rect -4886 114854 58000 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 58000 114854
rect -4886 114586 58000 114618
rect 541964 115174 588810 115206
rect 541964 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect 541964 114854 588810 114938
rect 541964 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect 541964 114586 588810 114618
rect -2966 111454 58000 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 58000 111454
rect -2966 111134 58000 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 58000 111134
rect -2966 110866 58000 110898
rect 541964 111454 586890 111486
rect 541964 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect 541964 111134 586890 111218
rect 541964 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect 541964 110866 586890 110898
rect -8726 104614 58000 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 58000 104614
rect -8726 104294 58000 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 58000 104294
rect -8726 104026 58000 104058
rect 541964 104614 592650 104646
rect 541964 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 541964 104294 592650 104378
rect 541964 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 541964 104026 592650 104058
rect -6806 100894 58000 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 58000 100894
rect -6806 100574 58000 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 58000 100574
rect -6806 100306 58000 100338
rect 541964 100894 590730 100926
rect 541964 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 541964 100574 590730 100658
rect 541964 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 541964 100306 590730 100338
rect -4886 97174 58000 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 58000 97174
rect -4886 96854 58000 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 58000 96854
rect -4886 96586 58000 96618
rect 541964 97174 588810 97206
rect 541964 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 541964 96854 588810 96938
rect 541964 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 541964 96586 588810 96618
rect -2966 93454 58000 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 58000 93454
rect -2966 93134 58000 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 58000 93134
rect -2966 92866 58000 92898
rect 541964 93454 586890 93486
rect 541964 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 541964 93134 586890 93218
rect 541964 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 541964 92866 586890 92898
rect -8726 86614 58000 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 58000 86614
rect -8726 86294 58000 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 58000 86294
rect -8726 86026 58000 86058
rect 541964 86614 592650 86646
rect 541964 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect 541964 86294 592650 86378
rect 541964 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect 541964 86026 592650 86058
rect -6806 82894 58000 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 58000 82894
rect -6806 82574 58000 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 58000 82574
rect -6806 82306 58000 82338
rect 541964 82894 590730 82926
rect 541964 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect 541964 82574 590730 82658
rect 541964 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect 541964 82306 590730 82338
rect -4886 79174 58000 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 58000 79174
rect -4886 78854 58000 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 58000 78854
rect -4886 78586 58000 78618
rect 541964 79174 588810 79206
rect 541964 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect 541964 78854 588810 78938
rect 541964 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect 541964 78586 588810 78618
rect -2966 75454 58000 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 58000 75454
rect -2966 75134 58000 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 58000 75134
rect -2966 74866 58000 74898
rect 541964 75454 586890 75486
rect 541964 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect 541964 75134 586890 75218
rect 541964 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect 541964 74866 586890 74898
rect -8726 68614 58000 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 58000 68614
rect -8726 68294 58000 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 58000 68294
rect -8726 68026 58000 68058
rect 541964 68614 592650 68646
rect 541964 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 541964 68294 592650 68378
rect 541964 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 541964 68026 592650 68058
rect -6806 64894 58000 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 58000 64894
rect -6806 64574 58000 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 58000 64574
rect -6806 64306 58000 64338
rect 541964 64894 590730 64926
rect 541964 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 541964 64574 590730 64658
rect 541964 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 541964 64306 590730 64338
rect -4886 61174 58000 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 58000 61174
rect -4886 60854 58000 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 58000 60854
rect -4886 60586 58000 60618
rect 541964 61174 588810 61206
rect 541964 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 541964 60854 588810 60938
rect 541964 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 541964 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use azadi_soc_top_caravel  mprj
timestamp 0
transform 1 0 60000 0 1 60000
box 0 0 479964 500004
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 692052 480 692292 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 598212 480 598452 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 504372 480 504612 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 410532 480 410772 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 316556 480 316796 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 222716 480 222956 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 15 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 16 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 17 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 18 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 19 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 20 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 21 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 23 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 24 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 25 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 26 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 27 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 28 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 29 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 30 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 31 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 32 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 33 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 34 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 35 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 36 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 37 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 38 nsew signal input
rlabel metal3 s -960 668524 480 668764 4 io_in[24]
port 39 nsew signal input
rlabel metal3 s -960 574684 480 574924 4 io_in[25]
port 40 nsew signal input
rlabel metal3 s -960 480844 480 481084 4 io_in[26]
port 41 nsew signal input
rlabel metal3 s -960 387004 480 387244 4 io_in[27]
port 42 nsew signal input
rlabel metal3 s -960 293164 480 293404 4 io_in[28]
port 43 nsew signal input
rlabel metal3 s -960 199324 480 199564 4 io_in[29]
port 44 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 45 nsew signal input
rlabel metal3 s -960 128876 480 129116 4 io_in[30]
port 46 nsew signal input
rlabel metal3 s -960 58564 480 58804 4 io_in[31]
port 47 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 48 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 49 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 50 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 51 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 52 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 53 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 54 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 55 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 56 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 57 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 58 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 59 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 60 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 61 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 62 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 63 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 64 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 65 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 66 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 67 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 68 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 69 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 70 nsew signal tristate
rlabel metal3 s -960 621604 480 621844 4 io_oeb[24]
port 71 nsew signal tristate
rlabel metal3 s -960 527764 480 528004 4 io_oeb[25]
port 72 nsew signal tristate
rlabel metal3 s -960 433924 480 434164 4 io_oeb[26]
port 73 nsew signal tristate
rlabel metal3 s -960 340084 480 340324 4 io_oeb[27]
port 74 nsew signal tristate
rlabel metal3 s -960 246244 480 246484 4 io_oeb[28]
port 75 nsew signal tristate
rlabel metal3 s -960 152404 480 152644 4 io_oeb[29]
port 76 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 77 nsew signal tristate
rlabel metal3 s -960 81956 480 82196 4 io_oeb[30]
port 78 nsew signal tristate
rlabel metal3 s -960 11644 480 11884 4 io_oeb[31]
port 79 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 80 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 81 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 82 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 83 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 84 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 85 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 86 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 87 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 88 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 89 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 90 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 91 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 92 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 93 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 94 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 95 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 96 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 97 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 98 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 99 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 100 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 101 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 102 nsew signal tristate
rlabel metal3 s -960 645132 480 645372 4 io_out[24]
port 103 nsew signal tristate
rlabel metal3 s -960 551292 480 551532 4 io_out[25]
port 104 nsew signal tristate
rlabel metal3 s -960 457452 480 457692 4 io_out[26]
port 105 nsew signal tristate
rlabel metal3 s -960 363612 480 363852 4 io_out[27]
port 106 nsew signal tristate
rlabel metal3 s -960 269636 480 269876 4 io_out[28]
port 107 nsew signal tristate
rlabel metal3 s -960 175796 480 176036 4 io_out[29]
port 108 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 109 nsew signal tristate
rlabel metal3 s -960 105484 480 105724 4 io_out[30]
port 110 nsew signal tristate
rlabel metal3 s -960 35036 480 35276 4 io_out[31]
port 111 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 112 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 113 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 114 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 115 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 116 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 117 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 118 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 119 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 120 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 121 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 122 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 123 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 124 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 125 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 126 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 127 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 128 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 129 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 130 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 131 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 132 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 133 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 134 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 135 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 136 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 137 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 138 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 139 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 140 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 141 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 142 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 143 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 144 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 145 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 146 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 147 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 148 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 149 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 150 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 151 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 152 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 153 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 154 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 155 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 156 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 157 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 158 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 159 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 160 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 161 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 162 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 163 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 164 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 165 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 166 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 167 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 168 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 169 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 170 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 171 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 172 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 173 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 174 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 175 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 176 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 177 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 178 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 179 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 180 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 181 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 182 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 183 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 184 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 185 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 186 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 187 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 188 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 189 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 190 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 191 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 192 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 193 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 194 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 195 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 196 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 197 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 198 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 199 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 200 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 201 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 202 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 203 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 204 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 205 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 206 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 207 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 208 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 209 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 210 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 211 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 212 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 213 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 214 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 215 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 216 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 217 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 218 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 219 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 220 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 221 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 222 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 223 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 224 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 225 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 226 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 227 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 228 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 229 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 230 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 231 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 232 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 233 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 234 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 235 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 236 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 237 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 238 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 239 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 240 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 241 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 242 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 243 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 244 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 245 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 246 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 247 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 248 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 249 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 250 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 251 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 252 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 253 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 254 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 255 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 256 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 257 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 258 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 259 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 260 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 261 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 262 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 263 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 264 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 265 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 266 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 267 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 268 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 269 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 270 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 271 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 272 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 273 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 274 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 275 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 276 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 277 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 278 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 279 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 280 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 281 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 282 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 283 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 284 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 285 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 286 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 287 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 288 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 289 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 290 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 291 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 292 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 293 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 294 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 295 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 296 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 297 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 298 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 299 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 300 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 301 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 302 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 303 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 304 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 305 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 306 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 307 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 308 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 309 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 310 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 311 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 312 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 313 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 314 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 315 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 316 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 317 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 318 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 319 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 320 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 321 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 322 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 323 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 324 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 325 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 326 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 327 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 328 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 329 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 330 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 331 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 332 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 333 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 334 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 335 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 336 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 337 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 338 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 339 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 340 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 341 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 342 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 343 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 344 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 345 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 346 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 347 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 348 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 349 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 350 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 351 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 352 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 353 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 354 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 355 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 356 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 357 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 358 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 359 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 360 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 361 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 362 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 363 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 364 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 365 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 366 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 367 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 368 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 369 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 370 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 371 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 372 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 373 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 374 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 375 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 376 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 377 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 378 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 379 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 380 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 381 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 382 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 383 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 384 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 385 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 386 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 387 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 388 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 389 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 390 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 391 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 392 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 393 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 394 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 395 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 396 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 397 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 398 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 399 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 400 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 401 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 402 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 403 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 404 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 405 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 406 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 407 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 408 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 409 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 410 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 411 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 412 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 413 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 414 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 415 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 416 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 417 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 418 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 419 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 420 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 421 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 422 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 423 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 424 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 425 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 426 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 427 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 428 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 429 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 430 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 431 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 432 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 433 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 434 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 435 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 436 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 437 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 438 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 439 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 440 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 441 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 442 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 443 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 444 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 445 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 446 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 447 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 448 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 449 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 450 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 451 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 452 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 453 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 454 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 455 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 456 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 457 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 458 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 459 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 460 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 461 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 462 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 463 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 464 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 465 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 466 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 467 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 468 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 469 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 470 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 471 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 472 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 473 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 474 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 475 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 476 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 477 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 478 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 479 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 480 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 481 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 482 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 483 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 484 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 485 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 486 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 487 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 488 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 489 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 490 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 491 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 492 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 493 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 494 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 495 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 496 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 497 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 498 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 499 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 500 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 501 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 502 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 503 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 504 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 505 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 506 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 507 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 74866 58000 75486 6 vccd1
port 507 nsew power input
rlabel metal5 s 541964 74866 586890 75486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 110866 58000 111486 6 vccd1
port 507 nsew power input
rlabel metal5 s 541964 110866 586890 111486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 146866 58000 147486 6 vccd1
port 507 nsew power input
rlabel metal5 s 541964 146866 586890 147486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 182866 58000 183486 6 vccd1
port 507 nsew power input
rlabel metal5 s 541964 182866 586890 183486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 218866 58000 219486 6 vccd1
port 507 nsew power input
rlabel metal5 s 541964 218866 586890 219486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 254866 58000 255486 6 vccd1
port 507 nsew power input
rlabel metal5 s 541964 254866 586890 255486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 290866 58000 291486 6 vccd1
port 507 nsew power input
rlabel metal5 s 541964 290866 586890 291486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 326866 58000 327486 6 vccd1
port 507 nsew power input
rlabel metal5 s 541964 326866 586890 327486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 362866 58000 363486 6 vccd1
port 507 nsew power input
rlabel metal5 s 541964 362866 586890 363486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 398866 58000 399486 6 vccd1
port 507 nsew power input
rlabel metal5 s 541964 398866 586890 399486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 434866 58000 435486 6 vccd1
port 507 nsew power input
rlabel metal5 s 541964 434866 586890 435486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 470866 58000 471486 6 vccd1
port 507 nsew power input
rlabel metal5 s 541964 470866 586890 471486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 506866 58000 507486 6 vccd1
port 507 nsew power input
rlabel metal5 s 541964 506866 586890 507486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 542866 58000 543486 6 vccd1
port 507 nsew power input
rlabel metal5 s 541964 542866 586890 543486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 507 nsew power input
rlabel metal4 s 73794 -1894 74414 58000 6 vccd1
port 507 nsew power input
rlabel metal4 s 109794 -1894 110414 58000 6 vccd1
port 507 nsew power input
rlabel metal4 s 145794 -1894 146414 58000 6 vccd1
port 507 nsew power input
rlabel metal4 s 181794 -1894 182414 58000 6 vccd1
port 507 nsew power input
rlabel metal4 s 217794 -1894 218414 58000 6 vccd1
port 507 nsew power input
rlabel metal4 s 253794 -1894 254414 58000 6 vccd1
port 507 nsew power input
rlabel metal4 s 289794 -1894 290414 58000 6 vccd1
port 507 nsew power input
rlabel metal4 s 325794 -1894 326414 58000 6 vccd1
port 507 nsew power input
rlabel metal4 s 361794 -1894 362414 58000 6 vccd1
port 507 nsew power input
rlabel metal4 s 397794 -1894 398414 58000 6 vccd1
port 507 nsew power input
rlabel metal4 s 433794 -1894 434414 58000 6 vccd1
port 507 nsew power input
rlabel metal4 s 469794 -1894 470414 58000 6 vccd1
port 507 nsew power input
rlabel metal4 s 505794 -1894 506414 58000 6 vccd1
port 507 nsew power input
rlabel metal4 s 541794 -1894 542414 58000 6 vccd1
port 507 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 507 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 507 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 73794 562004 74414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 109794 562004 110414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 145794 562004 146414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 181794 562004 182414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 217794 562004 218414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 253794 562004 254414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 289794 562004 290414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 325794 562004 326414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 361794 562004 362414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 397794 562004 398414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 433794 562004 434414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 469794 562004 470414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 505794 562004 506414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 541794 562004 542414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 507 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 508 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 78586 58000 79206 6 vccd2
port 508 nsew power input
rlabel metal5 s 541964 78586 588810 79206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 114586 58000 115206 6 vccd2
port 508 nsew power input
rlabel metal5 s 541964 114586 588810 115206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 150586 58000 151206 6 vccd2
port 508 nsew power input
rlabel metal5 s 541964 150586 588810 151206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 186586 58000 187206 6 vccd2
port 508 nsew power input
rlabel metal5 s 541964 186586 588810 187206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 222586 58000 223206 6 vccd2
port 508 nsew power input
rlabel metal5 s 541964 222586 588810 223206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 258586 58000 259206 6 vccd2
port 508 nsew power input
rlabel metal5 s 541964 258586 588810 259206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 294586 58000 295206 6 vccd2
port 508 nsew power input
rlabel metal5 s 541964 294586 588810 295206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 330586 58000 331206 6 vccd2
port 508 nsew power input
rlabel metal5 s 541964 330586 588810 331206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 366586 58000 367206 6 vccd2
port 508 nsew power input
rlabel metal5 s 541964 366586 588810 367206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 402586 58000 403206 6 vccd2
port 508 nsew power input
rlabel metal5 s 541964 402586 588810 403206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 438586 58000 439206 6 vccd2
port 508 nsew power input
rlabel metal5 s 541964 438586 588810 439206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 474586 58000 475206 6 vccd2
port 508 nsew power input
rlabel metal5 s 541964 474586 588810 475206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 510586 58000 511206 6 vccd2
port 508 nsew power input
rlabel metal5 s 541964 510586 588810 511206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 546586 58000 547206 6 vccd2
port 508 nsew power input
rlabel metal5 s 541964 546586 588810 547206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 508 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 508 nsew power input
rlabel metal4 s 77514 -3814 78134 58000 6 vccd2
port 508 nsew power input
rlabel metal4 s 113514 -3814 114134 58000 6 vccd2
port 508 nsew power input
rlabel metal4 s 149514 -3814 150134 58000 6 vccd2
port 508 nsew power input
rlabel metal4 s 185514 -3814 186134 58000 6 vccd2
port 508 nsew power input
rlabel metal4 s 221514 -3814 222134 58000 6 vccd2
port 508 nsew power input
rlabel metal4 s 257514 -3814 258134 58000 6 vccd2
port 508 nsew power input
rlabel metal4 s 293514 -3814 294134 58000 6 vccd2
port 508 nsew power input
rlabel metal4 s 329514 -3814 330134 58000 6 vccd2
port 508 nsew power input
rlabel metal4 s 365514 -3814 366134 58000 6 vccd2
port 508 nsew power input
rlabel metal4 s 401514 -3814 402134 58000 6 vccd2
port 508 nsew power input
rlabel metal4 s 437514 -3814 438134 58000 6 vccd2
port 508 nsew power input
rlabel metal4 s 473514 -3814 474134 58000 6 vccd2
port 508 nsew power input
rlabel metal4 s 509514 -3814 510134 58000 6 vccd2
port 508 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 508 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 508 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 77514 562004 78134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 113514 562004 114134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 149514 562004 150134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 185514 562004 186134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 221514 562004 222134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 257514 562004 258134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 293514 562004 294134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 329514 562004 330134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 365514 562004 366134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 401514 562004 402134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 437514 562004 438134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 473514 562004 474134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 509514 562004 510134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 508 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 509 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 82306 58000 82926 6 vdda1
port 509 nsew power input
rlabel metal5 s 541964 82306 590730 82926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 118306 58000 118926 6 vdda1
port 509 nsew power input
rlabel metal5 s 541964 118306 590730 118926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 154306 58000 154926 6 vdda1
port 509 nsew power input
rlabel metal5 s 541964 154306 590730 154926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 190306 58000 190926 6 vdda1
port 509 nsew power input
rlabel metal5 s 541964 190306 590730 190926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 226306 58000 226926 6 vdda1
port 509 nsew power input
rlabel metal5 s 541964 226306 590730 226926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 262306 58000 262926 6 vdda1
port 509 nsew power input
rlabel metal5 s 541964 262306 590730 262926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 298306 58000 298926 6 vdda1
port 509 nsew power input
rlabel metal5 s 541964 298306 590730 298926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 334306 58000 334926 6 vdda1
port 509 nsew power input
rlabel metal5 s 541964 334306 590730 334926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 370306 58000 370926 6 vdda1
port 509 nsew power input
rlabel metal5 s 541964 370306 590730 370926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 406306 58000 406926 6 vdda1
port 509 nsew power input
rlabel metal5 s 541964 406306 590730 406926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 442306 58000 442926 6 vdda1
port 509 nsew power input
rlabel metal5 s 541964 442306 590730 442926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 478306 58000 478926 6 vdda1
port 509 nsew power input
rlabel metal5 s 541964 478306 590730 478926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 514306 58000 514926 6 vdda1
port 509 nsew power input
rlabel metal5 s 541964 514306 590730 514926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 550306 58000 550926 6 vdda1
port 509 nsew power input
rlabel metal5 s 541964 550306 590730 550926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 509 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 509 nsew power input
rlabel metal4 s 81234 -5734 81854 58000 6 vdda1
port 509 nsew power input
rlabel metal4 s 117234 -5734 117854 58000 6 vdda1
port 509 nsew power input
rlabel metal4 s 153234 -5734 153854 58000 6 vdda1
port 509 nsew power input
rlabel metal4 s 189234 -5734 189854 58000 6 vdda1
port 509 nsew power input
rlabel metal4 s 225234 -5734 225854 58000 6 vdda1
port 509 nsew power input
rlabel metal4 s 261234 -5734 261854 58000 6 vdda1
port 509 nsew power input
rlabel metal4 s 297234 -5734 297854 58000 6 vdda1
port 509 nsew power input
rlabel metal4 s 333234 -5734 333854 58000 6 vdda1
port 509 nsew power input
rlabel metal4 s 369234 -5734 369854 58000 6 vdda1
port 509 nsew power input
rlabel metal4 s 405234 -5734 405854 58000 6 vdda1
port 509 nsew power input
rlabel metal4 s 441234 -5734 441854 58000 6 vdda1
port 509 nsew power input
rlabel metal4 s 477234 -5734 477854 58000 6 vdda1
port 509 nsew power input
rlabel metal4 s 513234 -5734 513854 58000 6 vdda1
port 509 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 509 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 509 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 81234 562004 81854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 117234 562004 117854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 153234 562004 153854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 189234 562004 189854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 225234 562004 225854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 261234 562004 261854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 297234 562004 297854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 333234 562004 333854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 369234 562004 369854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 405234 562004 405854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 441234 562004 441854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 477234 562004 477854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 513234 562004 513854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 509 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 510 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 86026 58000 86646 6 vdda2
port 510 nsew power input
rlabel metal5 s 541964 86026 592650 86646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 122026 58000 122646 6 vdda2
port 510 nsew power input
rlabel metal5 s 541964 122026 592650 122646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 158026 58000 158646 6 vdda2
port 510 nsew power input
rlabel metal5 s 541964 158026 592650 158646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 194026 58000 194646 6 vdda2
port 510 nsew power input
rlabel metal5 s 541964 194026 592650 194646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 230026 58000 230646 6 vdda2
port 510 nsew power input
rlabel metal5 s 541964 230026 592650 230646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 266026 58000 266646 6 vdda2
port 510 nsew power input
rlabel metal5 s 541964 266026 592650 266646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 302026 58000 302646 6 vdda2
port 510 nsew power input
rlabel metal5 s 541964 302026 592650 302646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 338026 58000 338646 6 vdda2
port 510 nsew power input
rlabel metal5 s 541964 338026 592650 338646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 374026 58000 374646 6 vdda2
port 510 nsew power input
rlabel metal5 s 541964 374026 592650 374646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 410026 58000 410646 6 vdda2
port 510 nsew power input
rlabel metal5 s 541964 410026 592650 410646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 446026 58000 446646 6 vdda2
port 510 nsew power input
rlabel metal5 s 541964 446026 592650 446646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 482026 58000 482646 6 vdda2
port 510 nsew power input
rlabel metal5 s 541964 482026 592650 482646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 518026 58000 518646 6 vdda2
port 510 nsew power input
rlabel metal5 s 541964 518026 592650 518646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 554026 58000 554646 6 vdda2
port 510 nsew power input
rlabel metal5 s 541964 554026 592650 554646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 510 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 510 nsew power input
rlabel metal4 s 84954 -7654 85574 58000 6 vdda2
port 510 nsew power input
rlabel metal4 s 120954 -7654 121574 58000 6 vdda2
port 510 nsew power input
rlabel metal4 s 156954 -7654 157574 58000 6 vdda2
port 510 nsew power input
rlabel metal4 s 192954 -7654 193574 58000 6 vdda2
port 510 nsew power input
rlabel metal4 s 228954 -7654 229574 58000 6 vdda2
port 510 nsew power input
rlabel metal4 s 264954 -7654 265574 58000 6 vdda2
port 510 nsew power input
rlabel metal4 s 300954 -7654 301574 58000 6 vdda2
port 510 nsew power input
rlabel metal4 s 336954 -7654 337574 58000 6 vdda2
port 510 nsew power input
rlabel metal4 s 372954 -7654 373574 58000 6 vdda2
port 510 nsew power input
rlabel metal4 s 408954 -7654 409574 58000 6 vdda2
port 510 nsew power input
rlabel metal4 s 444954 -7654 445574 58000 6 vdda2
port 510 nsew power input
rlabel metal4 s 480954 -7654 481574 58000 6 vdda2
port 510 nsew power input
rlabel metal4 s 516954 -7654 517574 58000 6 vdda2
port 510 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 510 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 510 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 84954 562004 85574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 120954 562004 121574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 156954 562004 157574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 192954 562004 193574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 228954 562004 229574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 264954 562004 265574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 300954 562004 301574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 336954 562004 337574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 372954 562004 373574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 408954 562004 409574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 444954 562004 445574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 480954 562004 481574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 516954 562004 517574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 510 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 64306 58000 64926 6 vssa1
port 511 nsew ground input
rlabel metal5 s 541964 64306 590730 64926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 100306 58000 100926 6 vssa1
port 511 nsew ground input
rlabel metal5 s 541964 100306 590730 100926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 136306 58000 136926 6 vssa1
port 511 nsew ground input
rlabel metal5 s 541964 136306 590730 136926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 172306 58000 172926 6 vssa1
port 511 nsew ground input
rlabel metal5 s 541964 172306 590730 172926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 208306 58000 208926 6 vssa1
port 511 nsew ground input
rlabel metal5 s 541964 208306 590730 208926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 244306 58000 244926 6 vssa1
port 511 nsew ground input
rlabel metal5 s 541964 244306 590730 244926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 280306 58000 280926 6 vssa1
port 511 nsew ground input
rlabel metal5 s 541964 280306 590730 280926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 316306 58000 316926 6 vssa1
port 511 nsew ground input
rlabel metal5 s 541964 316306 590730 316926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 352306 58000 352926 6 vssa1
port 511 nsew ground input
rlabel metal5 s 541964 352306 590730 352926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 388306 58000 388926 6 vssa1
port 511 nsew ground input
rlabel metal5 s 541964 388306 590730 388926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 424306 58000 424926 6 vssa1
port 511 nsew ground input
rlabel metal5 s 541964 424306 590730 424926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 460306 58000 460926 6 vssa1
port 511 nsew ground input
rlabel metal5 s 541964 460306 590730 460926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 496306 58000 496926 6 vssa1
port 511 nsew ground input
rlabel metal5 s 541964 496306 590730 496926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 532306 58000 532926 6 vssa1
port 511 nsew ground input
rlabel metal5 s 541964 532306 590730 532926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 63234 -5734 63854 58000 6 vssa1
port 511 nsew ground input
rlabel metal4 s 99234 -5734 99854 58000 6 vssa1
port 511 nsew ground input
rlabel metal4 s 135234 -5734 135854 58000 6 vssa1
port 511 nsew ground input
rlabel metal4 s 171234 -5734 171854 58000 6 vssa1
port 511 nsew ground input
rlabel metal4 s 207234 -5734 207854 58000 6 vssa1
port 511 nsew ground input
rlabel metal4 s 243234 -5734 243854 58000 6 vssa1
port 511 nsew ground input
rlabel metal4 s 279234 -5734 279854 58000 6 vssa1
port 511 nsew ground input
rlabel metal4 s 315234 -5734 315854 58000 6 vssa1
port 511 nsew ground input
rlabel metal4 s 351234 -5734 351854 58000 6 vssa1
port 511 nsew ground input
rlabel metal4 s 387234 -5734 387854 58000 6 vssa1
port 511 nsew ground input
rlabel metal4 s 423234 -5734 423854 58000 6 vssa1
port 511 nsew ground input
rlabel metal4 s 459234 -5734 459854 58000 6 vssa1
port 511 nsew ground input
rlabel metal4 s 495234 -5734 495854 58000 6 vssa1
port 511 nsew ground input
rlabel metal4 s 531234 -5734 531854 58000 6 vssa1
port 511 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 511 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 63234 562004 63854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 99234 562004 99854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 135234 562004 135854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 171234 562004 171854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 207234 562004 207854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 243234 562004 243854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 279234 562004 279854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 315234 562004 315854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 351234 562004 351854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 387234 562004 387854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 423234 562004 423854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 459234 562004 459854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 495234 562004 495854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 531234 562004 531854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 511 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 68026 58000 68646 6 vssa2
port 512 nsew ground input
rlabel metal5 s 541964 68026 592650 68646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 104026 58000 104646 6 vssa2
port 512 nsew ground input
rlabel metal5 s 541964 104026 592650 104646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 140026 58000 140646 6 vssa2
port 512 nsew ground input
rlabel metal5 s 541964 140026 592650 140646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 176026 58000 176646 6 vssa2
port 512 nsew ground input
rlabel metal5 s 541964 176026 592650 176646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 212026 58000 212646 6 vssa2
port 512 nsew ground input
rlabel metal5 s 541964 212026 592650 212646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 248026 58000 248646 6 vssa2
port 512 nsew ground input
rlabel metal5 s 541964 248026 592650 248646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 284026 58000 284646 6 vssa2
port 512 nsew ground input
rlabel metal5 s 541964 284026 592650 284646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 320026 58000 320646 6 vssa2
port 512 nsew ground input
rlabel metal5 s 541964 320026 592650 320646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 356026 58000 356646 6 vssa2
port 512 nsew ground input
rlabel metal5 s 541964 356026 592650 356646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 392026 58000 392646 6 vssa2
port 512 nsew ground input
rlabel metal5 s 541964 392026 592650 392646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 428026 58000 428646 6 vssa2
port 512 nsew ground input
rlabel metal5 s 541964 428026 592650 428646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 464026 58000 464646 6 vssa2
port 512 nsew ground input
rlabel metal5 s 541964 464026 592650 464646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 500026 58000 500646 6 vssa2
port 512 nsew ground input
rlabel metal5 s 541964 500026 592650 500646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 536026 58000 536646 6 vssa2
port 512 nsew ground input
rlabel metal5 s 541964 536026 592650 536646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 66954 -7654 67574 58000 6 vssa2
port 512 nsew ground input
rlabel metal4 s 102954 -7654 103574 58000 6 vssa2
port 512 nsew ground input
rlabel metal4 s 138954 -7654 139574 58000 6 vssa2
port 512 nsew ground input
rlabel metal4 s 174954 -7654 175574 58000 6 vssa2
port 512 nsew ground input
rlabel metal4 s 210954 -7654 211574 58000 6 vssa2
port 512 nsew ground input
rlabel metal4 s 246954 -7654 247574 58000 6 vssa2
port 512 nsew ground input
rlabel metal4 s 282954 -7654 283574 58000 6 vssa2
port 512 nsew ground input
rlabel metal4 s 318954 -7654 319574 58000 6 vssa2
port 512 nsew ground input
rlabel metal4 s 354954 -7654 355574 58000 6 vssa2
port 512 nsew ground input
rlabel metal4 s 390954 -7654 391574 58000 6 vssa2
port 512 nsew ground input
rlabel metal4 s 426954 -7654 427574 58000 6 vssa2
port 512 nsew ground input
rlabel metal4 s 462954 -7654 463574 58000 6 vssa2
port 512 nsew ground input
rlabel metal4 s 498954 -7654 499574 58000 6 vssa2
port 512 nsew ground input
rlabel metal4 s 534954 -7654 535574 58000 6 vssa2
port 512 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 512 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 66954 562004 67574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 102954 562004 103574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 138954 562004 139574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 174954 562004 175574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 210954 562004 211574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 246954 562004 247574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 282954 562004 283574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 318954 562004 319574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 354954 562004 355574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 390954 562004 391574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 426954 562004 427574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 462954 562004 463574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 498954 562004 499574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 534954 562004 535574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 512 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 92866 58000 93486 6 vssd1
port 513 nsew ground input
rlabel metal5 s 541964 92866 586890 93486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 128866 58000 129486 6 vssd1
port 513 nsew ground input
rlabel metal5 s 541964 128866 586890 129486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 164866 58000 165486 6 vssd1
port 513 nsew ground input
rlabel metal5 s 541964 164866 586890 165486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 200866 58000 201486 6 vssd1
port 513 nsew ground input
rlabel metal5 s 541964 200866 586890 201486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 236866 58000 237486 6 vssd1
port 513 nsew ground input
rlabel metal5 s 541964 236866 586890 237486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 272866 58000 273486 6 vssd1
port 513 nsew ground input
rlabel metal5 s 541964 272866 586890 273486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 308866 58000 309486 6 vssd1
port 513 nsew ground input
rlabel metal5 s 541964 308866 586890 309486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 344866 58000 345486 6 vssd1
port 513 nsew ground input
rlabel metal5 s 541964 344866 586890 345486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 380866 58000 381486 6 vssd1
port 513 nsew ground input
rlabel metal5 s 541964 380866 586890 381486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 416866 58000 417486 6 vssd1
port 513 nsew ground input
rlabel metal5 s 541964 416866 586890 417486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 452866 58000 453486 6 vssd1
port 513 nsew ground input
rlabel metal5 s 541964 452866 586890 453486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 488866 58000 489486 6 vssd1
port 513 nsew ground input
rlabel metal5 s 541964 488866 586890 489486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 524866 58000 525486 6 vssd1
port 513 nsew ground input
rlabel metal5 s 541964 524866 586890 525486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 560866 58000 561486 6 vssd1
port 513 nsew ground input
rlabel metal5 s 541964 560866 586890 561486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 91794 -1894 92414 58000 6 vssd1
port 513 nsew ground input
rlabel metal4 s 127794 -1894 128414 58000 6 vssd1
port 513 nsew ground input
rlabel metal4 s 163794 -1894 164414 58000 6 vssd1
port 513 nsew ground input
rlabel metal4 s 199794 -1894 200414 58000 6 vssd1
port 513 nsew ground input
rlabel metal4 s 235794 -1894 236414 58000 6 vssd1
port 513 nsew ground input
rlabel metal4 s 271794 -1894 272414 58000 6 vssd1
port 513 nsew ground input
rlabel metal4 s 307794 -1894 308414 58000 6 vssd1
port 513 nsew ground input
rlabel metal4 s 343794 -1894 344414 58000 6 vssd1
port 513 nsew ground input
rlabel metal4 s 379794 -1894 380414 58000 6 vssd1
port 513 nsew ground input
rlabel metal4 s 415794 -1894 416414 58000 6 vssd1
port 513 nsew ground input
rlabel metal4 s 451794 -1894 452414 58000 6 vssd1
port 513 nsew ground input
rlabel metal4 s 487794 -1894 488414 58000 6 vssd1
port 513 nsew ground input
rlabel metal4 s 523794 -1894 524414 58000 6 vssd1
port 513 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 513 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 91794 562004 92414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 127794 562004 128414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 163794 562004 164414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 199794 562004 200414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 235794 562004 236414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 271794 562004 272414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 307794 562004 308414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 343794 562004 344414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 379794 562004 380414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 415794 562004 416414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 451794 562004 452414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 487794 562004 488414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 523794 562004 524414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 513 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 60586 58000 61206 6 vssd2
port 514 nsew ground input
rlabel metal5 s 541964 60586 588810 61206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 96586 58000 97206 6 vssd2
port 514 nsew ground input
rlabel metal5 s 541964 96586 588810 97206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 132586 58000 133206 6 vssd2
port 514 nsew ground input
rlabel metal5 s 541964 132586 588810 133206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 168586 58000 169206 6 vssd2
port 514 nsew ground input
rlabel metal5 s 541964 168586 588810 169206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 204586 58000 205206 6 vssd2
port 514 nsew ground input
rlabel metal5 s 541964 204586 588810 205206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 240586 58000 241206 6 vssd2
port 514 nsew ground input
rlabel metal5 s 541964 240586 588810 241206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 276586 58000 277206 6 vssd2
port 514 nsew ground input
rlabel metal5 s 541964 276586 588810 277206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 312586 58000 313206 6 vssd2
port 514 nsew ground input
rlabel metal5 s 541964 312586 588810 313206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 348586 58000 349206 6 vssd2
port 514 nsew ground input
rlabel metal5 s 541964 348586 588810 349206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 384586 58000 385206 6 vssd2
port 514 nsew ground input
rlabel metal5 s 541964 384586 588810 385206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 420586 58000 421206 6 vssd2
port 514 nsew ground input
rlabel metal5 s 541964 420586 588810 421206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 456586 58000 457206 6 vssd2
port 514 nsew ground input
rlabel metal5 s 541964 456586 588810 457206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 492586 58000 493206 6 vssd2
port 514 nsew ground input
rlabel metal5 s 541964 492586 588810 493206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 528586 58000 529206 6 vssd2
port 514 nsew ground input
rlabel metal5 s 541964 528586 588810 529206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 59514 -3814 60134 58000 6 vssd2
port 514 nsew ground input
rlabel metal4 s 95514 -3814 96134 58000 6 vssd2
port 514 nsew ground input
rlabel metal4 s 131514 -3814 132134 58000 6 vssd2
port 514 nsew ground input
rlabel metal4 s 167514 -3814 168134 58000 6 vssd2
port 514 nsew ground input
rlabel metal4 s 203514 -3814 204134 58000 6 vssd2
port 514 nsew ground input
rlabel metal4 s 239514 -3814 240134 58000 6 vssd2
port 514 nsew ground input
rlabel metal4 s 275514 -3814 276134 58000 6 vssd2
port 514 nsew ground input
rlabel metal4 s 311514 -3814 312134 58000 6 vssd2
port 514 nsew ground input
rlabel metal4 s 347514 -3814 348134 58000 6 vssd2
port 514 nsew ground input
rlabel metal4 s 383514 -3814 384134 58000 6 vssd2
port 514 nsew ground input
rlabel metal4 s 419514 -3814 420134 58000 6 vssd2
port 514 nsew ground input
rlabel metal4 s 455514 -3814 456134 58000 6 vssd2
port 514 nsew ground input
rlabel metal4 s 491514 -3814 492134 58000 6 vssd2
port 514 nsew ground input
rlabel metal4 s 527514 -3814 528134 58000 6 vssd2
port 514 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 514 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 59514 562004 60134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 95514 562004 96134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 131514 562004 132134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 167514 562004 168134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 203514 562004 204134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 239514 562004 240134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 275514 562004 276134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 311514 562004 312134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 347514 562004 348134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 383514 562004 384134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 419514 562004 420134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 455514 562004 456134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 491514 562004 492134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 527514 562004 528134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 514 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 515 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 516 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 517 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 518 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 519 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 520 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 521 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 522 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 523 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 524 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 525 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 526 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 527 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 528 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 529 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 530 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 531 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 532 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 533 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 534 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 535 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 536 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 537 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 538 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 539 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 540 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 541 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 542 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 543 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 544 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 545 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 546 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 547 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 548 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 549 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 550 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 551 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 552 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 553 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 554 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 555 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 556 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 557 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 558 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 559 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 560 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 561 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 562 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 563 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 564 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 565 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 566 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 567 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 568 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 569 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 570 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 571 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 572 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 573 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 574 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 575 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 576 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 577 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 578 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 579 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 580 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 581 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 582 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 583 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 584 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 585 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 586 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 587 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 588 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 589 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 590 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 591 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 592 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 593 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 594 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 595 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 596 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 597 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 598 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 599 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 600 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 601 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 602 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 603 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 604 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 605 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 606 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 607 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 608 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 609 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 610 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 611 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 612 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 613 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 614 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 615 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 616 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 617 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 618 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 619 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 620 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
