##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Wed Jun  1 19:12:32 2022
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO azadi_soc_top_caravel
  CLASS BLOCK ;
  SIZE 2050.220000 BY 1949.900000 ;
  FOREIGN azadi_soc_top_caravel 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5386 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.0858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 48.928 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 4.010000 0.000000 4.310000 0.800000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 95.4106 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 4.72354 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 22.7465 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.132727 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1946.630000 0.800000 1946.930000 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 432.280000 0.000000 432.580000 0.800000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 145.380000 0.000000 145.680000 0.800000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.440000 0.000000 436.740000 0.800000 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 428.125000 0.000000 428.425000 0.800000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 423.965000 0.000000 424.265000 0.800000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 419.810000 0.000000 420.110000 0.800000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 415.650000 0.000000 415.950000 0.800000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 278.435000 0.000000 278.735000 0.800000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 274.280000 0.000000 274.580000 0.800000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.120000 0.000000 270.420000 0.800000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 265.960000 0.000000 266.260000 0.800000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 261.805000 0.000000 262.105000 0.800000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 257.645000 0.000000 257.945000 0.800000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 253.490000 0.000000 253.790000 0.800000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 249.330000 0.000000 249.630000 0.800000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 245.170000 0.000000 245.470000 0.800000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 241.015000 0.000000 241.315000 0.800000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.855000 0.000000 237.155000 0.800000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 232.700000 0.000000 233.000000 0.800000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 228.540000 0.000000 228.840000 0.800000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 224.380000 0.000000 224.680000 0.800000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 220.225000 0.000000 220.525000 0.800000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.065000 0.000000 216.365000 0.800000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 211.910000 0.000000 212.210000 0.800000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 207.750000 0.000000 208.050000 0.800000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 203.590000 0.000000 203.890000 0.800000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 199.435000 0.000000 199.735000 0.800000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 195.275000 0.000000 195.575000 0.800000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 191.120000 0.000000 191.420000 0.800000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 186.960000 0.000000 187.260000 0.800000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 182.800000 0.000000 183.100000 0.800000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.645000 0.000000 178.945000 0.800000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 174.485000 0.000000 174.785000 0.800000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 170.330000 0.000000 170.630000 0.800000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.170000 0.000000 166.470000 0.800000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 162.010000 0.000000 162.310000 0.800000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 157.855000 0.000000 158.155000 0.800000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 153.695000 0.000000 153.995000 0.800000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.540000 0.000000 149.840000 0.800000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 141.220000 0.000000 141.520000 0.800000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 137.065000 0.000000 137.365000 0.800000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 132.905000 0.000000 133.205000 0.800000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 128.750000 0.000000 129.050000 0.800000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 124.590000 0.000000 124.890000 0.800000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 120.430000 0.000000 120.730000 0.800000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.275000 0.000000 116.575000 0.800000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 112.115000 0.000000 112.415000 0.800000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 107.960000 0.000000 108.260000 0.800000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.800000 0.000000 104.100000 0.800000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 99.640000 0.000000 99.940000 0.800000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 95.485000 0.000000 95.785000 0.800000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.325000 0.000000 91.625000 0.800000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 87.170000 0.000000 87.470000 0.800000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.010000 0.000000 83.310000 0.800000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 78.850000 0.000000 79.150000 0.800000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.695000 0.000000 74.995000 0.800000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.535000 0.000000 70.835000 0.800000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 66.380000 0.000000 66.680000 0.800000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 62.220000 0.000000 62.520000 0.800000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 58.060000 0.000000 58.360000 0.800000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 53.905000 0.000000 54.205000 0.800000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 49.745000 0.000000 50.045000 0.800000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 45.590000 0.000000 45.890000 0.800000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 41.430000 0.000000 41.730000 0.800000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 37.270000 0.000000 37.570000 0.800000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 33.115000 0.000000 33.415000 0.800000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.955000 0.000000 29.255000 0.800000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 24.800000 0.000000 25.100000 0.800000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 20.640000 0.000000 20.940000 0.800000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 16.480000 0.000000 16.780000 0.800000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 12.325000 0.000000 12.625000 0.800000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 119.827 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 641.448 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 8.165000 0.000000 8.465000 0.800000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.95 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 411.490000 0.000000 411.790000 0.800000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.95 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 407.335000 0.000000 407.635000 0.800000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.95 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 403.175000 0.000000 403.475000 0.800000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.95 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 399.020000 0.000000 399.320000 0.800000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.95 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 394.860000 0.000000 395.160000 0.800000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.95 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 390.700000 0.000000 391.000000 0.800000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.95 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 386.545000 0.000000 386.845000 0.800000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.95 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 382.385000 0.000000 382.685000 0.800000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.95 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 378.230000 0.000000 378.530000 0.800000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.739 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.424 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.602 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3015.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 374.070000 0.000000 374.370000 0.800000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 119.872 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 641.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 369.910000 0.000000 370.210000 0.800000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 119.872 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 641.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 365.755000 0.000000 366.055000 0.800000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 119.872 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 641.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 361.595000 0.000000 361.895000 0.800000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 119.872 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 641.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 357.440000 0.000000 357.740000 0.800000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 119.872 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 641.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 353.280000 0.000000 353.580000 0.800000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 119.872 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 641.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 349.120000 0.000000 349.420000 0.800000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 119.872 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 641.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 344.965000 0.000000 345.265000 0.800000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 119.872 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 641.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 340.805000 0.000000 341.105000 0.800000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 119.872 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 641.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 336.650000 0.000000 336.950000 0.800000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 119.872 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 641.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 332.490000 0.000000 332.790000 0.800000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 119.872 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 641.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 328.330000 0.000000 328.630000 0.800000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 119.872 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 641.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 324.175000 0.000000 324.475000 0.800000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 119.872 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 641.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 320.015000 0.000000 320.315000 0.800000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 119.872 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 641.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 315.860000 0.000000 316.160000 0.800000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 119.872 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 641.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 311.700000 0.000000 312.000000 0.800000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 119.872 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 641.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 307.540000 0.000000 307.840000 0.800000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 119.872 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 641.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 303.385000 0.000000 303.685000 0.800000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 119.872 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 641.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 299.225000 0.000000 299.525000 0.800000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 119.872 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 641.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 295.070000 0.000000 295.370000 0.800000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 119.872 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 641.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 290.910000 0.000000 291.210000 0.800000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 119.872 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 641.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 286.750000 0.000000 287.050000 0.800000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 119.872 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 641.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 282.595000 0.000000 282.895000 0.800000 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 968.665000 0.000000 968.965000 0.800000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 964.505000 0.000000 964.805000 0.800000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 960.350000 0.000000 960.650000 0.800000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 956.190000 0.000000 956.490000 0.800000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 952.030000 0.000000 952.330000 0.800000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 947.875000 0.000000 948.175000 0.800000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 943.715000 0.000000 944.015000 0.800000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 939.560000 0.000000 939.860000 0.800000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 935.400000 0.000000 935.700000 0.800000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 931.240000 0.000000 931.540000 0.800000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 927.085000 0.000000 927.385000 0.800000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 922.925000 0.000000 923.225000 0.800000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 918.770000 0.000000 919.070000 0.800000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 914.610000 0.000000 914.910000 0.800000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 910.450000 0.000000 910.750000 0.800000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 906.295000 0.000000 906.595000 0.800000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 902.135000 0.000000 902.435000 0.800000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 897.980000 0.000000 898.280000 0.800000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 893.820000 0.000000 894.120000 0.800000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 889.660000 0.000000 889.960000 0.800000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 885.505000 0.000000 885.805000 0.800000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 881.345000 0.000000 881.645000 0.800000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 877.190000 0.000000 877.490000 0.800000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 873.030000 0.000000 873.330000 0.800000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 868.870000 0.000000 869.170000 0.800000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 864.715000 0.000000 865.015000 0.800000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 860.555000 0.000000 860.855000 0.800000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 856.400000 0.000000 856.700000 0.800000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 852.240000 0.000000 852.540000 0.800000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 848.080000 0.000000 848.380000 0.800000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 843.925000 0.000000 844.225000 0.800000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 839.765000 0.000000 840.065000 0.800000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.610000 0.000000 835.910000 0.800000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 831.450000 0.000000 831.750000 0.800000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 827.290000 0.000000 827.590000 0.800000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 823.135000 0.000000 823.435000 0.800000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 818.975000 0.000000 819.275000 0.800000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 814.820000 0.000000 815.120000 0.800000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 810.660000 0.000000 810.960000 0.800000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 806.500000 0.000000 806.800000 0.800000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 802.345000 0.000000 802.645000 0.800000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 798.185000 0.000000 798.485000 0.800000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.030000 0.000000 794.330000 0.800000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 789.870000 0.000000 790.170000 0.800000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 785.710000 0.000000 786.010000 0.800000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 781.555000 0.000000 781.855000 0.800000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 777.395000 0.000000 777.695000 0.800000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 773.240000 0.000000 773.540000 0.800000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 769.080000 0.000000 769.380000 0.800000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 764.920000 0.000000 765.220000 0.800000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 760.765000 0.000000 761.065000 0.800000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 756.605000 0.000000 756.905000 0.800000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 752.450000 0.000000 752.750000 0.800000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 748.290000 0.000000 748.590000 0.800000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 744.130000 0.000000 744.430000 0.800000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 739.975000 0.000000 740.275000 0.800000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 735.815000 0.000000 736.115000 0.800000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 731.660000 0.000000 731.960000 0.800000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 727.500000 0.000000 727.800000 0.800000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 723.340000 0.000000 723.640000 0.800000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 719.185000 0.000000 719.485000 0.800000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 715.025000 0.000000 715.325000 0.800000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 710.870000 0.000000 711.170000 0.800000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 706.710000 0.000000 707.010000 0.800000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 702.550000 0.000000 702.850000 0.800000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 698.395000 0.000000 698.695000 0.800000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 694.235000 0.000000 694.535000 0.800000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 690.080000 0.000000 690.380000 0.800000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 685.920000 0.000000 686.220000 0.800000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 681.760000 0.000000 682.060000 0.800000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 677.605000 0.000000 677.905000 0.800000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 673.445000 0.000000 673.745000 0.800000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.290000 0.000000 669.590000 0.800000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 665.130000 0.000000 665.430000 0.800000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 660.970000 0.000000 661.270000 0.800000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 656.815000 0.000000 657.115000 0.800000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 652.655000 0.000000 652.955000 0.800000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 648.500000 0.000000 648.800000 0.800000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 644.340000 0.000000 644.640000 0.800000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 640.180000 0.000000 640.480000 0.800000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 636.025000 0.000000 636.325000 0.800000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 631.865000 0.000000 632.165000 0.800000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 627.710000 0.000000 628.010000 0.800000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 623.550000 0.000000 623.850000 0.800000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 619.390000 0.000000 619.690000 0.800000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 615.235000 0.000000 615.535000 0.800000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 611.075000 0.000000 611.375000 0.800000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 606.920000 0.000000 607.220000 0.800000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 602.760000 0.000000 603.060000 0.800000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 598.600000 0.000000 598.900000 0.800000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 594.445000 0.000000 594.745000 0.800000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 590.285000 0.000000 590.585000 0.800000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.130000 0.000000 586.430000 0.800000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 581.970000 0.000000 582.270000 0.800000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 577.810000 0.000000 578.110000 0.800000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 573.655000 0.000000 573.955000 0.800000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 569.495000 0.000000 569.795000 0.800000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 565.340000 0.000000 565.640000 0.800000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 561.180000 0.000000 561.480000 0.800000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.020000 0.000000 557.320000 0.800000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 552.865000 0.000000 553.165000 0.800000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 548.705000 0.000000 549.005000 0.800000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 544.550000 0.000000 544.850000 0.800000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 540.390000 0.000000 540.690000 0.800000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 536.230000 0.000000 536.530000 0.800000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 532.075000 0.000000 532.375000 0.800000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 527.915000 0.000000 528.215000 0.800000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 523.760000 0.000000 524.060000 0.800000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 519.600000 0.000000 519.900000 0.800000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 515.440000 0.000000 515.740000 0.800000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 511.285000 0.000000 511.585000 0.800000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 507.125000 0.000000 507.425000 0.800000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 28.7841 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 154.456 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 502.970000 0.000000 503.270000 0.800000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 58.7733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 313.928 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 498.810000 0.000000 499.110000 0.800000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 88.1571 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 471.112 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 494.650000 0.000000 494.950000 0.800000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 55.5168 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 296.56 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 490.495000 0.000000 490.795000 0.800000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.9876 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 246.208 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 486.335000 0.000000 486.635000 0.800000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.5001 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.608 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 482.180000 0.000000 482.480000 0.800000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.0071 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.312 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 478.020000 0.000000 478.320000 0.800000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.8531 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 106.824 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 473.860000 0.000000 474.160000 0.800000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.6316 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 126.976 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 469.705000 0.000000 470.005000 0.800000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.1266 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 81.616 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 465.545000 0.000000 465.845000 0.800000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.6951 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 100.648 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 461.390000 0.000000 461.690000 0.800000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.9101 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 457.230000 0.000000 457.530000 0.800000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.5561 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 453.070000 0.000000 453.370000 0.800000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.0906 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 97.424 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 448.915000 0.000000 449.215000 0.800000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.5466 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 115.856 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 444.755000 0.000000 445.055000 0.800000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.0001 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123.608 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 440.600000 0.000000 440.900000 0.800000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.581 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.704 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.042 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2388.28 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1500.890000 0.000000 1501.190000 0.800000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1496.730000 0.000000 1497.030000 0.800000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1492.570000 0.000000 1492.870000 0.800000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 509.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2391.14 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1488.415000 0.000000 1488.715000 0.800000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 509.12 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2390.23 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1484.255000 0.000000 1484.555000 0.800000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1480.100000 0.000000 1480.400000 0.800000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1475.940000 0.000000 1476.240000 0.800000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1471.780000 0.000000 1472.080000 0.800000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1467.625000 0.000000 1467.925000 0.800000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1463.465000 0.000000 1463.765000 0.800000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1459.310000 0.000000 1459.610000 0.800000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1455.150000 0.000000 1455.450000 0.800000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1450.990000 0.000000 1451.290000 0.800000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 509.12 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2390.23 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1446.835000 0.000000 1447.135000 0.800000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 509.12 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2390.23 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1442.675000 0.000000 1442.975000 0.800000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1438.520000 0.000000 1438.820000 0.800000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1434.360000 0.000000 1434.660000 0.800000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1430.200000 0.000000 1430.500000 0.800000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1426.045000 0.000000 1426.345000 0.800000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1421.885000 0.000000 1422.185000 0.800000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1417.730000 0.000000 1418.030000 0.800000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1413.570000 0.000000 1413.870000 0.800000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1409.410000 0.000000 1409.710000 0.800000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1405.255000 0.000000 1405.555000 0.800000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1401.095000 0.000000 1401.395000 0.800000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1396.940000 0.000000 1397.240000 0.800000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1392.780000 0.000000 1393.080000 0.800000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1388.620000 0.000000 1388.920000 0.800000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1384.465000 0.000000 1384.765000 0.800000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1380.305000 0.000000 1380.605000 0.800000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1376.150000 0.000000 1376.450000 0.800000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1371.990000 0.000000 1372.290000 0.800000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1367.830000 0.000000 1368.130000 0.800000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 509.12 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2390.23 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1363.675000 0.000000 1363.975000 0.800000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 509.12 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2390.23 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1359.515000 0.000000 1359.815000 0.800000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1355.360000 0.000000 1355.660000 0.800000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1351.200000 0.000000 1351.500000 0.800000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1347.040000 0.000000 1347.340000 0.800000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1342.885000 0.000000 1343.185000 0.800000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1338.725000 0.000000 1339.025000 0.800000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1334.570000 0.000000 1334.870000 0.800000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 509.12 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2390.23 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1330.410000 0.000000 1330.710000 0.800000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 509.12 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2390.23 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1326.250000 0.000000 1326.550000 0.800000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1322.095000 0.000000 1322.395000 0.800000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1317.935000 0.000000 1318.235000 0.800000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1313.780000 0.000000 1314.080000 0.800000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1309.620000 0.000000 1309.920000 0.800000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1305.460000 0.000000 1305.760000 0.800000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1301.305000 0.000000 1301.605000 0.800000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1297.145000 0.000000 1297.445000 0.800000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1292.990000 0.000000 1293.290000 0.800000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1288.830000 0.000000 1289.130000 0.800000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1284.670000 0.000000 1284.970000 0.800000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.581 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.704 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.042 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2388.28 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1280.515000 0.000000 1280.815000 0.800000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 509.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2391.14 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1276.355000 0.000000 1276.655000 0.800000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 509.12 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2390.23 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1272.200000 0.000000 1272.500000 0.800000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 509.12 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2390.23 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1268.040000 0.000000 1268.340000 0.800000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 509.12 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2390.23 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1263.880000 0.000000 1264.180000 0.800000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 509.12 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2390.23 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1259.725000 0.000000 1260.025000 0.800000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 509.12 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2390.23 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1255.565000 0.000000 1255.865000 0.800000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 509.12 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2390.23 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1251.410000 0.000000 1251.710000 0.800000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 509.12 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2390.23 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1247.250000 0.000000 1247.550000 0.800000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 509.12 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2390.23 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1243.090000 0.000000 1243.390000 0.800000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 509.12 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2390.23 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1238.935000 0.000000 1239.235000 0.800000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.658 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 745.784 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.275 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3013.27 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1234.775000 0.000000 1235.075000 0.800000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 572.685 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3049.29 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1230.620000 0.000000 1230.920000 0.800000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1226.460000 0.000000 1226.760000 0.800000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1222.300000 0.000000 1222.600000 0.800000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1218.145000 0.000000 1218.445000 0.800000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1213.985000 0.000000 1214.285000 0.800000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1209.830000 0.000000 1210.130000 0.800000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1205.670000 0.000000 1205.970000 0.800000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.95 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1201.510000 0.000000 1201.810000 0.800000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.95 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1197.355000 0.000000 1197.655000 0.800000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1193.195000 0.000000 1193.495000 0.800000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1189.040000 0.000000 1189.340000 0.800000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1184.880000 0.000000 1185.180000 0.800000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1180.720000 0.000000 1181.020000 0.800000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1176.565000 0.000000 1176.865000 0.800000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1172.405000 0.000000 1172.705000 0.800000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1168.250000 0.000000 1168.550000 0.800000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1164.090000 0.000000 1164.390000 0.800000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1159.930000 0.000000 1160.230000 0.800000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1155.775000 0.000000 1156.075000 0.800000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1151.615000 0.000000 1151.915000 0.800000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1147.460000 0.000000 1147.760000 0.800000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1143.300000 0.000000 1143.600000 0.800000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1139.140000 0.000000 1139.440000 0.800000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1134.985000 0.000000 1135.285000 0.800000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1130.825000 0.000000 1131.125000 0.800000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1126.670000 0.000000 1126.970000 0.800000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1122.510000 0.000000 1122.810000 0.800000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.95 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1118.350000 0.000000 1118.650000 0.800000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.95 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1114.195000 0.000000 1114.495000 0.800000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1110.035000 0.000000 1110.335000 0.800000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1105.880000 0.000000 1106.180000 0.800000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1101.720000 0.000000 1102.020000 0.800000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1097.560000 0.000000 1097.860000 0.800000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1093.405000 0.000000 1093.705000 0.800000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1089.245000 0.000000 1089.545000 0.800000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1085.090000 0.000000 1085.390000 0.800000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1080.930000 0.000000 1081.230000 0.800000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1076.770000 0.000000 1077.070000 0.800000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.95 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1072.615000 0.000000 1072.915000 0.800000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.95 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1068.455000 0.000000 1068.755000 0.800000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1064.300000 0.000000 1064.600000 0.800000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1060.140000 0.000000 1060.440000 0.800000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1055.980000 0.000000 1056.280000 0.800000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1051.825000 0.000000 1052.125000 0.800000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1047.665000 0.000000 1047.965000 0.800000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1043.510000 0.000000 1043.810000 0.800000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1039.350000 0.000000 1039.650000 0.800000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.95 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1035.190000 0.000000 1035.490000 0.800000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.95 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1031.035000 0.000000 1031.335000 0.800000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1026.875000 0.000000 1027.175000 0.800000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1022.720000 0.000000 1023.020000 0.800000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1018.560000 0.000000 1018.860000 0.800000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1014.400000 0.000000 1014.700000 0.800000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1010.245000 0.000000 1010.545000 0.800000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1006.085000 0.000000 1006.385000 0.800000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1001.930000 0.000000 1002.230000 0.800000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 997.770000 0.000000 998.070000 0.800000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 993.610000 0.000000 993.910000 0.800000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 989.455000 0.000000 989.755000 0.800000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 985.295000 0.000000 985.595000 0.800000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 981.140000 0.000000 981.440000 0.800000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 976.980000 0.000000 977.280000 0.800000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 746.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 564.457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3014.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 972.820000 0.000000 973.120000 0.800000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2033.110000 0.000000 2033.410000 0.800000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2028.955000 0.000000 2029.255000 0.800000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2024.795000 0.000000 2025.095000 0.800000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2020.640000 0.000000 2020.940000 0.800000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2016.480000 0.000000 2016.780000 0.800000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2012.320000 0.000000 2012.620000 0.800000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2008.165000 0.000000 2008.465000 0.800000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2004.005000 0.000000 2004.305000 0.800000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1999.850000 0.000000 2000.150000 0.800000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1995.690000 0.000000 1995.990000 0.800000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1991.530000 0.000000 1991.830000 0.800000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1987.375000 0.000000 1987.675000 0.800000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1983.215000 0.000000 1983.515000 0.800000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1979.060000 0.000000 1979.360000 0.800000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1974.900000 0.000000 1975.200000 0.800000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1970.740000 0.000000 1971.040000 0.800000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1966.585000 0.000000 1966.885000 0.800000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1962.425000 0.000000 1962.725000 0.800000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1958.270000 0.000000 1958.570000 0.800000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1954.110000 0.000000 1954.410000 0.800000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1949.950000 0.000000 1950.250000 0.800000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1945.795000 0.000000 1946.095000 0.800000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1941.635000 0.000000 1941.935000 0.800000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1937.480000 0.000000 1937.780000 0.800000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1933.320000 0.000000 1933.620000 0.800000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1929.160000 0.000000 1929.460000 0.800000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1925.005000 0.000000 1925.305000 0.800000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1920.845000 0.000000 1921.145000 0.800000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1916.690000 0.000000 1916.990000 0.800000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1912.530000 0.000000 1912.830000 0.800000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1908.370000 0.000000 1908.670000 0.800000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1904.215000 0.000000 1904.515000 0.800000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1900.055000 0.000000 1900.355000 0.800000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1895.900000 0.000000 1896.200000 0.800000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1891.740000 0.000000 1892.040000 0.800000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1887.580000 0.000000 1887.880000 0.800000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1883.425000 0.000000 1883.725000 0.800000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1879.265000 0.000000 1879.565000 0.800000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1875.110000 0.000000 1875.410000 0.800000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1870.950000 0.000000 1871.250000 0.800000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1866.790000 0.000000 1867.090000 0.800000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1862.635000 0.000000 1862.935000 0.800000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1858.475000 0.000000 1858.775000 0.800000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1854.320000 0.000000 1854.620000 0.800000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1850.160000 0.000000 1850.460000 0.800000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1846.000000 0.000000 1846.300000 0.800000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1841.845000 0.000000 1842.145000 0.800000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1837.685000 0.000000 1837.985000 0.800000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1833.530000 0.000000 1833.830000 0.800000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1829.370000 0.000000 1829.670000 0.800000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1825.210000 0.000000 1825.510000 0.800000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1821.055000 0.000000 1821.355000 0.800000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1816.895000 0.000000 1817.195000 0.800000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1812.740000 0.000000 1813.040000 0.800000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1808.580000 0.000000 1808.880000 0.800000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1804.420000 0.000000 1804.720000 0.800000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1800.265000 0.000000 1800.565000 0.800000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.105000 0.000000 1796.405000 0.800000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1791.950000 0.000000 1792.250000 0.800000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1787.790000 0.000000 1788.090000 0.800000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1783.630000 0.000000 1783.930000 0.800000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1779.475000 0.000000 1779.775000 0.800000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1775.315000 0.000000 1775.615000 0.800000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1771.160000 0.000000 1771.460000 0.800000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1767.000000 0.000000 1767.300000 0.800000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1762.840000 0.000000 1763.140000 0.800000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1758.685000 0.000000 1758.985000 0.800000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1754.525000 0.000000 1754.825000 0.800000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1750.370000 0.000000 1750.670000 0.800000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1746.210000 0.000000 1746.510000 0.800000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1742.050000 0.000000 1742.350000 0.800000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1737.895000 0.000000 1738.195000 0.800000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1733.735000 0.000000 1734.035000 0.800000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1729.580000 0.000000 1729.880000 0.800000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1725.420000 0.000000 1725.720000 0.800000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1721.260000 0.000000 1721.560000 0.800000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1717.105000 0.000000 1717.405000 0.800000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1712.945000 0.000000 1713.245000 0.800000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1708.790000 0.000000 1709.090000 0.800000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1704.630000 0.000000 1704.930000 0.800000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1700.470000 0.000000 1700.770000 0.800000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.315000 0.000000 1696.615000 0.800000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1692.155000 0.000000 1692.455000 0.800000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1688.000000 0.000000 1688.300000 0.800000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1683.840000 0.000000 1684.140000 0.800000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1679.680000 0.000000 1679.980000 0.800000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1675.525000 0.000000 1675.825000 0.800000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1671.365000 0.000000 1671.665000 0.800000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1667.210000 0.000000 1667.510000 0.800000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1663.050000 0.000000 1663.350000 0.800000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1658.890000 0.000000 1659.190000 0.800000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1654.735000 0.000000 1655.035000 0.800000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1650.575000 0.000000 1650.875000 0.800000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1646.420000 0.000000 1646.720000 0.800000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1642.260000 0.000000 1642.560000 0.800000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1638.100000 0.000000 1638.400000 0.800000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1633.945000 0.000000 1634.245000 0.800000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1629.785000 0.000000 1630.085000 0.800000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1625.630000 0.000000 1625.930000 0.800000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1621.470000 0.000000 1621.770000 0.800000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1617.310000 0.000000 1617.610000 0.800000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1613.155000 0.000000 1613.455000 0.800000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1608.995000 0.000000 1609.295000 0.800000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1604.840000 0.000000 1605.140000 0.800000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1600.680000 0.000000 1600.980000 0.800000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.520000 0.000000 1596.820000 0.800000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1592.365000 0.000000 1592.665000 0.800000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1588.205000 0.000000 1588.505000 0.800000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1584.050000 0.000000 1584.350000 0.800000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1579.890000 0.000000 1580.190000 0.800000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1575.730000 0.000000 1576.030000 0.800000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1571.575000 0.000000 1571.875000 0.800000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1567.415000 0.000000 1567.715000 0.800000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1563.260000 0.000000 1563.560000 0.800000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1559.100000 0.000000 1559.400000 0.800000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1554.940000 0.000000 1555.240000 0.800000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1550.785000 0.000000 1551.085000 0.800000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1546.625000 0.000000 1546.925000 0.800000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1542.470000 0.000000 1542.770000 0.800000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1538.310000 0.000000 1538.610000 0.800000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1534.150000 0.000000 1534.450000 0.800000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1529.995000 0.000000 1530.295000 0.800000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1525.835000 0.000000 1526.135000 0.800000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1521.680000 0.000000 1521.980000 0.800000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1517.520000 0.000000 1517.820000 0.800000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1513.360000 0.000000 1513.660000 0.800000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1509.205000 0.000000 1509.505000 0.800000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1505.045000 0.000000 1505.345000 0.800000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 882.810000 0.800000 883.110000 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5063 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 846.020000 0.800000 846.320000 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.3124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 146.128 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 144.992 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 773.76 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 809.230000 0.800000 809.530000 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 46.1524 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 246.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 121.154 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 646.624 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 772.440000 0.800000 772.740000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.784 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 735.650000 0.800000 735.950000 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 698.860000 0.800000 699.160000 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 662.070000 0.800000 662.370000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 625.280000 0.800000 625.580000 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.9814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 93.9243 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 501.4 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 588.490000 0.800000 588.790000 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2386 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 118.61 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 633.056 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 551.700000 0.800000 552.000000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.4584 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.24 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.8943 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 101.24 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 514.910000 0.800000 515.210000 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5916 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 115.409 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 615.984 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 478.120000 0.800000 478.420000 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8044 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.0773 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 102.216 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 441.330000 0.800000 441.630000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.2111 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 103.4 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 404.540000 0.800000 404.840000 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2701 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.7758 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.608 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 117.005000 1949.100000 117.305000 1949.900000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3973 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.256 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 351.310000 1949.100000 351.610000 1949.900000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 86.7099 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 463.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 585.620000 1949.100000 585.920000 1949.900000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.8883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 192.248 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 819.930000 1949.100000 820.230000 1949.900000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 42.2646 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 226.352 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1054.235000 1949.100000 1054.535000 1949.900000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 49.9254 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 267.68 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1288.545000 1949.100000 1288.845000 1949.900000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 47.5389 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 254.952 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1522.850000 1949.100000 1523.150000 1949.900000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 28.2921 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 151.832 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1757.160000 1949.100000 1757.460000 1949.900000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1991.470000 1949.100000 1991.770000 1949.900000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 1087.290000 2050.220000 1087.590000 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8806 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 63.6438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 339.904 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 1124.790000 2050.220000 1125.090000 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1174 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.088 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 67.0968 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 358.32 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 1162.290000 2050.220000 1162.590000 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1508 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.608 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 1199.785000 2050.220000 1200.085000 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4738 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 73.3188 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 391.504 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 1237.285000 2050.220000 1237.585000 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 1274.780000 2050.220000 1275.080000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 1312.280000 2050.220000 1312.580000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 28.3521 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 152.152 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 1349.780000 2050.220000 1350.080000 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 1387.275000 2050.220000 1387.575000 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.7798 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.296 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 1424.775000 2050.220000 1425.075000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 1462.270000 2050.220000 1462.570000 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 1499.770000 2050.220000 1500.070000 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.9933 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 1537.270000 2050.220000 1537.570000 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 1574.765000 2050.220000 1575.065000 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 1612.265000 2050.220000 1612.565000 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 119.902 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 641.848 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1912.930000 0.800000 1913.230000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5573 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.776 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1876.140000 0.800000 1876.440000 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3383 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.608 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1839.350000 0.800000 1839.650000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.0873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.936 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1802.560000 0.800000 1802.860000 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2386 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 52.9608 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 282.928 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1765.770000 0.800000 1766.070000 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 81.9198 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 437.376 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1728.980000 0.800000 1729.280000 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.3684 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.76 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 30.9363 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 165.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1692.190000 0.800000 1692.490000 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9083 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.648 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1655.400000 0.800000 1655.700000 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2553 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.832 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1618.610000 0.800000 1618.910000 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2386 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.641 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1075.89 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1581.820000 0.800000 1582.120000 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.912 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1545.030000 0.800000 1545.330000 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.912 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1508.240000 0.800000 1508.540000 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4836 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 197.576 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1054.21 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1471.450000 0.800000 1471.750000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.0901 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 108.088 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1434.660000 0.800000 1434.960000 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 50.2266 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 268.816 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 58.425000 1949.100000 58.725000 1949.900000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.6046 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 94.832 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 292.735000 1949.100000 293.035000 1949.900000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 85.2172 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 455.88 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 527.045000 1949.100000 527.345000 1949.900000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3853 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.192 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 761.350000 1949.100000 761.650000 1949.900000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 92.6619 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 495.608 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 995.660000 1949.100000 995.960000 1949.900000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 38.7888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 207.344 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1229.965000 1949.100000 1230.265000 1949.900000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 42.5946 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 228.112 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1464.275000 1949.100000 1464.575000 1949.900000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2131 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.128 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9348 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.456 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1698.585000 1949.100000 1698.885000 1949.900000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 38.4394 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 205.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.9748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.336 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1932.890000 1949.100000 1933.190000 1949.900000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6463 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.584 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 9.880000 2050.220000 10.180000 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.656 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 509.104 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.394 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2390.16 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 37.350000 2050.220000 37.650000 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.656 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 509.104 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.394 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2390.16 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 74.845000 2050.220000 75.145000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.656 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 509.104 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.394 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2390.16 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 112.345000 2050.220000 112.645000 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.656 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 509.104 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.394 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2390.16 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 149.840000 2050.220000 150.140000 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.9093 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.32 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 187.340000 2050.220000 187.640000 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.3713 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.784 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 224.840000 2050.220000 225.140000 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.656 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 509.104 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 453.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2433.17 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 262.335000 2050.220000 262.635000 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8038 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.424 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 299.835000 2050.220000 300.135000 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.656 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 509.104 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.394 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2390.16 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 337.330000 2050.220000 337.630000 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1253 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.472 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 374.830000 2050.220000 375.130000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.6538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 142.624 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 412.330000 2050.220000 412.630000 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.656 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 509.104 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.394 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2390.16 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 449.825000 2050.220000 450.125000 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.928 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 487.325000 2050.220000 487.625000 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0273 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 275.351 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1469.01 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 524.820000 2050.220000 525.120000 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 119.827 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 641.448 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1.460000 0.000000 1.760000 0.800000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.56 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1397.870000 0.800000 1398.170000 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6354 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1361.080000 0.800000 1361.380000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5094 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.192 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1324.290000 0.800000 1324.590000 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5664 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.496 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1287.500000 0.800000 1287.800000 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 119.902 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 641.848 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1250.710000 0.800000 1251.010000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 119.902 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 641.848 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1213.920000 0.800000 1214.220000 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 119.902 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 641.848 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1177.130000 0.800000 1177.430000 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4914 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.616 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1140.340000 0.800000 1140.640000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4694 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.832 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1103.550000 0.800000 1103.850000 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.8814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.696 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1066.760000 0.800000 1067.060000 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6954 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1029.970000 0.800000 1030.270000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2034 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.08 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 993.180000 0.800000 993.480000 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.384 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 956.390000 0.800000 956.690000 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3174 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 919.600000 0.800000 919.900000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 234.160000 1949.100000 234.460000 1949.900000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 84.7599 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 452.048 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 468.465000 1949.100000 468.765000 1949.900000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2079 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.104 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 702.775000 1949.100000 703.075000 1949.900000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 33.0054 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 176.024 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 937.080000 1949.100000 937.380000 1949.900000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3354 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.784 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1171.390000 1949.100000 1171.690000 1949.900000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 59.9154 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 319.544 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1405.700000 1949.100000 1406.000000 1949.900000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 66.2199 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 353.168 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1640.005000 1949.100000 1640.305000 1949.900000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 46.5619 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 248.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.3258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.208 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met4  ;
    ANTENNAMAXAREACAR 1.52958 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 10.3662 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1874.315000 1949.100000 1874.615000 1949.900000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.89645 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 55.4547 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 296.629 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.910329 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.3258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.208 LAYER met4  ;
    ANTENNAGATEAREA 0.213 LAYER met4  ;
    ANTENNAMAXAREACAR 56.9843 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 306.995 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.910329 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 1941.750000 2050.220000 1942.050000 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8903 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.408 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 562.320000 2050.220000 562.620000 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8903 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.408 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 599.820000 2050.220000 600.120000 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8903 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.408 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 637.315000 2050.220000 637.615000 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8903 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.408 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 674.815000 2050.220000 675.115000 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4344 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.312 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 712.310000 2050.220000 712.610000 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.344 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 749.810000 2050.220000 750.110000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8903 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.408 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 787.310000 2050.220000 787.610000 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.89645 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 27.6829 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 165.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.3258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.208 LAYER met4  ;
    ANTENNAGATEAREA 0.213 LAYER met4  ;
    ANTENNAMAXAREACAR 29.2124 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 175.662 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 824.805000 2050.220000 825.105000 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8903 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.408 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 862.305000 2050.220000 862.605000 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.89645 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 27.6829 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 165.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.3258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.208 LAYER met4  ;
    ANTENNAGATEAREA 0.213 LAYER met4  ;
    ANTENNAMAXAREACAR 29.2124 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 175.662 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 899.800000 2050.220000 900.100000 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.89645 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 27.6829 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 165.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.3258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.208 LAYER met4  ;
    ANTENNAGATEAREA 0.213 LAYER met4  ;
    ANTENNAMAXAREACAR 29.2124 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 175.662 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 937.300000 2050.220000 937.600000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8453 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 974.800000 2050.220000 975.100000 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.728 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 1012.295000 2050.220000 1012.595000 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.89645 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 27.6829 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 165.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.3258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.208 LAYER met4  ;
    ANTENNAGATEAREA 0.213 LAYER met4  ;
    ANTENNAMAXAREACAR 29.2124 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 175.662 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 1049.795000 2050.220000 1050.095000 ;
    END
  END io_oeb[0]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 367.750000 0.800000 368.050000 ;
    END
  END analog_io[28]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 330.960000 0.800000 331.260000 ;
    END
  END analog_io[27]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 294.170000 0.800000 294.470000 ;
    END
  END analog_io[26]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 257.380000 0.800000 257.680000 ;
    END
  END analog_io[25]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 220.590000 0.800000 220.890000 ;
    END
  END analog_io[24]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 183.800000 0.800000 184.100000 ;
    END
  END analog_io[23]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 147.010000 0.800000 147.310000 ;
    END
  END analog_io[22]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 110.220000 0.800000 110.520000 ;
    END
  END analog_io[21]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 73.430000 0.800000 73.730000 ;
    END
  END analog_io[20]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 36.640000 0.800000 36.940000 ;
    END
  END analog_io[19]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 7.440000 0.800000 7.740000 ;
    END
  END analog_io[18]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3.760000 1949.100000 4.060000 1949.900000 ;
    END
  END analog_io[17]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 175.580000 1949.100000 175.880000 1949.900000 ;
    END
  END analog_io[16]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 409.890000 1949.100000 410.190000 1949.900000 ;
    END
  END analog_io[15]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 644.195000 1949.100000 644.495000 1949.900000 ;
    END
  END analog_io[14]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 878.505000 1949.100000 878.805000 1949.900000 ;
    END
  END analog_io[13]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1112.815000 1949.100000 1113.115000 1949.900000 ;
    END
  END analog_io[12]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1347.120000 1949.100000 1347.420000 1949.900000 ;
    END
  END analog_io[11]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.430000 1949.100000 1581.730000 1949.900000 ;
    END
  END analog_io[10]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1815.735000 1949.100000 1816.035000 1949.900000 ;
    END
  END analog_io[9]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 1649.760000 2050.220000 1650.060000 ;
    END
  END analog_io[8]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 1687.260000 2050.220000 1687.560000 ;
    END
  END analog_io[7]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 1724.760000 2050.220000 1725.060000 ;
    END
  END analog_io[6]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 1762.255000 2050.220000 1762.555000 ;
    END
  END analog_io[5]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 1799.755000 2050.220000 1800.055000 ;
    END
  END analog_io[4]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 1837.250000 2050.220000 1837.550000 ;
    END
  END analog_io[3]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 1874.750000 2050.220000 1875.050000 ;
    END
  END analog_io[2]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2049.420000 1912.250000 2050.220000 1912.550000 ;
    END
  END analog_io[1]
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2035.580000 1949.100000 2035.880000 1949.900000 ;
    END
  END analog_io[0]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2037.270000 0.000000 2037.570000 0.800000 ;
    END
  END user_clock2
  PIN user_irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2389.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2045.585000 0.000000 2045.885000 0.800000 ;
    END
  END user_irq[2]
  PIN user_irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.581 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.704 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.042 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2388.28 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2048.000000 0.000000 2048.300000 0.800000 ;
    END
  END user_irq[1]
  PIN user_irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.581 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 508.704 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 444.042 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2388.28 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2041.430000 0.000000 2041.730000 0.800000 ;
    END
  END user_irq[0]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2029.750000 19.275000 2031.550000 1933.595000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2038.300000 2.660000 2040.100000 1945.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2045.500000 2.660000 2047.300000 1945.540000 ;
      LAYER met3 ;
        RECT 2045.500000 2.660000 2047.300000 1945.540000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.070000 19.275000 2031.550000 21.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.920000 2.660000 2047.300000 4.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.920000 1943.740000 2047.300000 1945.540000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.070000 1931.795000 2031.550000 1933.595000 ;
    END
    PORT
      LAYER met4 ;
        RECT 17.070000 19.275000 18.870000 1933.595000 ;
    END
    PORT
      LAYER met4 ;
        RECT 13.720000 2.660000 15.520000 1945.520000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.920000 2.660000 4.720000 1945.540000 ;
    END

# P/G pin shape extracted from block 'azadi_soc_top'
    PORT
      LAYER met4 ;
        RECT 71.250000 84.380000 72.990000 479.160000 ;
      LAYER met4 ;
        RECT 546.570000 84.380000 548.310000 479.160000 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.250000 1015.380000 72.990000 1410.160000 ;
      LAYER met4 ;
        RECT 546.570000 1015.380000 548.310000 1410.160000 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.250000 1480.880000 72.990000 1875.660000 ;
      LAYER met4 ;
        RECT 546.570000 1480.880000 548.310000 1875.660000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1498.130000 78.840000 1499.870000 473.620000 ;
      LAYER met4 ;
        RECT 1973.450000 78.840000 1975.190000 473.620000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1498.130000 544.340000 1499.870000 939.120000 ;
      LAYER met4 ;
        RECT 1973.450000 544.340000 1975.190000 939.120000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1498.130000 1009.840000 1499.870000 1404.620000 ;
      LAYER met4 ;
        RECT 1973.450000 1009.840000 1975.190000 1404.620000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1498.130000 1475.340000 1499.870000 1870.120000 ;
      LAYER met4 ;
        RECT 1973.450000 1475.340000 1975.190000 1870.120000 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.250000 549.880000 72.990000 944.660000 ;
      LAYER met4 ;
        RECT 546.570000 549.880000 548.310000 944.660000 ;
    END
    PORT
      LAYER met4 ;
        RECT 27.190000 29.135000 28.990000 1923.055000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2019.630000 29.135000 2021.430000 1923.055000 ;
    END
# end of P/G pin shape extracted from block 'azadi_soc_top'

  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2041.900000 6.260000 2043.700000 1941.940000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2034.700000 6.260000 2036.500000 1941.940000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2026.150000 22.875000 2027.950000 1929.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.520000 6.260000 2043.700000 8.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.670000 22.875000 2027.950000 24.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.670000 1928.195000 2027.950000 1929.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.520000 1940.140000 2043.700000 1941.940000 ;
    END
    PORT
      LAYER met4 ;
        RECT 20.670000 22.875000 22.470000 1929.995000 ;
    END
    PORT
      LAYER met4 ;
        RECT 10.120000 6.260000 11.920000 1941.940000 ;
    END
    PORT
      LAYER met4 ;
        RECT 6.520000 6.260000 8.320000 1941.940000 ;
    END

# P/G pin shape extracted from block 'azadi_soc_top'
    PORT
      LAYER met4 ;
        RECT 543.170000 87.780000 544.910000 475.760000 ;
      LAYER met4 ;
        RECT 74.650000 87.780000 76.390000 475.760000 ;
    END
    PORT
      LAYER met4 ;
        RECT 543.170000 1018.780000 544.910000 1406.760000 ;
      LAYER met4 ;
        RECT 74.650000 1018.780000 76.390000 1406.760000 ;
    END
    PORT
      LAYER met4 ;
        RECT 543.170000 1484.280000 544.910000 1872.260000 ;
      LAYER met4 ;
        RECT 74.650000 1484.280000 76.390000 1872.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1970.050000 82.240000 1971.790000 470.220000 ;
      LAYER met4 ;
        RECT 1501.530000 82.240000 1503.270000 470.220000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1970.050000 547.740000 1971.790000 935.720000 ;
      LAYER met4 ;
        RECT 1501.530000 547.740000 1503.270000 935.720000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1970.050000 1013.240000 1971.790000 1401.220000 ;
      LAYER met4 ;
        RECT 1501.530000 1013.240000 1503.270000 1401.220000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1970.050000 1478.740000 1971.790000 1866.720000 ;
      LAYER met4 ;
        RECT 1501.530000 1478.740000 1503.270000 1866.720000 ;
    END
    PORT
      LAYER met4 ;
        RECT 543.170000 553.280000 544.910000 941.260000 ;
      LAYER met4 ;
        RECT 74.650000 553.280000 76.390000 941.260000 ;
    END
    PORT
      LAYER met4 ;
        RECT 30.790000 32.735000 32.590000 1919.455000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2016.030000 32.735000 2017.830000 1919.455000 ;
    END
# end of P/G pin shape extracted from block 'azadi_soc_top'

  END vccd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 2050.220000 1949.900000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 2050.220000 1949.900000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 2050.220000 1949.900000 ;
    LAYER met3 ;
      RECT 2036.180000 1948.800000 2050.220000 1949.900000 ;
      RECT 1992.070000 1948.800000 2035.280000 1949.900000 ;
      RECT 1933.490000 1948.800000 1991.170000 1949.900000 ;
      RECT 1874.915000 1948.800000 1932.590000 1949.900000 ;
      RECT 1816.335000 1948.800000 1874.015000 1949.900000 ;
      RECT 1757.760000 1948.800000 1815.435000 1949.900000 ;
      RECT 1699.185000 1948.800000 1756.860000 1949.900000 ;
      RECT 1640.605000 1948.800000 1698.285000 1949.900000 ;
      RECT 1582.030000 1948.800000 1639.705000 1949.900000 ;
      RECT 1523.450000 1948.800000 1581.130000 1949.900000 ;
      RECT 1464.875000 1948.800000 1522.550000 1949.900000 ;
      RECT 1406.300000 1948.800000 1463.975000 1949.900000 ;
      RECT 1347.720000 1948.800000 1405.400000 1949.900000 ;
      RECT 1289.145000 1948.800000 1346.820000 1949.900000 ;
      RECT 1230.565000 1948.800000 1288.245000 1949.900000 ;
      RECT 1171.990000 1948.800000 1229.665000 1949.900000 ;
      RECT 1113.415000 1948.800000 1171.090000 1949.900000 ;
      RECT 1054.835000 1948.800000 1112.515000 1949.900000 ;
      RECT 996.260000 1948.800000 1053.935000 1949.900000 ;
      RECT 937.680000 1948.800000 995.360000 1949.900000 ;
      RECT 879.105000 1948.800000 936.780000 1949.900000 ;
      RECT 820.530000 1948.800000 878.205000 1949.900000 ;
      RECT 761.950000 1948.800000 819.630000 1949.900000 ;
      RECT 703.375000 1948.800000 761.050000 1949.900000 ;
      RECT 644.795000 1948.800000 702.475000 1949.900000 ;
      RECT 586.220000 1948.800000 643.895000 1949.900000 ;
      RECT 527.645000 1948.800000 585.320000 1949.900000 ;
      RECT 469.065000 1948.800000 526.745000 1949.900000 ;
      RECT 410.490000 1948.800000 468.165000 1949.900000 ;
      RECT 351.910000 1948.800000 409.590000 1949.900000 ;
      RECT 293.335000 1948.800000 351.010000 1949.900000 ;
      RECT 234.760000 1948.800000 292.435000 1949.900000 ;
      RECT 176.180000 1948.800000 233.860000 1949.900000 ;
      RECT 117.605000 1948.800000 175.280000 1949.900000 ;
      RECT 59.025000 1948.800000 116.705000 1949.900000 ;
      RECT 4.360000 1948.800000 58.125000 1949.900000 ;
      RECT 0.000000 1948.800000 3.460000 1949.900000 ;
      RECT 0.000000 1947.230000 2050.220000 1948.800000 ;
      RECT 1.100000 1946.330000 2050.220000 1947.230000 ;
      RECT 0.000000 1945.940000 2050.220000 1946.330000 ;
      RECT 0.000000 1945.840000 2045.100000 1945.940000 ;
      RECT 0.000000 1943.440000 2.620000 1945.840000 ;
      RECT 2047.700000 1942.350000 2050.220000 1945.940000 ;
      RECT 0.000000 1942.240000 2045.100000 1943.440000 ;
      RECT 2047.700000 1941.450000 2049.120000 1942.350000 ;
      RECT 2044.000000 1939.840000 2045.100000 1942.240000 ;
      RECT 0.000000 1939.840000 6.220000 1942.240000 ;
      RECT 0.000000 1933.895000 2045.100000 1939.840000 ;
      RECT 2031.850000 1931.495000 2045.100000 1933.895000 ;
      RECT 0.000000 1931.495000 16.770000 1933.895000 ;
      RECT 0.000000 1930.295000 2045.100000 1931.495000 ;
      RECT 2028.250000 1927.895000 2045.100000 1930.295000 ;
      RECT 0.000000 1927.895000 20.370000 1930.295000 ;
      RECT 0.000000 1913.530000 2045.100000 1927.895000 ;
      RECT 2047.700000 1912.850000 2050.220000 1941.450000 ;
      RECT 1.100000 1912.630000 2045.100000 1913.530000 ;
      RECT 2047.700000 1911.950000 2049.120000 1912.850000 ;
      RECT 0.000000 1876.740000 2045.100000 1912.630000 ;
      RECT 1.100000 1875.840000 2045.100000 1876.740000 ;
      RECT 2047.700000 1875.350000 2050.220000 1911.950000 ;
      RECT 2047.700000 1874.450000 2049.120000 1875.350000 ;
      RECT 0.000000 1839.950000 2045.100000 1875.840000 ;
      RECT 1.100000 1839.050000 2045.100000 1839.950000 ;
      RECT 2047.700000 1837.850000 2050.220000 1874.450000 ;
      RECT 2047.700000 1836.950000 2049.120000 1837.850000 ;
      RECT 0.000000 1803.160000 2045.100000 1839.050000 ;
      RECT 1.100000 1802.260000 2045.100000 1803.160000 ;
      RECT 2047.700000 1800.355000 2050.220000 1836.950000 ;
      RECT 2047.700000 1799.455000 2049.120000 1800.355000 ;
      RECT 0.000000 1766.370000 2045.100000 1802.260000 ;
      RECT 1.100000 1765.470000 2045.100000 1766.370000 ;
      RECT 2047.700000 1762.855000 2050.220000 1799.455000 ;
      RECT 2047.700000 1761.955000 2049.120000 1762.855000 ;
      RECT 0.000000 1729.580000 2045.100000 1765.470000 ;
      RECT 1.100000 1728.680000 2045.100000 1729.580000 ;
      RECT 2047.700000 1725.360000 2050.220000 1761.955000 ;
      RECT 2047.700000 1724.460000 2049.120000 1725.360000 ;
      RECT 0.000000 1692.790000 2045.100000 1728.680000 ;
      RECT 1.100000 1691.890000 2045.100000 1692.790000 ;
      RECT 2047.700000 1687.860000 2050.220000 1724.460000 ;
      RECT 2047.700000 1686.960000 2049.120000 1687.860000 ;
      RECT 0.000000 1656.000000 2045.100000 1691.890000 ;
      RECT 1.100000 1655.100000 2045.100000 1656.000000 ;
      RECT 2047.700000 1650.360000 2050.220000 1686.960000 ;
      RECT 2047.700000 1649.460000 2049.120000 1650.360000 ;
      RECT 0.000000 1619.210000 2045.100000 1655.100000 ;
      RECT 1.100000 1618.310000 2045.100000 1619.210000 ;
      RECT 2047.700000 1612.865000 2050.220000 1649.460000 ;
      RECT 2047.700000 1611.965000 2049.120000 1612.865000 ;
      RECT 0.000000 1582.420000 2045.100000 1618.310000 ;
      RECT 1.100000 1581.520000 2045.100000 1582.420000 ;
      RECT 2047.700000 1575.365000 2050.220000 1611.965000 ;
      RECT 2047.700000 1574.465000 2049.120000 1575.365000 ;
      RECT 0.000000 1545.630000 2045.100000 1581.520000 ;
      RECT 1.100000 1544.730000 2045.100000 1545.630000 ;
      RECT 2047.700000 1537.870000 2050.220000 1574.465000 ;
      RECT 2047.700000 1536.970000 2049.120000 1537.870000 ;
      RECT 0.000000 1508.840000 2045.100000 1544.730000 ;
      RECT 1.100000 1507.940000 2045.100000 1508.840000 ;
      RECT 2047.700000 1500.370000 2050.220000 1536.970000 ;
      RECT 2047.700000 1499.470000 2049.120000 1500.370000 ;
      RECT 0.000000 1472.050000 2045.100000 1507.940000 ;
      RECT 1.100000 1471.150000 2045.100000 1472.050000 ;
      RECT 2047.700000 1462.870000 2050.220000 1499.470000 ;
      RECT 2047.700000 1461.970000 2049.120000 1462.870000 ;
      RECT 0.000000 1435.260000 2045.100000 1471.150000 ;
      RECT 1.100000 1434.360000 2045.100000 1435.260000 ;
      RECT 2047.700000 1425.375000 2050.220000 1461.970000 ;
      RECT 2047.700000 1424.475000 2049.120000 1425.375000 ;
      RECT 0.000000 1398.470000 2045.100000 1434.360000 ;
      RECT 1.100000 1397.570000 2045.100000 1398.470000 ;
      RECT 2047.700000 1387.875000 2050.220000 1424.475000 ;
      RECT 2047.700000 1386.975000 2049.120000 1387.875000 ;
      RECT 0.000000 1361.680000 2045.100000 1397.570000 ;
      RECT 1.100000 1360.780000 2045.100000 1361.680000 ;
      RECT 2047.700000 1350.380000 2050.220000 1386.975000 ;
      RECT 2047.700000 1349.480000 2049.120000 1350.380000 ;
      RECT 0.000000 1324.890000 2045.100000 1360.780000 ;
      RECT 1.100000 1323.990000 2045.100000 1324.890000 ;
      RECT 2047.700000 1312.880000 2050.220000 1349.480000 ;
      RECT 2047.700000 1311.980000 2049.120000 1312.880000 ;
      RECT 0.000000 1288.100000 2045.100000 1323.990000 ;
      RECT 1.100000 1287.200000 2045.100000 1288.100000 ;
      RECT 2047.700000 1275.380000 2050.220000 1311.980000 ;
      RECT 2047.700000 1274.480000 2049.120000 1275.380000 ;
      RECT 0.000000 1251.310000 2045.100000 1287.200000 ;
      RECT 1.100000 1250.410000 2045.100000 1251.310000 ;
      RECT 2047.700000 1237.885000 2050.220000 1274.480000 ;
      RECT 2047.700000 1236.985000 2049.120000 1237.885000 ;
      RECT 0.000000 1214.520000 2045.100000 1250.410000 ;
      RECT 1.100000 1213.620000 2045.100000 1214.520000 ;
      RECT 2047.700000 1200.385000 2050.220000 1236.985000 ;
      RECT 2047.700000 1199.485000 2049.120000 1200.385000 ;
      RECT 0.000000 1177.730000 2045.100000 1213.620000 ;
      RECT 1.100000 1176.830000 2045.100000 1177.730000 ;
      RECT 2047.700000 1162.890000 2050.220000 1199.485000 ;
      RECT 2047.700000 1161.990000 2049.120000 1162.890000 ;
      RECT 0.000000 1140.940000 2045.100000 1176.830000 ;
      RECT 1.100000 1140.040000 2045.100000 1140.940000 ;
      RECT 2047.700000 1125.390000 2050.220000 1161.990000 ;
      RECT 2047.700000 1124.490000 2049.120000 1125.390000 ;
      RECT 0.000000 1104.150000 2045.100000 1140.040000 ;
      RECT 1.100000 1103.250000 2045.100000 1104.150000 ;
      RECT 2047.700000 1087.890000 2050.220000 1124.490000 ;
      RECT 2047.700000 1086.990000 2049.120000 1087.890000 ;
      RECT 0.000000 1067.360000 2045.100000 1103.250000 ;
      RECT 1.100000 1066.460000 2045.100000 1067.360000 ;
      RECT 2047.700000 1050.395000 2050.220000 1086.990000 ;
      RECT 2047.700000 1049.495000 2049.120000 1050.395000 ;
      RECT 0.000000 1030.570000 2045.100000 1066.460000 ;
      RECT 1.100000 1029.670000 2045.100000 1030.570000 ;
      RECT 2047.700000 1012.895000 2050.220000 1049.495000 ;
      RECT 2047.700000 1011.995000 2049.120000 1012.895000 ;
      RECT 0.000000 993.780000 2045.100000 1029.670000 ;
      RECT 1.100000 992.880000 2045.100000 993.780000 ;
      RECT 2047.700000 975.400000 2050.220000 1011.995000 ;
      RECT 2047.700000 974.500000 2049.120000 975.400000 ;
      RECT 0.000000 956.990000 2045.100000 992.880000 ;
      RECT 1.100000 956.090000 2045.100000 956.990000 ;
      RECT 2047.700000 937.900000 2050.220000 974.500000 ;
      RECT 2047.700000 937.000000 2049.120000 937.900000 ;
      RECT 0.000000 920.200000 2045.100000 956.090000 ;
      RECT 1.100000 919.300000 2045.100000 920.200000 ;
      RECT 2047.700000 900.400000 2050.220000 937.000000 ;
      RECT 2047.700000 899.500000 2049.120000 900.400000 ;
      RECT 0.000000 883.410000 2045.100000 919.300000 ;
      RECT 1.100000 882.510000 2045.100000 883.410000 ;
      RECT 2047.700000 862.905000 2050.220000 899.500000 ;
      RECT 2047.700000 862.005000 2049.120000 862.905000 ;
      RECT 0.000000 846.620000 2045.100000 882.510000 ;
      RECT 1.100000 845.720000 2045.100000 846.620000 ;
      RECT 2047.700000 825.405000 2050.220000 862.005000 ;
      RECT 2047.700000 824.505000 2049.120000 825.405000 ;
      RECT 0.000000 809.830000 2045.100000 845.720000 ;
      RECT 1.100000 808.930000 2045.100000 809.830000 ;
      RECT 2047.700000 787.910000 2050.220000 824.505000 ;
      RECT 2047.700000 787.010000 2049.120000 787.910000 ;
      RECT 0.000000 773.040000 2045.100000 808.930000 ;
      RECT 1.100000 772.140000 2045.100000 773.040000 ;
      RECT 2047.700000 750.410000 2050.220000 787.010000 ;
      RECT 2047.700000 749.510000 2049.120000 750.410000 ;
      RECT 0.000000 736.250000 2045.100000 772.140000 ;
      RECT 1.100000 735.350000 2045.100000 736.250000 ;
      RECT 2047.700000 712.910000 2050.220000 749.510000 ;
      RECT 2047.700000 712.010000 2049.120000 712.910000 ;
      RECT 0.000000 699.460000 2045.100000 735.350000 ;
      RECT 1.100000 698.560000 2045.100000 699.460000 ;
      RECT 2047.700000 675.415000 2050.220000 712.010000 ;
      RECT 2047.700000 674.515000 2049.120000 675.415000 ;
      RECT 0.000000 662.670000 2045.100000 698.560000 ;
      RECT 1.100000 661.770000 2045.100000 662.670000 ;
      RECT 2047.700000 637.915000 2050.220000 674.515000 ;
      RECT 2047.700000 637.015000 2049.120000 637.915000 ;
      RECT 0.000000 625.880000 2045.100000 661.770000 ;
      RECT 1.100000 624.980000 2045.100000 625.880000 ;
      RECT 2047.700000 600.420000 2050.220000 637.015000 ;
      RECT 2047.700000 599.520000 2049.120000 600.420000 ;
      RECT 0.000000 589.090000 2045.100000 624.980000 ;
      RECT 1.100000 588.190000 2045.100000 589.090000 ;
      RECT 2047.700000 562.920000 2050.220000 599.520000 ;
      RECT 2047.700000 562.020000 2049.120000 562.920000 ;
      RECT 0.000000 552.300000 2045.100000 588.190000 ;
      RECT 1.100000 551.400000 2045.100000 552.300000 ;
      RECT 2047.700000 525.420000 2050.220000 562.020000 ;
      RECT 2047.700000 524.520000 2049.120000 525.420000 ;
      RECT 0.000000 515.510000 2045.100000 551.400000 ;
      RECT 1.100000 514.610000 2045.100000 515.510000 ;
      RECT 2047.700000 487.925000 2050.220000 524.520000 ;
      RECT 2047.700000 487.025000 2049.120000 487.925000 ;
      RECT 0.000000 478.720000 2045.100000 514.610000 ;
      RECT 1.100000 477.820000 2045.100000 478.720000 ;
      RECT 2047.700000 450.425000 2050.220000 487.025000 ;
      RECT 2047.700000 449.525000 2049.120000 450.425000 ;
      RECT 0.000000 441.930000 2045.100000 477.820000 ;
      RECT 1.100000 441.030000 2045.100000 441.930000 ;
      RECT 2047.700000 412.930000 2050.220000 449.525000 ;
      RECT 2047.700000 412.030000 2049.120000 412.930000 ;
      RECT 0.000000 405.140000 2045.100000 441.030000 ;
      RECT 1.100000 404.240000 2045.100000 405.140000 ;
      RECT 2047.700000 375.430000 2050.220000 412.030000 ;
      RECT 2047.700000 374.530000 2049.120000 375.430000 ;
      RECT 0.000000 368.350000 2045.100000 404.240000 ;
      RECT 1.100000 367.450000 2045.100000 368.350000 ;
      RECT 2047.700000 337.930000 2050.220000 374.530000 ;
      RECT 2047.700000 337.030000 2049.120000 337.930000 ;
      RECT 0.000000 331.560000 2045.100000 367.450000 ;
      RECT 1.100000 330.660000 2045.100000 331.560000 ;
      RECT 2047.700000 300.435000 2050.220000 337.030000 ;
      RECT 2047.700000 299.535000 2049.120000 300.435000 ;
      RECT 0.000000 294.770000 2045.100000 330.660000 ;
      RECT 1.100000 293.870000 2045.100000 294.770000 ;
      RECT 2047.700000 262.935000 2050.220000 299.535000 ;
      RECT 2047.700000 262.035000 2049.120000 262.935000 ;
      RECT 0.000000 257.980000 2045.100000 293.870000 ;
      RECT 1.100000 257.080000 2045.100000 257.980000 ;
      RECT 2047.700000 225.440000 2050.220000 262.035000 ;
      RECT 2047.700000 224.540000 2049.120000 225.440000 ;
      RECT 0.000000 221.190000 2045.100000 257.080000 ;
      RECT 1.100000 220.290000 2045.100000 221.190000 ;
      RECT 2047.700000 187.940000 2050.220000 224.540000 ;
      RECT 2047.700000 187.040000 2049.120000 187.940000 ;
      RECT 0.000000 184.400000 2045.100000 220.290000 ;
      RECT 1.100000 183.500000 2045.100000 184.400000 ;
      RECT 2047.700000 150.440000 2050.220000 187.040000 ;
      RECT 2047.700000 149.540000 2049.120000 150.440000 ;
      RECT 0.000000 147.610000 2045.100000 183.500000 ;
      RECT 1.100000 146.710000 2045.100000 147.610000 ;
      RECT 2047.700000 112.945000 2050.220000 149.540000 ;
      RECT 2047.700000 112.045000 2049.120000 112.945000 ;
      RECT 0.000000 110.820000 2045.100000 146.710000 ;
      RECT 1.100000 109.920000 2045.100000 110.820000 ;
      RECT 2047.700000 75.445000 2050.220000 112.045000 ;
      RECT 2047.700000 74.545000 2049.120000 75.445000 ;
      RECT 0.000000 74.030000 2045.100000 109.920000 ;
      RECT 1.100000 73.130000 2045.100000 74.030000 ;
      RECT 2047.700000 37.950000 2050.220000 74.545000 ;
      RECT 0.000000 37.240000 2045.100000 73.130000 ;
      RECT 2047.700000 37.050000 2049.120000 37.950000 ;
      RECT 1.100000 36.340000 2045.100000 37.240000 ;
      RECT 0.000000 24.975000 2045.100000 36.340000 ;
      RECT 2028.250000 22.575000 2045.100000 24.975000 ;
      RECT 0.000000 22.575000 20.370000 24.975000 ;
      RECT 0.000000 21.375000 2045.100000 22.575000 ;
      RECT 2031.850000 18.975000 2045.100000 21.375000 ;
      RECT 0.000000 18.975000 16.770000 21.375000 ;
      RECT 2047.700000 10.480000 2050.220000 37.050000 ;
      RECT 2047.700000 9.580000 2049.120000 10.480000 ;
      RECT 0.000000 8.360000 2045.100000 18.975000 ;
      RECT 0.000000 8.040000 6.220000 8.360000 ;
      RECT 1.100000 7.140000 6.220000 8.040000 ;
      RECT 2044.000000 5.960000 2045.100000 8.360000 ;
      RECT 0.000000 5.960000 6.220000 7.140000 ;
      RECT 0.000000 4.760000 2045.100000 5.960000 ;
      RECT 0.000000 2.360000 2.620000 4.760000 ;
      RECT 2047.700000 2.260000 2050.220000 9.580000 ;
      RECT 0.000000 2.260000 2045.100000 2.360000 ;
      RECT 0.000000 1.100000 2050.220000 2.260000 ;
      RECT 2048.600000 0.000000 2050.220000 1.100000 ;
      RECT 2046.185000 0.000000 2047.700000 1.100000 ;
      RECT 2042.030000 0.000000 2045.285000 1.100000 ;
      RECT 2037.870000 0.000000 2041.130000 1.100000 ;
      RECT 2033.710000 0.000000 2036.970000 1.100000 ;
      RECT 2029.555000 0.000000 2032.810000 1.100000 ;
      RECT 2025.395000 0.000000 2028.655000 1.100000 ;
      RECT 2021.240000 0.000000 2024.495000 1.100000 ;
      RECT 2017.080000 0.000000 2020.340000 1.100000 ;
      RECT 2012.920000 0.000000 2016.180000 1.100000 ;
      RECT 2008.765000 0.000000 2012.020000 1.100000 ;
      RECT 2004.605000 0.000000 2007.865000 1.100000 ;
      RECT 2000.450000 0.000000 2003.705000 1.100000 ;
      RECT 1996.290000 0.000000 1999.550000 1.100000 ;
      RECT 1992.130000 0.000000 1995.390000 1.100000 ;
      RECT 1987.975000 0.000000 1991.230000 1.100000 ;
      RECT 1983.815000 0.000000 1987.075000 1.100000 ;
      RECT 1979.660000 0.000000 1982.915000 1.100000 ;
      RECT 1975.500000 0.000000 1978.760000 1.100000 ;
      RECT 1971.340000 0.000000 1974.600000 1.100000 ;
      RECT 1967.185000 0.000000 1970.440000 1.100000 ;
      RECT 1963.025000 0.000000 1966.285000 1.100000 ;
      RECT 1958.870000 0.000000 1962.125000 1.100000 ;
      RECT 1954.710000 0.000000 1957.970000 1.100000 ;
      RECT 1950.550000 0.000000 1953.810000 1.100000 ;
      RECT 1946.395000 0.000000 1949.650000 1.100000 ;
      RECT 1942.235000 0.000000 1945.495000 1.100000 ;
      RECT 1938.080000 0.000000 1941.335000 1.100000 ;
      RECT 1933.920000 0.000000 1937.180000 1.100000 ;
      RECT 1929.760000 0.000000 1933.020000 1.100000 ;
      RECT 1925.605000 0.000000 1928.860000 1.100000 ;
      RECT 1921.445000 0.000000 1924.705000 1.100000 ;
      RECT 1917.290000 0.000000 1920.545000 1.100000 ;
      RECT 1913.130000 0.000000 1916.390000 1.100000 ;
      RECT 1908.970000 0.000000 1912.230000 1.100000 ;
      RECT 1904.815000 0.000000 1908.070000 1.100000 ;
      RECT 1900.655000 0.000000 1903.915000 1.100000 ;
      RECT 1896.500000 0.000000 1899.755000 1.100000 ;
      RECT 1892.340000 0.000000 1895.600000 1.100000 ;
      RECT 1888.180000 0.000000 1891.440000 1.100000 ;
      RECT 1884.025000 0.000000 1887.280000 1.100000 ;
      RECT 1879.865000 0.000000 1883.125000 1.100000 ;
      RECT 1875.710000 0.000000 1878.965000 1.100000 ;
      RECT 1871.550000 0.000000 1874.810000 1.100000 ;
      RECT 1867.390000 0.000000 1870.650000 1.100000 ;
      RECT 1863.235000 0.000000 1866.490000 1.100000 ;
      RECT 1859.075000 0.000000 1862.335000 1.100000 ;
      RECT 1854.920000 0.000000 1858.175000 1.100000 ;
      RECT 1850.760000 0.000000 1854.020000 1.100000 ;
      RECT 1846.600000 0.000000 1849.860000 1.100000 ;
      RECT 1842.445000 0.000000 1845.700000 1.100000 ;
      RECT 1838.285000 0.000000 1841.545000 1.100000 ;
      RECT 1834.130000 0.000000 1837.385000 1.100000 ;
      RECT 1829.970000 0.000000 1833.230000 1.100000 ;
      RECT 1825.810000 0.000000 1829.070000 1.100000 ;
      RECT 1821.655000 0.000000 1824.910000 1.100000 ;
      RECT 1817.495000 0.000000 1820.755000 1.100000 ;
      RECT 1813.340000 0.000000 1816.595000 1.100000 ;
      RECT 1809.180000 0.000000 1812.440000 1.100000 ;
      RECT 1805.020000 0.000000 1808.280000 1.100000 ;
      RECT 1800.865000 0.000000 1804.120000 1.100000 ;
      RECT 1796.705000 0.000000 1799.965000 1.100000 ;
      RECT 1792.550000 0.000000 1795.805000 1.100000 ;
      RECT 1788.390000 0.000000 1791.650000 1.100000 ;
      RECT 1784.230000 0.000000 1787.490000 1.100000 ;
      RECT 1780.075000 0.000000 1783.330000 1.100000 ;
      RECT 1775.915000 0.000000 1779.175000 1.100000 ;
      RECT 1771.760000 0.000000 1775.015000 1.100000 ;
      RECT 1767.600000 0.000000 1770.860000 1.100000 ;
      RECT 1763.440000 0.000000 1766.700000 1.100000 ;
      RECT 1759.285000 0.000000 1762.540000 1.100000 ;
      RECT 1755.125000 0.000000 1758.385000 1.100000 ;
      RECT 1750.970000 0.000000 1754.225000 1.100000 ;
      RECT 1746.810000 0.000000 1750.070000 1.100000 ;
      RECT 1742.650000 0.000000 1745.910000 1.100000 ;
      RECT 1738.495000 0.000000 1741.750000 1.100000 ;
      RECT 1734.335000 0.000000 1737.595000 1.100000 ;
      RECT 1730.180000 0.000000 1733.435000 1.100000 ;
      RECT 1726.020000 0.000000 1729.280000 1.100000 ;
      RECT 1721.860000 0.000000 1725.120000 1.100000 ;
      RECT 1717.705000 0.000000 1720.960000 1.100000 ;
      RECT 1713.545000 0.000000 1716.805000 1.100000 ;
      RECT 1709.390000 0.000000 1712.645000 1.100000 ;
      RECT 1705.230000 0.000000 1708.490000 1.100000 ;
      RECT 1701.070000 0.000000 1704.330000 1.100000 ;
      RECT 1696.915000 0.000000 1700.170000 1.100000 ;
      RECT 1692.755000 0.000000 1696.015000 1.100000 ;
      RECT 1688.600000 0.000000 1691.855000 1.100000 ;
      RECT 1684.440000 0.000000 1687.700000 1.100000 ;
      RECT 1680.280000 0.000000 1683.540000 1.100000 ;
      RECT 1676.125000 0.000000 1679.380000 1.100000 ;
      RECT 1671.965000 0.000000 1675.225000 1.100000 ;
      RECT 1667.810000 0.000000 1671.065000 1.100000 ;
      RECT 1663.650000 0.000000 1666.910000 1.100000 ;
      RECT 1659.490000 0.000000 1662.750000 1.100000 ;
      RECT 1655.335000 0.000000 1658.590000 1.100000 ;
      RECT 1651.175000 0.000000 1654.435000 1.100000 ;
      RECT 1647.020000 0.000000 1650.275000 1.100000 ;
      RECT 1642.860000 0.000000 1646.120000 1.100000 ;
      RECT 1638.700000 0.000000 1641.960000 1.100000 ;
      RECT 1634.545000 0.000000 1637.800000 1.100000 ;
      RECT 1630.385000 0.000000 1633.645000 1.100000 ;
      RECT 1626.230000 0.000000 1629.485000 1.100000 ;
      RECT 1622.070000 0.000000 1625.330000 1.100000 ;
      RECT 1617.910000 0.000000 1621.170000 1.100000 ;
      RECT 1613.755000 0.000000 1617.010000 1.100000 ;
      RECT 1609.595000 0.000000 1612.855000 1.100000 ;
      RECT 1605.440000 0.000000 1608.695000 1.100000 ;
      RECT 1601.280000 0.000000 1604.540000 1.100000 ;
      RECT 1597.120000 0.000000 1600.380000 1.100000 ;
      RECT 1592.965000 0.000000 1596.220000 1.100000 ;
      RECT 1588.805000 0.000000 1592.065000 1.100000 ;
      RECT 1584.650000 0.000000 1587.905000 1.100000 ;
      RECT 1580.490000 0.000000 1583.750000 1.100000 ;
      RECT 1576.330000 0.000000 1579.590000 1.100000 ;
      RECT 1572.175000 0.000000 1575.430000 1.100000 ;
      RECT 1568.015000 0.000000 1571.275000 1.100000 ;
      RECT 1563.860000 0.000000 1567.115000 1.100000 ;
      RECT 1559.700000 0.000000 1562.960000 1.100000 ;
      RECT 1555.540000 0.000000 1558.800000 1.100000 ;
      RECT 1551.385000 0.000000 1554.640000 1.100000 ;
      RECT 1547.225000 0.000000 1550.485000 1.100000 ;
      RECT 1543.070000 0.000000 1546.325000 1.100000 ;
      RECT 1538.910000 0.000000 1542.170000 1.100000 ;
      RECT 1534.750000 0.000000 1538.010000 1.100000 ;
      RECT 1530.595000 0.000000 1533.850000 1.100000 ;
      RECT 1526.435000 0.000000 1529.695000 1.100000 ;
      RECT 1522.280000 0.000000 1525.535000 1.100000 ;
      RECT 1518.120000 0.000000 1521.380000 1.100000 ;
      RECT 1513.960000 0.000000 1517.220000 1.100000 ;
      RECT 1509.805000 0.000000 1513.060000 1.100000 ;
      RECT 1505.645000 0.000000 1508.905000 1.100000 ;
      RECT 1501.490000 0.000000 1504.745000 1.100000 ;
      RECT 1497.330000 0.000000 1500.590000 1.100000 ;
      RECT 1493.170000 0.000000 1496.430000 1.100000 ;
      RECT 1489.015000 0.000000 1492.270000 1.100000 ;
      RECT 1484.855000 0.000000 1488.115000 1.100000 ;
      RECT 1480.700000 0.000000 1483.955000 1.100000 ;
      RECT 1476.540000 0.000000 1479.800000 1.100000 ;
      RECT 1472.380000 0.000000 1475.640000 1.100000 ;
      RECT 1468.225000 0.000000 1471.480000 1.100000 ;
      RECT 1464.065000 0.000000 1467.325000 1.100000 ;
      RECT 1459.910000 0.000000 1463.165000 1.100000 ;
      RECT 1455.750000 0.000000 1459.010000 1.100000 ;
      RECT 1451.590000 0.000000 1454.850000 1.100000 ;
      RECT 1447.435000 0.000000 1450.690000 1.100000 ;
      RECT 1443.275000 0.000000 1446.535000 1.100000 ;
      RECT 1439.120000 0.000000 1442.375000 1.100000 ;
      RECT 1434.960000 0.000000 1438.220000 1.100000 ;
      RECT 1430.800000 0.000000 1434.060000 1.100000 ;
      RECT 1426.645000 0.000000 1429.900000 1.100000 ;
      RECT 1422.485000 0.000000 1425.745000 1.100000 ;
      RECT 1418.330000 0.000000 1421.585000 1.100000 ;
      RECT 1414.170000 0.000000 1417.430000 1.100000 ;
      RECT 1410.010000 0.000000 1413.270000 1.100000 ;
      RECT 1405.855000 0.000000 1409.110000 1.100000 ;
      RECT 1401.695000 0.000000 1404.955000 1.100000 ;
      RECT 1397.540000 0.000000 1400.795000 1.100000 ;
      RECT 1393.380000 0.000000 1396.640000 1.100000 ;
      RECT 1389.220000 0.000000 1392.480000 1.100000 ;
      RECT 1385.065000 0.000000 1388.320000 1.100000 ;
      RECT 1380.905000 0.000000 1384.165000 1.100000 ;
      RECT 1376.750000 0.000000 1380.005000 1.100000 ;
      RECT 1372.590000 0.000000 1375.850000 1.100000 ;
      RECT 1368.430000 0.000000 1371.690000 1.100000 ;
      RECT 1364.275000 0.000000 1367.530000 1.100000 ;
      RECT 1360.115000 0.000000 1363.375000 1.100000 ;
      RECT 1355.960000 0.000000 1359.215000 1.100000 ;
      RECT 1351.800000 0.000000 1355.060000 1.100000 ;
      RECT 1347.640000 0.000000 1350.900000 1.100000 ;
      RECT 1343.485000 0.000000 1346.740000 1.100000 ;
      RECT 1339.325000 0.000000 1342.585000 1.100000 ;
      RECT 1335.170000 0.000000 1338.425000 1.100000 ;
      RECT 1331.010000 0.000000 1334.270000 1.100000 ;
      RECT 1326.850000 0.000000 1330.110000 1.100000 ;
      RECT 1322.695000 0.000000 1325.950000 1.100000 ;
      RECT 1318.535000 0.000000 1321.795000 1.100000 ;
      RECT 1314.380000 0.000000 1317.635000 1.100000 ;
      RECT 1310.220000 0.000000 1313.480000 1.100000 ;
      RECT 1306.060000 0.000000 1309.320000 1.100000 ;
      RECT 1301.905000 0.000000 1305.160000 1.100000 ;
      RECT 1297.745000 0.000000 1301.005000 1.100000 ;
      RECT 1293.590000 0.000000 1296.845000 1.100000 ;
      RECT 1289.430000 0.000000 1292.690000 1.100000 ;
      RECT 1285.270000 0.000000 1288.530000 1.100000 ;
      RECT 1281.115000 0.000000 1284.370000 1.100000 ;
      RECT 1276.955000 0.000000 1280.215000 1.100000 ;
      RECT 1272.800000 0.000000 1276.055000 1.100000 ;
      RECT 1268.640000 0.000000 1271.900000 1.100000 ;
      RECT 1264.480000 0.000000 1267.740000 1.100000 ;
      RECT 1260.325000 0.000000 1263.580000 1.100000 ;
      RECT 1256.165000 0.000000 1259.425000 1.100000 ;
      RECT 1252.010000 0.000000 1255.265000 1.100000 ;
      RECT 1247.850000 0.000000 1251.110000 1.100000 ;
      RECT 1243.690000 0.000000 1246.950000 1.100000 ;
      RECT 1239.535000 0.000000 1242.790000 1.100000 ;
      RECT 1235.375000 0.000000 1238.635000 1.100000 ;
      RECT 1231.220000 0.000000 1234.475000 1.100000 ;
      RECT 1227.060000 0.000000 1230.320000 1.100000 ;
      RECT 1222.900000 0.000000 1226.160000 1.100000 ;
      RECT 1218.745000 0.000000 1222.000000 1.100000 ;
      RECT 1214.585000 0.000000 1217.845000 1.100000 ;
      RECT 1210.430000 0.000000 1213.685000 1.100000 ;
      RECT 1206.270000 0.000000 1209.530000 1.100000 ;
      RECT 1202.110000 0.000000 1205.370000 1.100000 ;
      RECT 1197.955000 0.000000 1201.210000 1.100000 ;
      RECT 1193.795000 0.000000 1197.055000 1.100000 ;
      RECT 1189.640000 0.000000 1192.895000 1.100000 ;
      RECT 1185.480000 0.000000 1188.740000 1.100000 ;
      RECT 1181.320000 0.000000 1184.580000 1.100000 ;
      RECT 1177.165000 0.000000 1180.420000 1.100000 ;
      RECT 1173.005000 0.000000 1176.265000 1.100000 ;
      RECT 1168.850000 0.000000 1172.105000 1.100000 ;
      RECT 1164.690000 0.000000 1167.950000 1.100000 ;
      RECT 1160.530000 0.000000 1163.790000 1.100000 ;
      RECT 1156.375000 0.000000 1159.630000 1.100000 ;
      RECT 1152.215000 0.000000 1155.475000 1.100000 ;
      RECT 1148.060000 0.000000 1151.315000 1.100000 ;
      RECT 1143.900000 0.000000 1147.160000 1.100000 ;
      RECT 1139.740000 0.000000 1143.000000 1.100000 ;
      RECT 1135.585000 0.000000 1138.840000 1.100000 ;
      RECT 1131.425000 0.000000 1134.685000 1.100000 ;
      RECT 1127.270000 0.000000 1130.525000 1.100000 ;
      RECT 1123.110000 0.000000 1126.370000 1.100000 ;
      RECT 1118.950000 0.000000 1122.210000 1.100000 ;
      RECT 1114.795000 0.000000 1118.050000 1.100000 ;
      RECT 1110.635000 0.000000 1113.895000 1.100000 ;
      RECT 1106.480000 0.000000 1109.735000 1.100000 ;
      RECT 1102.320000 0.000000 1105.580000 1.100000 ;
      RECT 1098.160000 0.000000 1101.420000 1.100000 ;
      RECT 1094.005000 0.000000 1097.260000 1.100000 ;
      RECT 1089.845000 0.000000 1093.105000 1.100000 ;
      RECT 1085.690000 0.000000 1088.945000 1.100000 ;
      RECT 1081.530000 0.000000 1084.790000 1.100000 ;
      RECT 1077.370000 0.000000 1080.630000 1.100000 ;
      RECT 1073.215000 0.000000 1076.470000 1.100000 ;
      RECT 1069.055000 0.000000 1072.315000 1.100000 ;
      RECT 1064.900000 0.000000 1068.155000 1.100000 ;
      RECT 1060.740000 0.000000 1064.000000 1.100000 ;
      RECT 1056.580000 0.000000 1059.840000 1.100000 ;
      RECT 1052.425000 0.000000 1055.680000 1.100000 ;
      RECT 1048.265000 0.000000 1051.525000 1.100000 ;
      RECT 1044.110000 0.000000 1047.365000 1.100000 ;
      RECT 1039.950000 0.000000 1043.210000 1.100000 ;
      RECT 1035.790000 0.000000 1039.050000 1.100000 ;
      RECT 1031.635000 0.000000 1034.890000 1.100000 ;
      RECT 1027.475000 0.000000 1030.735000 1.100000 ;
      RECT 1023.320000 0.000000 1026.575000 1.100000 ;
      RECT 1019.160000 0.000000 1022.420000 1.100000 ;
      RECT 1015.000000 0.000000 1018.260000 1.100000 ;
      RECT 1010.845000 0.000000 1014.100000 1.100000 ;
      RECT 1006.685000 0.000000 1009.945000 1.100000 ;
      RECT 1002.530000 0.000000 1005.785000 1.100000 ;
      RECT 998.370000 0.000000 1001.630000 1.100000 ;
      RECT 994.210000 0.000000 997.470000 1.100000 ;
      RECT 990.055000 0.000000 993.310000 1.100000 ;
      RECT 985.895000 0.000000 989.155000 1.100000 ;
      RECT 981.740000 0.000000 984.995000 1.100000 ;
      RECT 977.580000 0.000000 980.840000 1.100000 ;
      RECT 973.420000 0.000000 976.680000 1.100000 ;
      RECT 969.265000 0.000000 972.520000 1.100000 ;
      RECT 965.105000 0.000000 968.365000 1.100000 ;
      RECT 960.950000 0.000000 964.205000 1.100000 ;
      RECT 956.790000 0.000000 960.050000 1.100000 ;
      RECT 952.630000 0.000000 955.890000 1.100000 ;
      RECT 948.475000 0.000000 951.730000 1.100000 ;
      RECT 944.315000 0.000000 947.575000 1.100000 ;
      RECT 940.160000 0.000000 943.415000 1.100000 ;
      RECT 936.000000 0.000000 939.260000 1.100000 ;
      RECT 931.840000 0.000000 935.100000 1.100000 ;
      RECT 927.685000 0.000000 930.940000 1.100000 ;
      RECT 923.525000 0.000000 926.785000 1.100000 ;
      RECT 919.370000 0.000000 922.625000 1.100000 ;
      RECT 915.210000 0.000000 918.470000 1.100000 ;
      RECT 911.050000 0.000000 914.310000 1.100000 ;
      RECT 906.895000 0.000000 910.150000 1.100000 ;
      RECT 902.735000 0.000000 905.995000 1.100000 ;
      RECT 898.580000 0.000000 901.835000 1.100000 ;
      RECT 894.420000 0.000000 897.680000 1.100000 ;
      RECT 890.260000 0.000000 893.520000 1.100000 ;
      RECT 886.105000 0.000000 889.360000 1.100000 ;
      RECT 881.945000 0.000000 885.205000 1.100000 ;
      RECT 877.790000 0.000000 881.045000 1.100000 ;
      RECT 873.630000 0.000000 876.890000 1.100000 ;
      RECT 869.470000 0.000000 872.730000 1.100000 ;
      RECT 865.315000 0.000000 868.570000 1.100000 ;
      RECT 861.155000 0.000000 864.415000 1.100000 ;
      RECT 857.000000 0.000000 860.255000 1.100000 ;
      RECT 852.840000 0.000000 856.100000 1.100000 ;
      RECT 848.680000 0.000000 851.940000 1.100000 ;
      RECT 844.525000 0.000000 847.780000 1.100000 ;
      RECT 840.365000 0.000000 843.625000 1.100000 ;
      RECT 836.210000 0.000000 839.465000 1.100000 ;
      RECT 832.050000 0.000000 835.310000 1.100000 ;
      RECT 827.890000 0.000000 831.150000 1.100000 ;
      RECT 823.735000 0.000000 826.990000 1.100000 ;
      RECT 819.575000 0.000000 822.835000 1.100000 ;
      RECT 815.420000 0.000000 818.675000 1.100000 ;
      RECT 811.260000 0.000000 814.520000 1.100000 ;
      RECT 807.100000 0.000000 810.360000 1.100000 ;
      RECT 802.945000 0.000000 806.200000 1.100000 ;
      RECT 798.785000 0.000000 802.045000 1.100000 ;
      RECT 794.630000 0.000000 797.885000 1.100000 ;
      RECT 790.470000 0.000000 793.730000 1.100000 ;
      RECT 786.310000 0.000000 789.570000 1.100000 ;
      RECT 782.155000 0.000000 785.410000 1.100000 ;
      RECT 777.995000 0.000000 781.255000 1.100000 ;
      RECT 773.840000 0.000000 777.095000 1.100000 ;
      RECT 769.680000 0.000000 772.940000 1.100000 ;
      RECT 765.520000 0.000000 768.780000 1.100000 ;
      RECT 761.365000 0.000000 764.620000 1.100000 ;
      RECT 757.205000 0.000000 760.465000 1.100000 ;
      RECT 753.050000 0.000000 756.305000 1.100000 ;
      RECT 748.890000 0.000000 752.150000 1.100000 ;
      RECT 744.730000 0.000000 747.990000 1.100000 ;
      RECT 740.575000 0.000000 743.830000 1.100000 ;
      RECT 736.415000 0.000000 739.675000 1.100000 ;
      RECT 732.260000 0.000000 735.515000 1.100000 ;
      RECT 728.100000 0.000000 731.360000 1.100000 ;
      RECT 723.940000 0.000000 727.200000 1.100000 ;
      RECT 719.785000 0.000000 723.040000 1.100000 ;
      RECT 715.625000 0.000000 718.885000 1.100000 ;
      RECT 711.470000 0.000000 714.725000 1.100000 ;
      RECT 707.310000 0.000000 710.570000 1.100000 ;
      RECT 703.150000 0.000000 706.410000 1.100000 ;
      RECT 698.995000 0.000000 702.250000 1.100000 ;
      RECT 694.835000 0.000000 698.095000 1.100000 ;
      RECT 690.680000 0.000000 693.935000 1.100000 ;
      RECT 686.520000 0.000000 689.780000 1.100000 ;
      RECT 682.360000 0.000000 685.620000 1.100000 ;
      RECT 678.205000 0.000000 681.460000 1.100000 ;
      RECT 674.045000 0.000000 677.305000 1.100000 ;
      RECT 669.890000 0.000000 673.145000 1.100000 ;
      RECT 665.730000 0.000000 668.990000 1.100000 ;
      RECT 661.570000 0.000000 664.830000 1.100000 ;
      RECT 657.415000 0.000000 660.670000 1.100000 ;
      RECT 653.255000 0.000000 656.515000 1.100000 ;
      RECT 649.100000 0.000000 652.355000 1.100000 ;
      RECT 644.940000 0.000000 648.200000 1.100000 ;
      RECT 640.780000 0.000000 644.040000 1.100000 ;
      RECT 636.625000 0.000000 639.880000 1.100000 ;
      RECT 632.465000 0.000000 635.725000 1.100000 ;
      RECT 628.310000 0.000000 631.565000 1.100000 ;
      RECT 624.150000 0.000000 627.410000 1.100000 ;
      RECT 619.990000 0.000000 623.250000 1.100000 ;
      RECT 615.835000 0.000000 619.090000 1.100000 ;
      RECT 611.675000 0.000000 614.935000 1.100000 ;
      RECT 607.520000 0.000000 610.775000 1.100000 ;
      RECT 603.360000 0.000000 606.620000 1.100000 ;
      RECT 599.200000 0.000000 602.460000 1.100000 ;
      RECT 595.045000 0.000000 598.300000 1.100000 ;
      RECT 590.885000 0.000000 594.145000 1.100000 ;
      RECT 586.730000 0.000000 589.985000 1.100000 ;
      RECT 582.570000 0.000000 585.830000 1.100000 ;
      RECT 578.410000 0.000000 581.670000 1.100000 ;
      RECT 574.255000 0.000000 577.510000 1.100000 ;
      RECT 570.095000 0.000000 573.355000 1.100000 ;
      RECT 565.940000 0.000000 569.195000 1.100000 ;
      RECT 561.780000 0.000000 565.040000 1.100000 ;
      RECT 557.620000 0.000000 560.880000 1.100000 ;
      RECT 553.465000 0.000000 556.720000 1.100000 ;
      RECT 549.305000 0.000000 552.565000 1.100000 ;
      RECT 545.150000 0.000000 548.405000 1.100000 ;
      RECT 540.990000 0.000000 544.250000 1.100000 ;
      RECT 536.830000 0.000000 540.090000 1.100000 ;
      RECT 532.675000 0.000000 535.930000 1.100000 ;
      RECT 528.515000 0.000000 531.775000 1.100000 ;
      RECT 524.360000 0.000000 527.615000 1.100000 ;
      RECT 520.200000 0.000000 523.460000 1.100000 ;
      RECT 516.040000 0.000000 519.300000 1.100000 ;
      RECT 511.885000 0.000000 515.140000 1.100000 ;
      RECT 507.725000 0.000000 510.985000 1.100000 ;
      RECT 503.570000 0.000000 506.825000 1.100000 ;
      RECT 499.410000 0.000000 502.670000 1.100000 ;
      RECT 495.250000 0.000000 498.510000 1.100000 ;
      RECT 491.095000 0.000000 494.350000 1.100000 ;
      RECT 486.935000 0.000000 490.195000 1.100000 ;
      RECT 482.780000 0.000000 486.035000 1.100000 ;
      RECT 478.620000 0.000000 481.880000 1.100000 ;
      RECT 474.460000 0.000000 477.720000 1.100000 ;
      RECT 470.305000 0.000000 473.560000 1.100000 ;
      RECT 466.145000 0.000000 469.405000 1.100000 ;
      RECT 461.990000 0.000000 465.245000 1.100000 ;
      RECT 457.830000 0.000000 461.090000 1.100000 ;
      RECT 453.670000 0.000000 456.930000 1.100000 ;
      RECT 449.515000 0.000000 452.770000 1.100000 ;
      RECT 445.355000 0.000000 448.615000 1.100000 ;
      RECT 441.200000 0.000000 444.455000 1.100000 ;
      RECT 437.040000 0.000000 440.300000 1.100000 ;
      RECT 432.880000 0.000000 436.140000 1.100000 ;
      RECT 428.725000 0.000000 431.980000 1.100000 ;
      RECT 424.565000 0.000000 427.825000 1.100000 ;
      RECT 420.410000 0.000000 423.665000 1.100000 ;
      RECT 416.250000 0.000000 419.510000 1.100000 ;
      RECT 412.090000 0.000000 415.350000 1.100000 ;
      RECT 407.935000 0.000000 411.190000 1.100000 ;
      RECT 403.775000 0.000000 407.035000 1.100000 ;
      RECT 399.620000 0.000000 402.875000 1.100000 ;
      RECT 395.460000 0.000000 398.720000 1.100000 ;
      RECT 391.300000 0.000000 394.560000 1.100000 ;
      RECT 387.145000 0.000000 390.400000 1.100000 ;
      RECT 382.985000 0.000000 386.245000 1.100000 ;
      RECT 378.830000 0.000000 382.085000 1.100000 ;
      RECT 374.670000 0.000000 377.930000 1.100000 ;
      RECT 370.510000 0.000000 373.770000 1.100000 ;
      RECT 366.355000 0.000000 369.610000 1.100000 ;
      RECT 362.195000 0.000000 365.455000 1.100000 ;
      RECT 358.040000 0.000000 361.295000 1.100000 ;
      RECT 353.880000 0.000000 357.140000 1.100000 ;
      RECT 349.720000 0.000000 352.980000 1.100000 ;
      RECT 345.565000 0.000000 348.820000 1.100000 ;
      RECT 341.405000 0.000000 344.665000 1.100000 ;
      RECT 337.250000 0.000000 340.505000 1.100000 ;
      RECT 333.090000 0.000000 336.350000 1.100000 ;
      RECT 328.930000 0.000000 332.190000 1.100000 ;
      RECT 324.775000 0.000000 328.030000 1.100000 ;
      RECT 320.615000 0.000000 323.875000 1.100000 ;
      RECT 316.460000 0.000000 319.715000 1.100000 ;
      RECT 312.300000 0.000000 315.560000 1.100000 ;
      RECT 308.140000 0.000000 311.400000 1.100000 ;
      RECT 303.985000 0.000000 307.240000 1.100000 ;
      RECT 299.825000 0.000000 303.085000 1.100000 ;
      RECT 295.670000 0.000000 298.925000 1.100000 ;
      RECT 291.510000 0.000000 294.770000 1.100000 ;
      RECT 287.350000 0.000000 290.610000 1.100000 ;
      RECT 283.195000 0.000000 286.450000 1.100000 ;
      RECT 279.035000 0.000000 282.295000 1.100000 ;
      RECT 274.880000 0.000000 278.135000 1.100000 ;
      RECT 270.720000 0.000000 273.980000 1.100000 ;
      RECT 266.560000 0.000000 269.820000 1.100000 ;
      RECT 262.405000 0.000000 265.660000 1.100000 ;
      RECT 258.245000 0.000000 261.505000 1.100000 ;
      RECT 254.090000 0.000000 257.345000 1.100000 ;
      RECT 249.930000 0.000000 253.190000 1.100000 ;
      RECT 245.770000 0.000000 249.030000 1.100000 ;
      RECT 241.615000 0.000000 244.870000 1.100000 ;
      RECT 237.455000 0.000000 240.715000 1.100000 ;
      RECT 233.300000 0.000000 236.555000 1.100000 ;
      RECT 229.140000 0.000000 232.400000 1.100000 ;
      RECT 224.980000 0.000000 228.240000 1.100000 ;
      RECT 220.825000 0.000000 224.080000 1.100000 ;
      RECT 216.665000 0.000000 219.925000 1.100000 ;
      RECT 212.510000 0.000000 215.765000 1.100000 ;
      RECT 208.350000 0.000000 211.610000 1.100000 ;
      RECT 204.190000 0.000000 207.450000 1.100000 ;
      RECT 200.035000 0.000000 203.290000 1.100000 ;
      RECT 195.875000 0.000000 199.135000 1.100000 ;
      RECT 191.720000 0.000000 194.975000 1.100000 ;
      RECT 187.560000 0.000000 190.820000 1.100000 ;
      RECT 183.400000 0.000000 186.660000 1.100000 ;
      RECT 179.245000 0.000000 182.500000 1.100000 ;
      RECT 175.085000 0.000000 178.345000 1.100000 ;
      RECT 170.930000 0.000000 174.185000 1.100000 ;
      RECT 166.770000 0.000000 170.030000 1.100000 ;
      RECT 162.610000 0.000000 165.870000 1.100000 ;
      RECT 158.455000 0.000000 161.710000 1.100000 ;
      RECT 154.295000 0.000000 157.555000 1.100000 ;
      RECT 150.140000 0.000000 153.395000 1.100000 ;
      RECT 145.980000 0.000000 149.240000 1.100000 ;
      RECT 141.820000 0.000000 145.080000 1.100000 ;
      RECT 137.665000 0.000000 140.920000 1.100000 ;
      RECT 133.505000 0.000000 136.765000 1.100000 ;
      RECT 129.350000 0.000000 132.605000 1.100000 ;
      RECT 125.190000 0.000000 128.450000 1.100000 ;
      RECT 121.030000 0.000000 124.290000 1.100000 ;
      RECT 116.875000 0.000000 120.130000 1.100000 ;
      RECT 112.715000 0.000000 115.975000 1.100000 ;
      RECT 108.560000 0.000000 111.815000 1.100000 ;
      RECT 104.400000 0.000000 107.660000 1.100000 ;
      RECT 100.240000 0.000000 103.500000 1.100000 ;
      RECT 96.085000 0.000000 99.340000 1.100000 ;
      RECT 91.925000 0.000000 95.185000 1.100000 ;
      RECT 87.770000 0.000000 91.025000 1.100000 ;
      RECT 83.610000 0.000000 86.870000 1.100000 ;
      RECT 79.450000 0.000000 82.710000 1.100000 ;
      RECT 75.295000 0.000000 78.550000 1.100000 ;
      RECT 71.135000 0.000000 74.395000 1.100000 ;
      RECT 66.980000 0.000000 70.235000 1.100000 ;
      RECT 62.820000 0.000000 66.080000 1.100000 ;
      RECT 58.660000 0.000000 61.920000 1.100000 ;
      RECT 54.505000 0.000000 57.760000 1.100000 ;
      RECT 50.345000 0.000000 53.605000 1.100000 ;
      RECT 46.190000 0.000000 49.445000 1.100000 ;
      RECT 42.030000 0.000000 45.290000 1.100000 ;
      RECT 37.870000 0.000000 41.130000 1.100000 ;
      RECT 33.715000 0.000000 36.970000 1.100000 ;
      RECT 29.555000 0.000000 32.815000 1.100000 ;
      RECT 25.400000 0.000000 28.655000 1.100000 ;
      RECT 21.240000 0.000000 24.500000 1.100000 ;
      RECT 17.080000 0.000000 20.340000 1.100000 ;
      RECT 12.925000 0.000000 16.180000 1.100000 ;
      RECT 8.765000 0.000000 12.025000 1.100000 ;
      RECT 4.610000 0.000000 7.865000 1.100000 ;
      RECT 2.060000 0.000000 3.710000 1.100000 ;
      RECT 0.000000 0.000000 1.160000 1.100000 ;
    LAYER met4 ;
      RECT 0.000000 1945.840000 2050.220000 1949.900000 ;
      RECT 5.020000 1945.820000 2038.000000 1945.840000 ;
      RECT 2040.400000 1942.240000 2045.200000 1945.840000 ;
      RECT 15.820000 1942.240000 2038.000000 1945.820000 ;
      RECT 5.020000 1942.240000 13.420000 1945.820000 ;
      RECT 15.820000 1933.895000 2034.400000 1942.240000 ;
      RECT 19.170000 1930.295000 2029.450000 1933.895000 ;
      RECT 2028.250000 22.575000 2029.450000 1930.295000 ;
      RECT 22.770000 22.575000 2025.850000 1930.295000 ;
      RECT 19.170000 22.575000 20.370000 1930.295000 ;
      RECT 2031.850000 18.975000 2034.400000 1933.895000 ;
      RECT 19.170000 18.975000 2029.450000 22.575000 ;
      RECT 15.820000 18.975000 16.770000 1933.895000 ;
      RECT 2044.000000 5.960000 2045.200000 1942.240000 ;
      RECT 2040.400000 5.960000 2041.600000 1942.240000 ;
      RECT 2036.800000 5.960000 2038.000000 1942.240000 ;
      RECT 15.820000 5.960000 2034.400000 18.975000 ;
      RECT 12.220000 5.960000 13.420000 1942.240000 ;
      RECT 8.620000 5.960000 9.820000 1942.240000 ;
      RECT 5.020000 5.960000 6.220000 1942.240000 ;
      RECT 2047.600000 2.360000 2050.220000 1945.840000 ;
      RECT 2040.400000 2.360000 2045.200000 5.960000 ;
      RECT 15.820000 2.360000 2038.000000 5.960000 ;
      RECT 5.020000 2.360000 13.420000 5.960000 ;
      RECT 0.000000 2.360000 2.620000 1945.840000 ;
      RECT 0.000000 0.000000 2050.220000 2.360000 ;
    LAYER met5 ;
      RECT 0.000000 0.000000 2050.220000 1949.900000 ;
  END
END azadi_soc_top_caravel

END LIBRARY
