##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Fri Jun  3 13:54:56 2022
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO azadi_soc_top_caravel
  CLASS BLOCK ;
  SIZE 2029.980000 BY 1929.840000 ;
  FOREIGN azadi_soc_top_caravel 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1853 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.792 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 428.340000 0.000000 428.640000 0.800000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.0724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met3  ;
    ANTENNAMAXAREACAR 10.1697 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 51.5131 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.0923232 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1927.240000 0.800000 1927.540000 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 4.220000 0.000000 4.520000 0.800000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 288.500000 0.000000 288.800000 0.800000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.460000 0.000000 1.760000 0.800000 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 8.360000 0.000000 8.660000 0.800000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 12.500000 0.000000 12.800000 0.800000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 16.640000 0.000000 16.940000 0.800000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 20.780000 0.000000 21.080000 0.800000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.940000 0.000000 157.240000 0.800000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.080000 0.000000 161.380000 0.800000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 164.760000 0.000000 165.060000 0.800000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 168.900000 0.000000 169.200000 0.800000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 173.040000 0.000000 173.340000 0.800000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 177.180000 0.000000 177.480000 0.800000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 181.320000 0.000000 181.620000 0.800000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 185.460000 0.000000 185.760000 0.800000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 189.600000 0.000000 189.900000 0.800000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 193.740000 0.000000 194.040000 0.800000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 197.880000 0.000000 198.180000 0.800000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 202.020000 0.000000 202.320000 0.800000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.160000 0.000000 206.460000 0.800000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.300000 0.000000 210.600000 0.800000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.440000 0.000000 214.740000 0.800000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.580000 0.000000 218.880000 0.800000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 222.720000 0.000000 223.020000 0.800000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 226.860000 0.000000 227.160000 0.800000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 231.000000 0.000000 231.300000 0.800000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 235.140000 0.000000 235.440000 0.800000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.280000 0.000000 239.580000 0.800000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 243.420000 0.000000 243.720000 0.800000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 247.100000 0.000000 247.400000 0.800000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 251.240000 0.000000 251.540000 0.800000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 255.380000 0.000000 255.680000 0.800000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 259.520000 0.000000 259.820000 0.800000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 263.660000 0.000000 263.960000 0.800000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 267.800000 0.000000 268.100000 0.800000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 271.940000 0.000000 272.240000 0.800000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 276.080000 0.000000 276.380000 0.800000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 280.220000 0.000000 280.520000 0.800000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 284.360000 0.000000 284.660000 0.800000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 292.640000 0.000000 292.940000 0.800000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.780000 0.000000 297.080000 0.800000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 300.920000 0.000000 301.220000 0.800000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 305.060000 0.000000 305.360000 0.800000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 309.200000 0.000000 309.500000 0.800000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.340000 0.000000 313.640000 0.800000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 317.480000 0.000000 317.780000 0.800000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 321.620000 0.000000 321.920000 0.800000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 325.300000 0.000000 325.600000 0.800000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 329.440000 0.000000 329.740000 0.800000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 333.580000 0.000000 333.880000 0.800000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 337.720000 0.000000 338.020000 0.800000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 341.860000 0.000000 342.160000 0.800000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000000 0.000000 346.300000 0.800000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 350.140000 0.000000 350.440000 0.800000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 354.280000 0.000000 354.580000 0.800000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 358.420000 0.000000 358.720000 0.800000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 362.560000 0.000000 362.860000 0.800000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.700000 0.000000 367.000000 0.800000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 370.840000 0.000000 371.140000 0.800000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 374.980000 0.000000 375.280000 0.800000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 379.120000 0.000000 379.420000 0.800000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.260000 0.000000 383.560000 0.800000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 387.400000 0.000000 387.700000 0.800000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 391.540000 0.000000 391.840000 0.800000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.680000 0.000000 395.980000 0.800000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 399.820000 0.000000 400.120000 0.800000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 403.960000 0.000000 404.260000 0.800000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 407.640000 0.000000 407.940000 0.800000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 411.780000 0.000000 412.080000 0.800000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 415.920000 0.000000 416.220000 0.800000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 420.060000 0.000000 420.360000 0.800000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.748 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 549.88 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 424.200000 0.000000 424.500000 0.800000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.748 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 549.88 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 24.920000 0.000000 25.220000 0.800000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.296 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.060000 0.000000 29.360000 0.800000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.296 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 33.200000 0.000000 33.500000 0.800000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.296 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 37.340000 0.000000 37.640000 0.800000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.488 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 41.480000 0.000000 41.780000 0.800000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.748 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 549.88 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 45.620000 0.000000 45.920000 0.800000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 49.760000 0.000000 50.060000 0.800000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 53.900000 0.000000 54.200000 0.800000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 58.040000 0.000000 58.340000 0.800000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 62.180000 0.000000 62.480000 0.800000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 66.320000 0.000000 66.620000 0.800000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 70.460000 0.000000 70.760000 0.800000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 74.600000 0.000000 74.900000 0.800000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 78.740000 0.000000 79.040000 0.800000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 82.420000 0.000000 82.720000 0.800000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 86.560000 0.000000 86.860000 0.800000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 90.700000 0.000000 91.000000 0.800000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 94.840000 0.000000 95.140000 0.800000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 98.980000 0.000000 99.280000 0.800000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 103.120000 0.000000 103.420000 0.800000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 107.260000 0.000000 107.560000 0.800000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 111.400000 0.000000 111.700000 0.800000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 115.540000 0.000000 115.840000 0.800000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 119.680000 0.000000 119.980000 0.800000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 123.820000 0.000000 124.120000 0.800000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 127.960000 0.000000 128.260000 0.800000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 132.100000 0.000000 132.400000 0.800000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 136.240000 0.000000 136.540000 0.800000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 140.380000 0.000000 140.680000 0.800000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 144.520000 0.000000 144.820000 0.800000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 148.660000 0.000000 148.960000 0.800000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.296 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 152.800000 0.000000 153.100000 0.800000 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1502.900000 0.000000 1503.200000 0.800000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1507.040000 0.000000 1507.340000 0.800000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1511.180000 0.000000 1511.480000 0.800000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1515.320000 0.000000 1515.620000 0.800000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1519.460000 0.000000 1519.760000 0.800000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1523.600000 0.000000 1523.900000 0.800000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1527.740000 0.000000 1528.040000 0.800000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1531.880000 0.000000 1532.180000 0.800000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1536.020000 0.000000 1536.320000 0.800000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1540.160000 0.000000 1540.460000 0.800000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1543.840000 0.000000 1544.140000 0.800000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1547.980000 0.000000 1548.280000 0.800000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1552.120000 0.000000 1552.420000 0.800000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1556.260000 0.000000 1556.560000 0.800000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1560.400000 0.000000 1560.700000 0.800000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1564.540000 0.000000 1564.840000 0.800000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1568.680000 0.000000 1568.980000 0.800000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1572.820000 0.000000 1573.120000 0.800000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1576.960000 0.000000 1577.260000 0.800000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.100000 0.000000 1581.400000 0.800000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1585.240000 0.000000 1585.540000 0.800000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1589.380000 0.000000 1589.680000 0.800000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1593.520000 0.000000 1593.820000 0.800000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1597.660000 0.000000 1597.960000 0.800000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1601.800000 0.000000 1602.100000 0.800000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1605.940000 0.000000 1606.240000 0.800000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1610.080000 0.000000 1610.380000 0.800000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1614.220000 0.000000 1614.520000 0.800000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1618.360000 0.000000 1618.660000 0.800000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1622.500000 0.000000 1622.800000 0.800000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1626.180000 0.000000 1626.480000 0.800000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1630.320000 0.000000 1630.620000 0.800000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1634.460000 0.000000 1634.760000 0.800000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1638.600000 0.000000 1638.900000 0.800000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1642.740000 0.000000 1643.040000 0.800000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1646.880000 0.000000 1647.180000 0.800000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1651.020000 0.000000 1651.320000 0.800000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1655.160000 0.000000 1655.460000 0.800000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1659.300000 0.000000 1659.600000 0.800000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1663.440000 0.000000 1663.740000 0.800000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1667.580000 0.000000 1667.880000 0.800000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1671.720000 0.000000 1672.020000 0.800000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1675.860000 0.000000 1676.160000 0.800000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1680.000000 0.000000 1680.300000 0.800000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1684.140000 0.000000 1684.440000 0.800000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1688.280000 0.000000 1688.580000 0.800000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1692.420000 0.000000 1692.720000 0.800000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.560000 0.000000 1696.860000 0.800000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1700.700000 0.000000 1701.000000 0.800000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1704.840000 0.000000 1705.140000 0.800000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1708.520000 0.000000 1708.820000 0.800000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1712.660000 0.000000 1712.960000 0.800000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1716.800000 0.000000 1717.100000 0.800000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1720.940000 0.000000 1721.240000 0.800000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1725.080000 0.000000 1725.380000 0.800000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1729.220000 0.000000 1729.520000 0.800000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1733.360000 0.000000 1733.660000 0.800000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1737.500000 0.000000 1737.800000 0.800000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.640000 0.000000 1741.940000 0.800000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1745.780000 0.000000 1746.080000 0.800000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1749.920000 0.000000 1750.220000 0.800000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1754.060000 0.000000 1754.360000 0.800000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1758.200000 0.000000 1758.500000 0.800000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1762.340000 0.000000 1762.640000 0.800000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1766.480000 0.000000 1766.780000 0.800000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1770.620000 0.000000 1770.920000 0.800000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1774.760000 0.000000 1775.060000 0.800000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1778.900000 0.000000 1779.200000 0.800000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1783.040000 0.000000 1783.340000 0.800000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1786.720000 0.000000 1787.020000 0.800000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1790.860000 0.000000 1791.160000 0.800000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1795.000000 0.000000 1795.300000 0.800000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1799.140000 0.000000 1799.440000 0.800000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1803.280000 0.000000 1803.580000 0.800000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1807.420000 0.000000 1807.720000 0.800000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1811.560000 0.000000 1811.860000 0.800000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1815.700000 0.000000 1816.000000 0.800000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1819.840000 0.000000 1820.140000 0.800000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1823.980000 0.000000 1824.280000 0.800000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1828.120000 0.000000 1828.420000 0.800000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1832.260000 0.000000 1832.560000 0.800000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1836.400000 0.000000 1836.700000 0.800000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1840.540000 0.000000 1840.840000 0.800000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1844.680000 0.000000 1844.980000 0.800000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1848.820000 0.000000 1849.120000 0.800000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1852.960000 0.000000 1853.260000 0.800000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1857.100000 0.000000 1857.400000 0.800000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1861.240000 0.000000 1861.540000 0.800000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1865.380000 0.000000 1865.680000 0.800000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1869.060000 0.000000 1869.360000 0.800000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1873.200000 0.000000 1873.500000 0.800000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1877.340000 0.000000 1877.640000 0.800000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1881.480000 0.000000 1881.780000 0.800000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1885.620000 0.000000 1885.920000 0.800000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1889.760000 0.000000 1890.060000 0.800000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1893.900000 0.000000 1894.200000 0.800000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1898.040000 0.000000 1898.340000 0.800000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1902.180000 0.000000 1902.480000 0.800000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1906.320000 0.000000 1906.620000 0.800000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1910.460000 0.000000 1910.760000 0.800000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1914.600000 0.000000 1914.900000 0.800000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1918.740000 0.000000 1919.040000 0.800000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1922.880000 0.000000 1923.180000 0.800000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1927.020000 0.000000 1927.320000 0.800000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1931.160000 0.000000 1931.460000 0.800000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1935.300000 0.000000 1935.600000 0.800000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1939.440000 0.000000 1939.740000 0.800000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1943.580000 0.000000 1943.880000 0.800000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1947.720000 0.000000 1948.020000 0.800000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1951.400000 0.000000 1951.700000 0.800000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1955.540000 0.000000 1955.840000 0.800000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1959.680000 0.000000 1959.980000 0.800000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 29.2701 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 157.048 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1963.820000 0.000000 1964.120000 0.800000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.2001 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 146.008 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1967.960000 0.000000 1968.260000 0.800000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.6601 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 127.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1972.100000 0.000000 1972.400000 0.800000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.4341 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 99.256 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1976.240000 0.000000 1976.540000 0.800000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.8621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 170.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1980.380000 0.000000 1980.680000 0.800000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.1641 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 129.816 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1984.520000 0.000000 1984.820000 0.800000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7241 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 170.136 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1988.660000 0.000000 1988.960000 0.800000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 29.6541 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 159.096 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1992.800000 0.000000 1993.100000 0.800000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.3761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 136.28 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1996.940000 0.000000 1997.240000 0.800000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.0181 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123.704 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2001.080000 0.000000 2001.380000 0.800000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9856 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.248 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.3148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.816 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2005.220000 0.000000 2005.520000 0.800000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 113.376 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 605.144 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2009.360000 0.000000 2009.660000 0.800000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9856 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.248 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.0468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.72 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2013.500000 0.000000 2013.800000 0.800000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9856 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.248 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.9618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2017.640000 0.000000 2017.940000 0.800000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 30.6501 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 164.408 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2021.780000 0.000000 2022.080000 0.800000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.7993 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.4 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2025.920000 0.000000 2026.220000 0.800000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.296 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 975.740000 0.000000 976.040000 0.800000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 979.880000 0.000000 980.180000 0.800000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 984.020000 0.000000 984.320000 0.800000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 988.160000 0.000000 988.460000 0.800000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 992.300000 0.000000 992.600000 0.800000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.296 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 996.440000 0.000000 996.740000 0.800000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1000.580000 0.000000 1000.880000 0.800000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1004.720000 0.000000 1005.020000 0.800000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1008.860000 0.000000 1009.160000 0.800000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1013.000000 0.000000 1013.300000 0.800000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1017.140000 0.000000 1017.440000 0.800000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1021.280000 0.000000 1021.580000 0.800000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1025.420000 0.000000 1025.720000 0.800000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1029.560000 0.000000 1029.860000 0.800000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1033.700000 0.000000 1034.000000 0.800000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.296 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1037.840000 0.000000 1038.140000 0.800000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.296 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1041.980000 0.000000 1042.280000 0.800000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1046.120000 0.000000 1046.420000 0.800000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1050.260000 0.000000 1050.560000 0.800000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1054.400000 0.000000 1054.700000 0.800000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1058.080000 0.000000 1058.380000 0.800000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.296 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1062.220000 0.000000 1062.520000 0.800000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.296 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1066.360000 0.000000 1066.660000 0.800000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1070.500000 0.000000 1070.800000 0.800000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1074.640000 0.000000 1074.940000 0.800000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1078.780000 0.000000 1079.080000 0.800000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1082.920000 0.000000 1083.220000 0.800000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1087.060000 0.000000 1087.360000 0.800000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1091.200000 0.000000 1091.500000 0.800000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1095.340000 0.000000 1095.640000 0.800000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1099.480000 0.000000 1099.780000 0.800000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1103.620000 0.000000 1103.920000 0.800000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1107.760000 0.000000 1108.060000 0.800000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1111.900000 0.000000 1112.200000 0.800000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1116.040000 0.000000 1116.340000 0.800000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.296 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1120.180000 0.000000 1120.480000 0.800000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.488 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1124.320000 0.000000 1124.620000 0.800000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.488 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1128.460000 0.000000 1128.760000 0.800000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.748 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 549.88 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1132.600000 0.000000 1132.900000 0.800000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.416 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2560.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1136.740000 0.000000 1137.040000 0.800000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.416 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2560.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1140.420000 0.000000 1140.720000 0.800000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.416 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2560.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1144.560000 0.000000 1144.860000 0.800000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.416 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2560.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1148.700000 0.000000 1149.000000 0.800000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.416 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2560.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1152.840000 0.000000 1153.140000 0.800000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.416 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2560.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1156.980000 0.000000 1157.280000 0.800000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.416 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2560.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1161.120000 0.000000 1161.420000 0.800000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1165.260000 0.000000 1165.560000 0.800000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1169.400000 0.000000 1169.700000 0.800000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1173.540000 0.000000 1173.840000 0.800000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1177.680000 0.000000 1177.980000 0.800000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1181.820000 0.000000 1182.120000 0.800000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1185.960000 0.000000 1186.260000 0.800000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1190.100000 0.000000 1190.400000 0.800000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1194.240000 0.000000 1194.540000 0.800000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1198.380000 0.000000 1198.680000 0.800000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.416 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2560.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1202.520000 0.000000 1202.820000 0.800000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.416 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2560.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1206.660000 0.000000 1206.960000 0.800000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1210.800000 0.000000 1211.100000 0.800000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1214.940000 0.000000 1215.240000 0.800000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1218.620000 0.000000 1218.920000 0.800000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1222.760000 0.000000 1223.060000 0.800000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1226.900000 0.000000 1227.200000 0.800000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1231.040000 0.000000 1231.340000 0.800000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1235.180000 0.000000 1235.480000 0.800000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1239.320000 0.000000 1239.620000 0.800000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1243.460000 0.000000 1243.760000 0.800000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1247.600000 0.000000 1247.900000 0.800000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1251.740000 0.000000 1252.040000 0.800000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1255.880000 0.000000 1256.180000 0.800000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1260.020000 0.000000 1260.320000 0.800000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1264.160000 0.000000 1264.460000 0.800000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1268.300000 0.000000 1268.600000 0.800000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1272.440000 0.000000 1272.740000 0.800000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1276.580000 0.000000 1276.880000 0.800000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1280.720000 0.000000 1281.020000 0.800000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.416 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2560.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1284.860000 0.000000 1285.160000 0.800000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.416 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2560.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1289.000000 0.000000 1289.300000 0.800000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1293.140000 0.000000 1293.440000 0.800000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1297.280000 0.000000 1297.580000 0.800000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1300.960000 0.000000 1301.260000 0.800000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1305.100000 0.000000 1305.400000 0.800000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1309.240000 0.000000 1309.540000 0.800000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1313.380000 0.000000 1313.680000 0.800000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1317.520000 0.000000 1317.820000 0.800000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1321.660000 0.000000 1321.960000 0.800000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1325.800000 0.000000 1326.100000 0.800000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1329.940000 0.000000 1330.240000 0.800000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1334.080000 0.000000 1334.380000 0.800000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1338.220000 0.000000 1338.520000 0.800000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1342.360000 0.000000 1342.660000 0.800000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1346.500000 0.000000 1346.800000 0.800000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.416 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2560.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1350.640000 0.000000 1350.940000 0.800000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.416 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2560.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1354.780000 0.000000 1355.080000 0.800000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1358.920000 0.000000 1359.220000 0.800000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1363.060000 0.000000 1363.360000 0.800000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.416 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2560.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1367.200000 0.000000 1367.500000 0.800000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.416 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2560.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1371.340000 0.000000 1371.640000 0.800000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1375.480000 0.000000 1375.780000 0.800000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1379.620000 0.000000 1379.920000 0.800000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1383.300000 0.000000 1383.600000 0.800000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1387.440000 0.000000 1387.740000 0.800000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1391.580000 0.000000 1391.880000 0.800000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1395.720000 0.000000 1396.020000 0.800000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1399.860000 0.000000 1400.160000 0.800000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1404.000000 0.000000 1404.300000 0.800000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1408.140000 0.000000 1408.440000 0.800000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1412.280000 0.000000 1412.580000 0.800000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1416.420000 0.000000 1416.720000 0.800000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1420.560000 0.000000 1420.860000 0.800000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2559.81 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1424.700000 0.000000 1425.000000 0.800000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.416 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2560.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1428.840000 0.000000 1429.140000 0.800000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 490.692 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2610.53 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1432.980000 0.000000 1433.280000 0.800000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.099 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 545 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 479.339 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2558.69 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1437.120000 0.000000 1437.420000 0.800000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.6195 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123.176 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 132.131 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 668.321 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 293.471 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1566.08 LAYER met4  ;
    ANTENNAGATEAREA 0.6915 LAYER met4  ;
    ANTENNAMAXAREACAR 556.528 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2933.08 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1441.260000 0.000000 1441.560000 0.800000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.6195 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123.176 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 115.112 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 626.85 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 293.471 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1566.08 LAYER met4  ;
    ANTENNAGATEAREA 0.6915 LAYER met4  ;
    ANTENNAMAXAREACAR 539.509 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2891.61 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1445.400000 0.000000 1445.700000 0.800000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.6195 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123.176 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 115.112 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 626.85 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 293.471 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1566.08 LAYER met4  ;
    ANTENNAGATEAREA 0.6915 LAYER met4  ;
    ANTENNAMAXAREACAR 539.509 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2891.61 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1449.540000 0.000000 1449.840000 0.800000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.6195 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 115.112 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 625.954 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 293.471 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1566.08 LAYER met4  ;
    ANTENNAGATEAREA 0.6915 LAYER met4  ;
    ANTENNAMAXAREACAR 539.509 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2890.71 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1453.680000 0.000000 1453.980000 0.800000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.6195 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 115.112 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 625.954 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 293.471 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1566.08 LAYER met4  ;
    ANTENNAGATEAREA 0.6915 LAYER met4  ;
    ANTENNAMAXAREACAR 539.509 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2890.71 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1457.820000 0.000000 1458.120000 0.800000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.6195 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 115.112 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 625.954 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 293.471 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1566.08 LAYER met4  ;
    ANTENNAGATEAREA 0.6915 LAYER met4  ;
    ANTENNAMAXAREACAR 539.509 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2890.71 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1461.500000 0.000000 1461.800000 0.800000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.6195 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 115.112 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 625.954 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 293.471 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1566.08 LAYER met4  ;
    ANTENNAGATEAREA 0.6915 LAYER met4  ;
    ANTENNAMAXAREACAR 539.509 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2890.71 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1465.640000 0.000000 1465.940000 0.800000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.6195 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 115.112 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 625.954 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 293.471 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1566.08 LAYER met4  ;
    ANTENNAGATEAREA 0.6915 LAYER met4  ;
    ANTENNAMAXAREACAR 539.509 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2890.71 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1469.780000 0.000000 1470.080000 0.800000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.6195 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 115.112 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 625.954 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 293.471 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1566.08 LAYER met4  ;
    ANTENNAGATEAREA 0.6915 LAYER met4  ;
    ANTENNAMAXAREACAR 539.509 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2890.71 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1473.920000 0.000000 1474.220000 0.800000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.6195 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 115.112 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 625.954 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 293.471 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1566.08 LAYER met4  ;
    ANTENNAGATEAREA 0.6915 LAYER met4  ;
    ANTENNAMAXAREACAR 539.509 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2890.71 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1478.060000 0.000000 1478.360000 0.800000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.6195 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 115.112 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 625.954 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 293.471 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1566.08 LAYER met4  ;
    ANTENNAGATEAREA 0.6915 LAYER met4  ;
    ANTENNAMAXAREACAR 539.509 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2890.71 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1482.200000 0.000000 1482.500000 0.800000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.6195 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123.176 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 115.112 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 626.85 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 293.471 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1566.08 LAYER met4  ;
    ANTENNAGATEAREA 0.6915 LAYER met4  ;
    ANTENNAMAXAREACAR 539.509 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2891.61 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1486.340000 0.000000 1486.640000 0.800000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.5745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 122.76 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 114.883 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 624.733 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 293.471 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1566.08 LAYER met4  ;
    ANTENNAGATEAREA 0.6915 LAYER met4  ;
    ANTENNAMAXAREACAR 539.28 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2889.49 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1490.480000 0.000000 1490.780000 0.800000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.6195 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123.368 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 115.112 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 627.827 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 293.471 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1566.08 LAYER met4  ;
    ANTENNAGATEAREA 0.6915 LAYER met4  ;
    ANTENNAMAXAREACAR 539.509 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2892.58 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1494.620000 0.000000 1494.920000 0.800000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.5745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 122.76 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 114.883 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 624.733 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 293.471 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1566.08 LAYER met4  ;
    ANTENNAGATEAREA 0.6915 LAYER met4  ;
    ANTENNAMAXAREACAR 539.28 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2889.49 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1498.760000 0.000000 1499.060000 0.800000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 449.040000 0.000000 449.340000 0.800000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 453.180000 0.000000 453.480000 0.800000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 457.320000 0.000000 457.620000 0.800000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.460000 0.000000 461.760000 0.800000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 465.600000 0.000000 465.900000 0.800000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 469.740000 0.000000 470.040000 0.800000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 473.880000 0.000000 474.180000 0.800000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 478.020000 0.000000 478.320000 0.800000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 482.160000 0.000000 482.460000 0.800000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 486.300000 0.000000 486.600000 0.800000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 489.980000 0.000000 490.280000 0.800000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 494.120000 0.000000 494.420000 0.800000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 498.260000 0.000000 498.560000 0.800000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 502.400000 0.000000 502.700000 0.800000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 506.540000 0.000000 506.840000 0.800000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 510.680000 0.000000 510.980000 0.800000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 514.820000 0.000000 515.120000 0.800000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 518.960000 0.000000 519.260000 0.800000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 523.100000 0.000000 523.400000 0.800000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 527.240000 0.000000 527.540000 0.800000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 531.380000 0.000000 531.680000 0.800000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 535.520000 0.000000 535.820000 0.800000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 539.660000 0.000000 539.960000 0.800000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 543.800000 0.000000 544.100000 0.800000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 547.940000 0.000000 548.240000 0.800000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 552.080000 0.000000 552.380000 0.800000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 556.220000 0.000000 556.520000 0.800000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 560.360000 0.000000 560.660000 0.800000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 564.500000 0.000000 564.800000 0.800000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 568.640000 0.000000 568.940000 0.800000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 572.320000 0.000000 572.620000 0.800000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 576.460000 0.000000 576.760000 0.800000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 580.600000 0.000000 580.900000 0.800000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 584.740000 0.000000 585.040000 0.800000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 588.880000 0.000000 589.180000 0.800000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 593.020000 0.000000 593.320000 0.800000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 597.160000 0.000000 597.460000 0.800000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 601.300000 0.000000 601.600000 0.800000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 605.440000 0.000000 605.740000 0.800000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 609.580000 0.000000 609.880000 0.800000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.720000 0.000000 614.020000 0.800000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 617.860000 0.000000 618.160000 0.800000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 622.000000 0.000000 622.300000 0.800000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 626.140000 0.000000 626.440000 0.800000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 630.280000 0.000000 630.580000 0.800000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 634.420000 0.000000 634.720000 0.800000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 638.560000 0.000000 638.860000 0.800000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 642.700000 0.000000 643.000000 0.800000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.840000 0.000000 647.140000 0.800000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 650.520000 0.000000 650.820000 0.800000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 654.660000 0.000000 654.960000 0.800000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 658.800000 0.000000 659.100000 0.800000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 662.940000 0.000000 663.240000 0.800000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 667.080000 0.000000 667.380000 0.800000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 671.220000 0.000000 671.520000 0.800000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 675.360000 0.000000 675.660000 0.800000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 679.500000 0.000000 679.800000 0.800000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 683.640000 0.000000 683.940000 0.800000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 687.780000 0.000000 688.080000 0.800000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 691.920000 0.000000 692.220000 0.800000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.060000 0.000000 696.360000 0.800000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 700.200000 0.000000 700.500000 0.800000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 704.340000 0.000000 704.640000 0.800000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 708.480000 0.000000 708.780000 0.800000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 712.620000 0.000000 712.920000 0.800000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 716.760000 0.000000 717.060000 0.800000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 720.900000 0.000000 721.200000 0.800000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 725.040000 0.000000 725.340000 0.800000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 729.180000 0.000000 729.480000 0.800000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 732.860000 0.000000 733.160000 0.800000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 737.000000 0.000000 737.300000 0.800000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 741.140000 0.000000 741.440000 0.800000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 745.280000 0.000000 745.580000 0.800000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 749.420000 0.000000 749.720000 0.800000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 753.560000 0.000000 753.860000 0.800000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 757.700000 0.000000 758.000000 0.800000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 761.840000 0.000000 762.140000 0.800000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 765.980000 0.000000 766.280000 0.800000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 770.120000 0.000000 770.420000 0.800000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 774.260000 0.000000 774.560000 0.800000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 778.400000 0.000000 778.700000 0.800000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 782.540000 0.000000 782.840000 0.800000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 786.680000 0.000000 786.980000 0.800000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 790.820000 0.000000 791.120000 0.800000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.960000 0.000000 795.260000 0.800000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 799.100000 0.000000 799.400000 0.800000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 803.240000 0.000000 803.540000 0.800000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 807.380000 0.000000 807.680000 0.800000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 811.520000 0.000000 811.820000 0.800000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 815.200000 0.000000 815.500000 0.800000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.340000 0.000000 819.640000 0.800000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 823.480000 0.000000 823.780000 0.800000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 827.620000 0.000000 827.920000 0.800000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 831.760000 0.000000 832.060000 0.800000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.900000 0.000000 836.200000 0.800000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 840.040000 0.000000 840.340000 0.800000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 844.180000 0.000000 844.480000 0.800000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 848.320000 0.000000 848.620000 0.800000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 852.460000 0.000000 852.760000 0.800000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 856.600000 0.000000 856.900000 0.800000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 860.740000 0.000000 861.040000 0.800000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 864.880000 0.000000 865.180000 0.800000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 869.020000 0.000000 869.320000 0.800000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 873.160000 0.000000 873.460000 0.800000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 877.300000 0.000000 877.600000 0.800000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 881.440000 0.000000 881.740000 0.800000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 885.580000 0.000000 885.880000 0.800000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 889.720000 0.000000 890.020000 0.800000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 893.400000 0.000000 893.700000 0.800000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 897.540000 0.000000 897.840000 0.800000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 901.680000 0.000000 901.980000 0.800000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 905.820000 0.000000 906.120000 0.800000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 909.960000 0.000000 910.260000 0.800000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 914.100000 0.000000 914.400000 0.800000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 918.240000 0.000000 918.540000 0.800000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 922.380000 0.000000 922.680000 0.800000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 926.520000 0.000000 926.820000 0.800000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 930.660000 0.000000 930.960000 0.800000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 934.800000 0.000000 935.100000 0.800000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 938.940000 0.000000 939.240000 0.800000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 943.080000 0.000000 943.380000 0.800000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 947.220000 0.000000 947.520000 0.800000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 951.360000 0.000000 951.660000 0.800000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 955.500000 0.000000 955.800000 0.800000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 959.640000 0.000000 959.940000 0.800000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 963.780000 0.000000 964.080000 0.800000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 967.920000 0.000000 968.220000 0.800000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 972.060000 0.000000 972.360000 0.800000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 873.770000 0.800000 874.070000 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.2766 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 34.416 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 430.132 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2295.84 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 837.170000 0.800000 837.470000 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 176.598 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 942.776 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.7398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 800.570000 0.800000 800.870000 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.0112 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.6808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.768 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 764.580000 0.800000 764.880000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 543.484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2899.99 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 727.980000 0.800000 728.280000 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 691.380000 0.800000 691.680000 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 655.390000 0.800000 655.690000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 618.790000 0.800000 619.090000 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.7213 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.984 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 582.190000 0.800000 582.490000 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9673 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.296 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 546.200000 0.800000 546.500000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3253 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 509.600000 0.800000 509.900000 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.7213 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.984 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 473.000000 0.800000 473.300000 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.2803 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.632 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 437.010000 0.800000 437.310000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.7658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.888 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.562 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.4 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 400.410000 0.800000 400.710000 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.0131 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.344 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 985.400000 1929.040000 985.700000 1929.840000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.5361 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 115.8 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 927.440000 1929.040000 927.740000 1929.840000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.5673 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 131.496 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 869.480000 1929.040000 869.780000 1929.840000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.8341 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 128.056 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 811.520000 1929.040000 811.820000 1929.840000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.8073 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 148.776 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 753.560000 1929.040000 753.860000 1929.840000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 26.7321 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 143.512 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 695.600000 1929.040000 695.900000 1929.840000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.4503 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 130.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 637.640000 1929.040000 637.940000 1929.840000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2026 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.7608 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.528 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 579.680000 1929.040000 579.980000 1929.840000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 521.720000 1929.040000 522.020000 1929.840000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 1076.290000 2029.980000 1076.590000 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3713 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.784 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 1113.500000 2029.980000 1113.800000 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3713 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.784 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 1150.710000 2029.980000 1151.010000 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1466 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 134.45 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 717.536 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 1187.920000 2029.980000 1188.220000 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8633 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.408 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 1225.130000 2029.980000 1225.430000 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 1262.340000 2029.980000 1262.640000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 1298.940000 2029.980000 1299.240000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.2361 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 114.2 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 1336.150000 2029.980000 1336.450000 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 1373.360000 2029.980000 1373.660000 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7483 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 1410.570000 2029.980000 1410.870000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 1447.780000 2029.980000 1448.080000 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 1484.990000 2029.980000 1485.290000 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5543 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.76 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 1521.590000 2029.980000 1521.890000 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 1558.800000 2029.980000 1559.100000 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 1596.010000 2029.980000 1596.310000 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.47025 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.128 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 197.797 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1056.8 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1893.080000 0.800000 1893.380000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.6774 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.261 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 54.096 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1856.480000 0.800000 1856.780000 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 291.139 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1554.15 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1819.880000 0.800000 1820.180000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 606.711 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3236.26 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 198.746 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1060.45 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1783.890000 0.800000 1784.190000 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 310.305 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1655.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 179.849 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 959.664 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1747.290000 0.800000 1747.590000 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1403 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.552 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1710.690000 0.800000 1710.990000 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.36 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1674.700000 0.800000 1675.000000 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.7874 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 58.944 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.3174 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.136 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1638.100000 0.800000 1638.400000 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4686 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.101 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1073.01 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1601.500000 0.800000 1601.800000 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.4633 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.608 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1565.510000 0.800000 1565.810000 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1623 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.336 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1528.910000 0.800000 1529.210000 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.136 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1492.310000 0.800000 1492.610000 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6013 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.344 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1456.320000 0.800000 1456.620000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.3983 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 103.928 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1419.720000 0.800000 1420.020000 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 29.3935 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 157.696 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2019.940000 1929.040000 2020.240000 1929.840000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 28.8218 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 154.616 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1971.180000 1929.040000 1971.480000 1929.840000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.9233 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 138.728 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1913.220000 1929.040000 1913.520000 1929.840000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.2261 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 119.48 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1855.260000 1929.040000 1855.560000 1929.840000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2534 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.3258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.208 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1797.300000 1929.040000 1797.600000 1929.840000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 34.5813 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 184.904 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1739.340000 1929.040000 1739.640000 1929.840000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.3563 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.704 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1681.380000 1929.040000 1681.680000 1929.840000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.1194 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 124.224 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1623.420000 1929.040000 1623.720000 1929.840000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 134.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 719.112 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1565.460000 1929.040000 1565.760000 1929.840000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2003 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 4.520000 2029.980000 4.820000 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.5745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 122.76 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 114.883 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 624.733 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 293.471 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1566.08 LAYER met4  ;
    ANTENNAGATEAREA 0.6915 LAYER met4  ;
    ANTENNAMAXAREACAR 539.28 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2889.49 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 37.460000 2029.980000 37.760000 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.6195 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 115.112 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 625.954 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 293.471 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1566.08 LAYER met4  ;
    ANTENNAGATEAREA 0.6915 LAYER met4  ;
    ANTENNAMAXAREACAR 539.509 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2890.71 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 74.670000 2029.980000 74.970000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2116 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 293.471 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1566.08 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6915 LAYER met4  ;
    ANTENNAMAXAREACAR 424.397 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2264.76 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 111.880000 2029.980000 112.180000 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3946 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 293.471 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1566.08 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6915 LAYER met4  ;
    ANTENNAMAXAREACAR 424.397 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2264.76 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 149.090000 2029.980000 149.390000 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0963 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.984 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 186.300000 2029.980000 186.600000 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3353 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.592 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 222.900000 2029.980000 223.200000 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3946 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 293.471 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1566.08 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6915 LAYER met4  ;
    ANTENNAMAXAREACAR 424.397 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2264.76 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 260.110000 2029.980000 260.410000 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2333 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.048 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 297.320000 2029.980000 297.620000 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7756 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.128 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 293.471 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1566.08 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6915 LAYER met4  ;
    ANTENNAMAXAREACAR 424.397 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2264.76 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 334.530000 2029.980000 334.830000 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7035 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.752 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 371.740000 2029.980000 372.040000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5663 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.824 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 408.950000 2029.980000 409.250000 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0302 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 293.471 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1566.08 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6915 LAYER met4  ;
    ANTENNAMAXAREACAR 424.397 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2264.76 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 445.550000 2029.980000 445.850000 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 62.5458 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 334.048 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 482.760000 2029.980000 483.060000 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5293 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.96 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 519.970000 2029.980000 520.270000 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.5745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 122.76 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 114.883 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 624.733 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 293.471 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1566.08 LAYER met4  ;
    ANTENNAGATEAREA 0.6915 LAYER met4  ;
    ANTENNAMAXAREACAR 539.28 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2889.49 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2027.760000 0.000000 2028.060000 0.800000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.7184 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.16 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1383.120000 0.800000 1383.420000 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.6144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.272 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1347.130000 0.800000 1347.430000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.8994 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.792 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1310.530000 0.800000 1310.830000 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.9584 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.44 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1273.930000 0.800000 1274.230000 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4483 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 197.797 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1056.8 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1237.940000 0.800000 1238.240000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5503 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 197.797 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1056.8 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1201.340000 0.800000 1201.640000 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5503 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 197.797 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1056.8 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1164.740000 0.800000 1165.040000 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.0144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.072 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1128.750000 0.800000 1129.050000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.8904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.744 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1092.150000 0.800000 1092.450000 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.5194 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.432 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1055.550000 0.800000 1055.850000 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.4284 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.28 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1019.560000 0.800000 1019.860000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.0624 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 982.960000 0.800000 983.260000 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3804 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.024 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 946.360000 0.800000 946.660000 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8204 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.704 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 909.760000 0.800000 910.060000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3714 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.976 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1507.500000 1929.040000 1507.800000 1929.840000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.1884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1449.540000 1929.040000 1449.840000 1929.840000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.544 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1391.580000 1929.040000 1391.880000 1929.840000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.1764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.936 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1333.620000 1929.040000 1333.920000 1929.840000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.1764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.936 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1275.660000 1929.040000 1275.960000 1929.840000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.1764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.936 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1217.700000 1929.040000 1218.000000 1929.840000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.1764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.936 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1159.740000 1929.040000 1160.040000 1929.840000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.57765 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 197.797 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1056.8 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1101.780000 1929.040000 1102.080000 1929.840000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.97065 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 197.797 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1056.8 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1043.820000 1929.040000 1044.120000 1929.840000 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4773 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 557.180000 2029.980000 557.480000 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4773 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 594.390000 2029.980000 594.690000 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4773 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 631.600000 2029.980000 631.900000 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5523 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 668.200000 2029.980000 668.500000 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.0624 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 705.410000 2029.980000 705.710000 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.9924 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.288 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 742.620000 2029.980000 742.920000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4773 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 779.830000 2029.980000 780.130000 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3776 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 293.471 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1566.08 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6915 LAYER met4  ;
    ANTENNAMAXAREACAR 424.397 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2264.76 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 817.040000 2029.980000 817.340000 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4323 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 854.250000 2029.980000 854.550000 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3776 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 293.471 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1566.08 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6915 LAYER met4  ;
    ANTENNAMAXAREACAR 424.397 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2264.76 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 890.850000 2029.980000 891.150000 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3776 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 293.471 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1566.08 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6915 LAYER met4  ;
    ANTENNAMAXAREACAR 424.397 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2264.76 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 928.060000 2029.980000 928.360000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2116 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 965.270000 2029.980000 965.570000 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.5104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.384 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 1002.480000 2029.980000 1002.780000 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3005 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.736 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 7.79071 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 39.1495 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 293.471 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1566.08 LAYER met4  ;
    ANTENNAGATEAREA 0.6915 LAYER met4  ;
    ANTENNAMAXAREACAR 432.188 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2303.91 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 1039.690000 2029.980000 1039.990000 ;
    END
  END io_oeb[0]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 363.810000 0.800000 364.110000 ;
    END
  END analog_io[28]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 327.820000 0.800000 328.120000 ;
    END
  END analog_io[27]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 291.220000 0.800000 291.520000 ;
    END
  END analog_io[26]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 254.620000 0.800000 254.920000 ;
    END
  END analog_io[25]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 218.630000 0.800000 218.930000 ;
    END
  END analog_io[24]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 182.030000 0.800000 182.330000 ;
    END
  END analog_io[23]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 145.430000 0.800000 145.730000 ;
    END
  END analog_io[22]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 109.440000 0.800000 109.740000 ;
    END
  END analog_io[21]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 72.840000 0.800000 73.140000 ;
    END
  END analog_io[20]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 36.240000 0.800000 36.540000 ;
    END
  END analog_io[19]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 4.520000 0.800000 4.820000 ;
    END
  END analog_io[18]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 463.760000 1929.040000 464.060000 1929.840000 ;
    END
  END analog_io[17]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 405.800000 1929.040000 406.100000 1929.840000 ;
    END
  END analog_io[16]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 347.840000 1929.040000 348.140000 1929.840000 ;
    END
  END analog_io[15]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 289.880000 1929.040000 290.180000 1929.840000 ;
    END
  END analog_io[14]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 231.920000 1929.040000 232.220000 1929.840000 ;
    END
  END analog_io[13]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 173.960000 1929.040000 174.260000 1929.840000 ;
    END
  END analog_io[12]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000000 1929.040000 116.300000 1929.840000 ;
    END
  END analog_io[11]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 58.040000 1929.040000 58.340000 1929.840000 ;
    END
  END analog_io[10]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.460000 1929.040000 1.760000 1929.840000 ;
    END
  END analog_io[9]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 1633.220000 2029.980000 1633.520000 ;
    END
  END analog_io[8]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 1670.430000 2029.980000 1670.730000 ;
    END
  END analog_io[7]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 1707.640000 2029.980000 1707.940000 ;
    END
  END analog_io[6]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 1744.240000 2029.980000 1744.540000 ;
    END
  END analog_io[5]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 1781.450000 2029.980000 1781.750000 ;
    END
  END analog_io[4]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 1818.660000 2029.980000 1818.960000 ;
    END
  END analog_io[3]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 1855.870000 2029.980000 1856.170000 ;
    END
  END analog_io[2]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 1893.080000 2029.980000 1893.380000 ;
    END
  END analog_io[1]
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2029.180000 1926.020000 2029.980000 1926.320000 ;
    END
  END analog_io[0]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 444.900000 0.000000 445.200000 0.800000 ;
    END
  END user_clock2
  PIN user_irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.296 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 432.480000 0.000000 432.780000 0.800000 ;
    END
  END user_irq[2]
  PIN user_irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 436.620000 0.000000 436.920000 0.800000 ;
    END
  END user_irq[1]
  PIN user_irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 102.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 550.296 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 440.760000 0.000000 441.060000 0.800000 ;
    END
  END user_irq[0]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2023.760000 4.960000 2025.360000 1923.520000 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.620000 4.960000 6.220000 1923.520000 ;
    END

# P/G pin shape extracted from block 'azadi_soc_top'
    PORT
      LAYER met4 ;
        RECT 536.510000 76.020000 538.250000 464.000000 ;
      LAYER met4 ;
        RECT 67.990000 76.020000 69.730000 464.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 536.510000 1007.020000 538.250000 1395.000000 ;
      LAYER met4 ;
        RECT 67.990000 1007.020000 69.730000 1395.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 536.510000 1472.520000 538.250000 1860.500000 ;
      LAYER met4 ;
        RECT 67.990000 1472.520000 69.730000 1860.500000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1963.390000 70.480000 1965.130000 458.460000 ;
      LAYER met4 ;
        RECT 1494.870000 70.480000 1496.610000 458.460000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1963.390000 535.980000 1965.130000 923.960000 ;
      LAYER met4 ;
        RECT 1494.870000 535.980000 1496.610000 923.960000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1963.390000 1001.480000 1965.130000 1389.460000 ;
      LAYER met4 ;
        RECT 1494.870000 1001.480000 1496.610000 1389.460000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1963.390000 1466.980000 1965.130000 1854.960000 ;
      LAYER met4 ;
        RECT 1494.870000 1466.980000 1496.610000 1854.960000 ;
    END
    PORT
      LAYER met4 ;
        RECT 536.510000 541.520000 538.250000 929.500000 ;
      LAYER met4 ;
        RECT 67.990000 541.520000 69.730000 929.500000 ;
    END
    PORT
      LAYER met4 ;
        RECT 24.130000 20.975000 25.930000 1907.695000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2009.370000 20.975000 2011.170000 1907.695000 ;
    END
# end of P/G pin shape extracted from block 'azadi_soc_top'

  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2026.960000 1.760000 2028.560000 1926.720000 ;
    END

# P/G pin shape extracted from block 'azadi_soc_top'
    PORT
      LAYER met4 ;
        RECT 64.590000 72.620000 66.330000 467.400000 ;
      LAYER met4 ;
        RECT 539.910000 72.620000 541.650000 467.400000 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.590000 1003.620000 66.330000 1398.400000 ;
      LAYER met4 ;
        RECT 539.910000 1003.620000 541.650000 1398.400000 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.590000 1469.120000 66.330000 1863.900000 ;
      LAYER met4 ;
        RECT 539.910000 1469.120000 541.650000 1863.900000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1491.470000 67.080000 1493.210000 461.860000 ;
      LAYER met4 ;
        RECT 1966.790000 67.080000 1968.530000 461.860000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1491.470000 532.580000 1493.210000 927.360000 ;
      LAYER met4 ;
        RECT 1966.790000 532.580000 1968.530000 927.360000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1491.470000 998.080000 1493.210000 1392.860000 ;
      LAYER met4 ;
        RECT 1966.790000 998.080000 1968.530000 1392.860000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1491.470000 1463.580000 1493.210000 1858.360000 ;
      LAYER met4 ;
        RECT 1966.790000 1463.580000 1968.530000 1858.360000 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.590000 538.120000 66.330000 932.900000 ;
      LAYER met4 ;
        RECT 539.910000 538.120000 541.650000 932.900000 ;
    END
    PORT
      LAYER met4 ;
        RECT 20.530000 17.375000 22.330000 1911.295000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2012.970000 17.375000 2014.770000 1911.295000 ;
    END
# end of P/G pin shape extracted from block 'azadi_soc_top'

  END vssd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 2029.980000 1929.840000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 2029.980000 1929.840000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 2029.980000 1929.840000 ;
    LAYER met3 ;
      RECT 2020.540000 1928.740000 2029.980000 1929.840000 ;
      RECT 1971.780000 1928.740000 2019.640000 1929.840000 ;
      RECT 1913.820000 1928.740000 1970.880000 1929.840000 ;
      RECT 1855.860000 1928.740000 1912.920000 1929.840000 ;
      RECT 1797.900000 1928.740000 1854.960000 1929.840000 ;
      RECT 1739.940000 1928.740000 1797.000000 1929.840000 ;
      RECT 1681.980000 1928.740000 1739.040000 1929.840000 ;
      RECT 1624.020000 1928.740000 1681.080000 1929.840000 ;
      RECT 1566.060000 1928.740000 1623.120000 1929.840000 ;
      RECT 1508.100000 1928.740000 1565.160000 1929.840000 ;
      RECT 1450.140000 1928.740000 1507.200000 1929.840000 ;
      RECT 1392.180000 1928.740000 1449.240000 1929.840000 ;
      RECT 1334.220000 1928.740000 1391.280000 1929.840000 ;
      RECT 1276.260000 1928.740000 1333.320000 1929.840000 ;
      RECT 1218.300000 1928.740000 1275.360000 1929.840000 ;
      RECT 1160.340000 1928.740000 1217.400000 1929.840000 ;
      RECT 1102.380000 1928.740000 1159.440000 1929.840000 ;
      RECT 1044.420000 1928.740000 1101.480000 1929.840000 ;
      RECT 986.000000 1928.740000 1043.520000 1929.840000 ;
      RECT 928.040000 1928.740000 985.100000 1929.840000 ;
      RECT 870.080000 1928.740000 927.140000 1929.840000 ;
      RECT 812.120000 1928.740000 869.180000 1929.840000 ;
      RECT 754.160000 1928.740000 811.220000 1929.840000 ;
      RECT 696.200000 1928.740000 753.260000 1929.840000 ;
      RECT 638.240000 1928.740000 695.300000 1929.840000 ;
      RECT 580.280000 1928.740000 637.340000 1929.840000 ;
      RECT 522.320000 1928.740000 579.380000 1929.840000 ;
      RECT 464.360000 1928.740000 521.420000 1929.840000 ;
      RECT 406.400000 1928.740000 463.460000 1929.840000 ;
      RECT 348.440000 1928.740000 405.500000 1929.840000 ;
      RECT 290.480000 1928.740000 347.540000 1929.840000 ;
      RECT 232.520000 1928.740000 289.580000 1929.840000 ;
      RECT 174.560000 1928.740000 231.620000 1929.840000 ;
      RECT 116.600000 1928.740000 173.660000 1929.840000 ;
      RECT 58.640000 1928.740000 115.700000 1929.840000 ;
      RECT 2.060000 1928.740000 57.740000 1929.840000 ;
      RECT 0.000000 1928.740000 1.160000 1929.840000 ;
      RECT 0.000000 1927.840000 2029.980000 1928.740000 ;
      RECT 1.100000 1926.940000 2029.980000 1927.840000 ;
      RECT 0.000000 1926.620000 2029.980000 1926.940000 ;
      RECT 0.000000 1925.720000 2028.880000 1926.620000 ;
      RECT 0.000000 1893.680000 2029.980000 1925.720000 ;
      RECT 1.100000 1892.780000 2028.880000 1893.680000 ;
      RECT 0.000000 1857.080000 2029.980000 1892.780000 ;
      RECT 1.100000 1856.470000 2029.980000 1857.080000 ;
      RECT 1.100000 1856.180000 2028.880000 1856.470000 ;
      RECT 0.000000 1855.570000 2028.880000 1856.180000 ;
      RECT 0.000000 1820.480000 2029.980000 1855.570000 ;
      RECT 1.100000 1819.580000 2029.980000 1820.480000 ;
      RECT 0.000000 1819.260000 2029.980000 1819.580000 ;
      RECT 0.000000 1818.360000 2028.880000 1819.260000 ;
      RECT 0.000000 1784.490000 2029.980000 1818.360000 ;
      RECT 1.100000 1783.590000 2029.980000 1784.490000 ;
      RECT 0.000000 1782.050000 2029.980000 1783.590000 ;
      RECT 0.000000 1781.150000 2028.880000 1782.050000 ;
      RECT 0.000000 1747.890000 2029.980000 1781.150000 ;
      RECT 1.100000 1746.990000 2029.980000 1747.890000 ;
      RECT 0.000000 1744.840000 2029.980000 1746.990000 ;
      RECT 0.000000 1743.940000 2028.880000 1744.840000 ;
      RECT 0.000000 1711.290000 2029.980000 1743.940000 ;
      RECT 1.100000 1710.390000 2029.980000 1711.290000 ;
      RECT 0.000000 1708.240000 2029.980000 1710.390000 ;
      RECT 0.000000 1707.340000 2028.880000 1708.240000 ;
      RECT 0.000000 1675.300000 2029.980000 1707.340000 ;
      RECT 1.100000 1674.400000 2029.980000 1675.300000 ;
      RECT 0.000000 1671.030000 2029.980000 1674.400000 ;
      RECT 0.000000 1670.130000 2028.880000 1671.030000 ;
      RECT 0.000000 1638.700000 2029.980000 1670.130000 ;
      RECT 1.100000 1637.800000 2029.980000 1638.700000 ;
      RECT 0.000000 1633.820000 2029.980000 1637.800000 ;
      RECT 0.000000 1632.920000 2028.880000 1633.820000 ;
      RECT 0.000000 1602.100000 2029.980000 1632.920000 ;
      RECT 1.100000 1601.200000 2029.980000 1602.100000 ;
      RECT 0.000000 1596.610000 2029.980000 1601.200000 ;
      RECT 0.000000 1595.710000 2028.880000 1596.610000 ;
      RECT 0.000000 1566.110000 2029.980000 1595.710000 ;
      RECT 1.100000 1565.210000 2029.980000 1566.110000 ;
      RECT 0.000000 1559.400000 2029.980000 1565.210000 ;
      RECT 0.000000 1558.500000 2028.880000 1559.400000 ;
      RECT 0.000000 1529.510000 2029.980000 1558.500000 ;
      RECT 1.100000 1528.610000 2029.980000 1529.510000 ;
      RECT 0.000000 1522.190000 2029.980000 1528.610000 ;
      RECT 0.000000 1521.290000 2028.880000 1522.190000 ;
      RECT 0.000000 1492.910000 2029.980000 1521.290000 ;
      RECT 1.100000 1492.010000 2029.980000 1492.910000 ;
      RECT 0.000000 1485.590000 2029.980000 1492.010000 ;
      RECT 0.000000 1484.690000 2028.880000 1485.590000 ;
      RECT 0.000000 1456.920000 2029.980000 1484.690000 ;
      RECT 1.100000 1456.020000 2029.980000 1456.920000 ;
      RECT 0.000000 1448.380000 2029.980000 1456.020000 ;
      RECT 0.000000 1447.480000 2028.880000 1448.380000 ;
      RECT 0.000000 1420.320000 2029.980000 1447.480000 ;
      RECT 1.100000 1419.420000 2029.980000 1420.320000 ;
      RECT 0.000000 1411.170000 2029.980000 1419.420000 ;
      RECT 0.000000 1410.270000 2028.880000 1411.170000 ;
      RECT 0.000000 1383.720000 2029.980000 1410.270000 ;
      RECT 1.100000 1382.820000 2029.980000 1383.720000 ;
      RECT 0.000000 1373.960000 2029.980000 1382.820000 ;
      RECT 0.000000 1373.060000 2028.880000 1373.960000 ;
      RECT 0.000000 1347.730000 2029.980000 1373.060000 ;
      RECT 1.100000 1346.830000 2029.980000 1347.730000 ;
      RECT 0.000000 1336.750000 2029.980000 1346.830000 ;
      RECT 0.000000 1335.850000 2028.880000 1336.750000 ;
      RECT 0.000000 1311.130000 2029.980000 1335.850000 ;
      RECT 1.100000 1310.230000 2029.980000 1311.130000 ;
      RECT 0.000000 1299.540000 2029.980000 1310.230000 ;
      RECT 0.000000 1298.640000 2028.880000 1299.540000 ;
      RECT 0.000000 1274.530000 2029.980000 1298.640000 ;
      RECT 1.100000 1273.630000 2029.980000 1274.530000 ;
      RECT 0.000000 1262.940000 2029.980000 1273.630000 ;
      RECT 0.000000 1262.040000 2028.880000 1262.940000 ;
      RECT 0.000000 1238.540000 2029.980000 1262.040000 ;
      RECT 1.100000 1237.640000 2029.980000 1238.540000 ;
      RECT 0.000000 1225.730000 2029.980000 1237.640000 ;
      RECT 0.000000 1224.830000 2028.880000 1225.730000 ;
      RECT 0.000000 1201.940000 2029.980000 1224.830000 ;
      RECT 1.100000 1201.040000 2029.980000 1201.940000 ;
      RECT 0.000000 1188.520000 2029.980000 1201.040000 ;
      RECT 0.000000 1187.620000 2028.880000 1188.520000 ;
      RECT 0.000000 1165.340000 2029.980000 1187.620000 ;
      RECT 1.100000 1164.440000 2029.980000 1165.340000 ;
      RECT 0.000000 1151.310000 2029.980000 1164.440000 ;
      RECT 0.000000 1150.410000 2028.880000 1151.310000 ;
      RECT 0.000000 1129.350000 2029.980000 1150.410000 ;
      RECT 1.100000 1128.450000 2029.980000 1129.350000 ;
      RECT 0.000000 1114.100000 2029.980000 1128.450000 ;
      RECT 0.000000 1113.200000 2028.880000 1114.100000 ;
      RECT 0.000000 1092.750000 2029.980000 1113.200000 ;
      RECT 1.100000 1091.850000 2029.980000 1092.750000 ;
      RECT 0.000000 1076.890000 2029.980000 1091.850000 ;
      RECT 0.000000 1075.990000 2028.880000 1076.890000 ;
      RECT 0.000000 1056.150000 2029.980000 1075.990000 ;
      RECT 1.100000 1055.250000 2029.980000 1056.150000 ;
      RECT 0.000000 1040.290000 2029.980000 1055.250000 ;
      RECT 0.000000 1039.390000 2028.880000 1040.290000 ;
      RECT 0.000000 1020.160000 2029.980000 1039.390000 ;
      RECT 1.100000 1019.260000 2029.980000 1020.160000 ;
      RECT 0.000000 1003.080000 2029.980000 1019.260000 ;
      RECT 0.000000 1002.180000 2028.880000 1003.080000 ;
      RECT 0.000000 983.560000 2029.980000 1002.180000 ;
      RECT 1.100000 982.660000 2029.980000 983.560000 ;
      RECT 0.000000 965.870000 2029.980000 982.660000 ;
      RECT 0.000000 964.970000 2028.880000 965.870000 ;
      RECT 0.000000 946.960000 2029.980000 964.970000 ;
      RECT 1.100000 946.060000 2029.980000 946.960000 ;
      RECT 0.000000 928.660000 2029.980000 946.060000 ;
      RECT 0.000000 927.760000 2028.880000 928.660000 ;
      RECT 0.000000 910.360000 2029.980000 927.760000 ;
      RECT 1.100000 909.460000 2029.980000 910.360000 ;
      RECT 0.000000 891.450000 2029.980000 909.460000 ;
      RECT 0.000000 890.550000 2028.880000 891.450000 ;
      RECT 0.000000 874.370000 2029.980000 890.550000 ;
      RECT 1.100000 873.470000 2029.980000 874.370000 ;
      RECT 0.000000 854.850000 2029.980000 873.470000 ;
      RECT 0.000000 853.950000 2028.880000 854.850000 ;
      RECT 0.000000 837.770000 2029.980000 853.950000 ;
      RECT 1.100000 836.870000 2029.980000 837.770000 ;
      RECT 0.000000 817.640000 2029.980000 836.870000 ;
      RECT 0.000000 816.740000 2028.880000 817.640000 ;
      RECT 0.000000 801.170000 2029.980000 816.740000 ;
      RECT 1.100000 800.270000 2029.980000 801.170000 ;
      RECT 0.000000 780.430000 2029.980000 800.270000 ;
      RECT 0.000000 779.530000 2028.880000 780.430000 ;
      RECT 0.000000 765.180000 2029.980000 779.530000 ;
      RECT 1.100000 764.280000 2029.980000 765.180000 ;
      RECT 0.000000 743.220000 2029.980000 764.280000 ;
      RECT 0.000000 742.320000 2028.880000 743.220000 ;
      RECT 0.000000 728.580000 2029.980000 742.320000 ;
      RECT 1.100000 727.680000 2029.980000 728.580000 ;
      RECT 0.000000 706.010000 2029.980000 727.680000 ;
      RECT 0.000000 705.110000 2028.880000 706.010000 ;
      RECT 0.000000 691.980000 2029.980000 705.110000 ;
      RECT 1.100000 691.080000 2029.980000 691.980000 ;
      RECT 0.000000 668.800000 2029.980000 691.080000 ;
      RECT 0.000000 667.900000 2028.880000 668.800000 ;
      RECT 0.000000 655.990000 2029.980000 667.900000 ;
      RECT 1.100000 655.090000 2029.980000 655.990000 ;
      RECT 0.000000 632.200000 2029.980000 655.090000 ;
      RECT 0.000000 631.300000 2028.880000 632.200000 ;
      RECT 0.000000 619.390000 2029.980000 631.300000 ;
      RECT 1.100000 618.490000 2029.980000 619.390000 ;
      RECT 0.000000 594.990000 2029.980000 618.490000 ;
      RECT 0.000000 594.090000 2028.880000 594.990000 ;
      RECT 0.000000 582.790000 2029.980000 594.090000 ;
      RECT 1.100000 581.890000 2029.980000 582.790000 ;
      RECT 0.000000 557.780000 2029.980000 581.890000 ;
      RECT 0.000000 556.880000 2028.880000 557.780000 ;
      RECT 0.000000 546.800000 2029.980000 556.880000 ;
      RECT 1.100000 545.900000 2029.980000 546.800000 ;
      RECT 0.000000 520.570000 2029.980000 545.900000 ;
      RECT 0.000000 519.670000 2028.880000 520.570000 ;
      RECT 0.000000 510.200000 2029.980000 519.670000 ;
      RECT 1.100000 509.300000 2029.980000 510.200000 ;
      RECT 0.000000 483.360000 2029.980000 509.300000 ;
      RECT 0.000000 482.460000 2028.880000 483.360000 ;
      RECT 0.000000 473.600000 2029.980000 482.460000 ;
      RECT 1.100000 472.700000 2029.980000 473.600000 ;
      RECT 0.000000 446.150000 2029.980000 472.700000 ;
      RECT 0.000000 445.250000 2028.880000 446.150000 ;
      RECT 0.000000 437.610000 2029.980000 445.250000 ;
      RECT 1.100000 436.710000 2029.980000 437.610000 ;
      RECT 0.000000 409.550000 2029.980000 436.710000 ;
      RECT 0.000000 408.650000 2028.880000 409.550000 ;
      RECT 0.000000 401.010000 2029.980000 408.650000 ;
      RECT 1.100000 400.110000 2029.980000 401.010000 ;
      RECT 0.000000 372.340000 2029.980000 400.110000 ;
      RECT 0.000000 371.440000 2028.880000 372.340000 ;
      RECT 0.000000 364.410000 2029.980000 371.440000 ;
      RECT 1.100000 363.510000 2029.980000 364.410000 ;
      RECT 0.000000 335.130000 2029.980000 363.510000 ;
      RECT 0.000000 334.230000 2028.880000 335.130000 ;
      RECT 0.000000 328.420000 2029.980000 334.230000 ;
      RECT 1.100000 327.520000 2029.980000 328.420000 ;
      RECT 0.000000 297.920000 2029.980000 327.520000 ;
      RECT 0.000000 297.020000 2028.880000 297.920000 ;
      RECT 0.000000 291.820000 2029.980000 297.020000 ;
      RECT 1.100000 290.920000 2029.980000 291.820000 ;
      RECT 0.000000 260.710000 2029.980000 290.920000 ;
      RECT 0.000000 259.810000 2028.880000 260.710000 ;
      RECT 0.000000 255.220000 2029.980000 259.810000 ;
      RECT 1.100000 254.320000 2029.980000 255.220000 ;
      RECT 0.000000 223.500000 2029.980000 254.320000 ;
      RECT 0.000000 222.600000 2028.880000 223.500000 ;
      RECT 0.000000 219.230000 2029.980000 222.600000 ;
      RECT 1.100000 218.330000 2029.980000 219.230000 ;
      RECT 0.000000 186.900000 2029.980000 218.330000 ;
      RECT 0.000000 186.000000 2028.880000 186.900000 ;
      RECT 0.000000 182.630000 2029.980000 186.000000 ;
      RECT 1.100000 181.730000 2029.980000 182.630000 ;
      RECT 0.000000 149.690000 2029.980000 181.730000 ;
      RECT 0.000000 148.790000 2028.880000 149.690000 ;
      RECT 0.000000 146.030000 2029.980000 148.790000 ;
      RECT 1.100000 145.130000 2029.980000 146.030000 ;
      RECT 0.000000 112.480000 2029.980000 145.130000 ;
      RECT 0.000000 111.580000 2028.880000 112.480000 ;
      RECT 0.000000 110.040000 2029.980000 111.580000 ;
      RECT 1.100000 109.140000 2029.980000 110.040000 ;
      RECT 0.000000 75.270000 2029.980000 109.140000 ;
      RECT 0.000000 74.370000 2028.880000 75.270000 ;
      RECT 0.000000 73.440000 2029.980000 74.370000 ;
      RECT 1.100000 72.540000 2029.980000 73.440000 ;
      RECT 0.000000 38.060000 2029.980000 72.540000 ;
      RECT 0.000000 37.160000 2028.880000 38.060000 ;
      RECT 0.000000 36.840000 2029.980000 37.160000 ;
      RECT 1.100000 35.940000 2029.980000 36.840000 ;
      RECT 0.000000 5.120000 2029.980000 35.940000 ;
      RECT 1.100000 4.220000 2028.880000 5.120000 ;
      RECT 0.000000 1.100000 2029.980000 4.220000 ;
      RECT 2028.360000 0.000000 2029.980000 1.100000 ;
      RECT 2026.520000 0.000000 2027.460000 1.100000 ;
      RECT 2022.380000 0.000000 2025.620000 1.100000 ;
      RECT 2018.240000 0.000000 2021.480000 1.100000 ;
      RECT 2014.100000 0.000000 2017.340000 1.100000 ;
      RECT 2009.960000 0.000000 2013.200000 1.100000 ;
      RECT 2005.820000 0.000000 2009.060000 1.100000 ;
      RECT 2001.680000 0.000000 2004.920000 1.100000 ;
      RECT 1997.540000 0.000000 2000.780000 1.100000 ;
      RECT 1993.400000 0.000000 1996.640000 1.100000 ;
      RECT 1989.260000 0.000000 1992.500000 1.100000 ;
      RECT 1985.120000 0.000000 1988.360000 1.100000 ;
      RECT 1980.980000 0.000000 1984.220000 1.100000 ;
      RECT 1976.840000 0.000000 1980.080000 1.100000 ;
      RECT 1972.700000 0.000000 1975.940000 1.100000 ;
      RECT 1968.560000 0.000000 1971.800000 1.100000 ;
      RECT 1964.420000 0.000000 1967.660000 1.100000 ;
      RECT 1960.280000 0.000000 1963.520000 1.100000 ;
      RECT 1956.140000 0.000000 1959.380000 1.100000 ;
      RECT 1952.000000 0.000000 1955.240000 1.100000 ;
      RECT 1948.320000 0.000000 1951.100000 1.100000 ;
      RECT 1944.180000 0.000000 1947.420000 1.100000 ;
      RECT 1940.040000 0.000000 1943.280000 1.100000 ;
      RECT 1935.900000 0.000000 1939.140000 1.100000 ;
      RECT 1931.760000 0.000000 1935.000000 1.100000 ;
      RECT 1927.620000 0.000000 1930.860000 1.100000 ;
      RECT 1923.480000 0.000000 1926.720000 1.100000 ;
      RECT 1919.340000 0.000000 1922.580000 1.100000 ;
      RECT 1915.200000 0.000000 1918.440000 1.100000 ;
      RECT 1911.060000 0.000000 1914.300000 1.100000 ;
      RECT 1906.920000 0.000000 1910.160000 1.100000 ;
      RECT 1902.780000 0.000000 1906.020000 1.100000 ;
      RECT 1898.640000 0.000000 1901.880000 1.100000 ;
      RECT 1894.500000 0.000000 1897.740000 1.100000 ;
      RECT 1890.360000 0.000000 1893.600000 1.100000 ;
      RECT 1886.220000 0.000000 1889.460000 1.100000 ;
      RECT 1882.080000 0.000000 1885.320000 1.100000 ;
      RECT 1877.940000 0.000000 1881.180000 1.100000 ;
      RECT 1873.800000 0.000000 1877.040000 1.100000 ;
      RECT 1869.660000 0.000000 1872.900000 1.100000 ;
      RECT 1865.980000 0.000000 1868.760000 1.100000 ;
      RECT 1861.840000 0.000000 1865.080000 1.100000 ;
      RECT 1857.700000 0.000000 1860.940000 1.100000 ;
      RECT 1853.560000 0.000000 1856.800000 1.100000 ;
      RECT 1849.420000 0.000000 1852.660000 1.100000 ;
      RECT 1845.280000 0.000000 1848.520000 1.100000 ;
      RECT 1841.140000 0.000000 1844.380000 1.100000 ;
      RECT 1837.000000 0.000000 1840.240000 1.100000 ;
      RECT 1832.860000 0.000000 1836.100000 1.100000 ;
      RECT 1828.720000 0.000000 1831.960000 1.100000 ;
      RECT 1824.580000 0.000000 1827.820000 1.100000 ;
      RECT 1820.440000 0.000000 1823.680000 1.100000 ;
      RECT 1816.300000 0.000000 1819.540000 1.100000 ;
      RECT 1812.160000 0.000000 1815.400000 1.100000 ;
      RECT 1808.020000 0.000000 1811.260000 1.100000 ;
      RECT 1803.880000 0.000000 1807.120000 1.100000 ;
      RECT 1799.740000 0.000000 1802.980000 1.100000 ;
      RECT 1795.600000 0.000000 1798.840000 1.100000 ;
      RECT 1791.460000 0.000000 1794.700000 1.100000 ;
      RECT 1787.320000 0.000000 1790.560000 1.100000 ;
      RECT 1783.640000 0.000000 1786.420000 1.100000 ;
      RECT 1779.500000 0.000000 1782.740000 1.100000 ;
      RECT 1775.360000 0.000000 1778.600000 1.100000 ;
      RECT 1771.220000 0.000000 1774.460000 1.100000 ;
      RECT 1767.080000 0.000000 1770.320000 1.100000 ;
      RECT 1762.940000 0.000000 1766.180000 1.100000 ;
      RECT 1758.800000 0.000000 1762.040000 1.100000 ;
      RECT 1754.660000 0.000000 1757.900000 1.100000 ;
      RECT 1750.520000 0.000000 1753.760000 1.100000 ;
      RECT 1746.380000 0.000000 1749.620000 1.100000 ;
      RECT 1742.240000 0.000000 1745.480000 1.100000 ;
      RECT 1738.100000 0.000000 1741.340000 1.100000 ;
      RECT 1733.960000 0.000000 1737.200000 1.100000 ;
      RECT 1729.820000 0.000000 1733.060000 1.100000 ;
      RECT 1725.680000 0.000000 1728.920000 1.100000 ;
      RECT 1721.540000 0.000000 1724.780000 1.100000 ;
      RECT 1717.400000 0.000000 1720.640000 1.100000 ;
      RECT 1713.260000 0.000000 1716.500000 1.100000 ;
      RECT 1709.120000 0.000000 1712.360000 1.100000 ;
      RECT 1705.440000 0.000000 1708.220000 1.100000 ;
      RECT 1701.300000 0.000000 1704.540000 1.100000 ;
      RECT 1697.160000 0.000000 1700.400000 1.100000 ;
      RECT 1693.020000 0.000000 1696.260000 1.100000 ;
      RECT 1688.880000 0.000000 1692.120000 1.100000 ;
      RECT 1684.740000 0.000000 1687.980000 1.100000 ;
      RECT 1680.600000 0.000000 1683.840000 1.100000 ;
      RECT 1676.460000 0.000000 1679.700000 1.100000 ;
      RECT 1672.320000 0.000000 1675.560000 1.100000 ;
      RECT 1668.180000 0.000000 1671.420000 1.100000 ;
      RECT 1664.040000 0.000000 1667.280000 1.100000 ;
      RECT 1659.900000 0.000000 1663.140000 1.100000 ;
      RECT 1655.760000 0.000000 1659.000000 1.100000 ;
      RECT 1651.620000 0.000000 1654.860000 1.100000 ;
      RECT 1647.480000 0.000000 1650.720000 1.100000 ;
      RECT 1643.340000 0.000000 1646.580000 1.100000 ;
      RECT 1639.200000 0.000000 1642.440000 1.100000 ;
      RECT 1635.060000 0.000000 1638.300000 1.100000 ;
      RECT 1630.920000 0.000000 1634.160000 1.100000 ;
      RECT 1626.780000 0.000000 1630.020000 1.100000 ;
      RECT 1623.100000 0.000000 1625.880000 1.100000 ;
      RECT 1618.960000 0.000000 1622.200000 1.100000 ;
      RECT 1614.820000 0.000000 1618.060000 1.100000 ;
      RECT 1610.680000 0.000000 1613.920000 1.100000 ;
      RECT 1606.540000 0.000000 1609.780000 1.100000 ;
      RECT 1602.400000 0.000000 1605.640000 1.100000 ;
      RECT 1598.260000 0.000000 1601.500000 1.100000 ;
      RECT 1594.120000 0.000000 1597.360000 1.100000 ;
      RECT 1589.980000 0.000000 1593.220000 1.100000 ;
      RECT 1585.840000 0.000000 1589.080000 1.100000 ;
      RECT 1581.700000 0.000000 1584.940000 1.100000 ;
      RECT 1577.560000 0.000000 1580.800000 1.100000 ;
      RECT 1573.420000 0.000000 1576.660000 1.100000 ;
      RECT 1569.280000 0.000000 1572.520000 1.100000 ;
      RECT 1565.140000 0.000000 1568.380000 1.100000 ;
      RECT 1561.000000 0.000000 1564.240000 1.100000 ;
      RECT 1556.860000 0.000000 1560.100000 1.100000 ;
      RECT 1552.720000 0.000000 1555.960000 1.100000 ;
      RECT 1548.580000 0.000000 1551.820000 1.100000 ;
      RECT 1544.440000 0.000000 1547.680000 1.100000 ;
      RECT 1540.760000 0.000000 1543.540000 1.100000 ;
      RECT 1536.620000 0.000000 1539.860000 1.100000 ;
      RECT 1532.480000 0.000000 1535.720000 1.100000 ;
      RECT 1528.340000 0.000000 1531.580000 1.100000 ;
      RECT 1524.200000 0.000000 1527.440000 1.100000 ;
      RECT 1520.060000 0.000000 1523.300000 1.100000 ;
      RECT 1515.920000 0.000000 1519.160000 1.100000 ;
      RECT 1511.780000 0.000000 1515.020000 1.100000 ;
      RECT 1507.640000 0.000000 1510.880000 1.100000 ;
      RECT 1503.500000 0.000000 1506.740000 1.100000 ;
      RECT 1499.360000 0.000000 1502.600000 1.100000 ;
      RECT 1495.220000 0.000000 1498.460000 1.100000 ;
      RECT 1491.080000 0.000000 1494.320000 1.100000 ;
      RECT 1486.940000 0.000000 1490.180000 1.100000 ;
      RECT 1482.800000 0.000000 1486.040000 1.100000 ;
      RECT 1478.660000 0.000000 1481.900000 1.100000 ;
      RECT 1474.520000 0.000000 1477.760000 1.100000 ;
      RECT 1470.380000 0.000000 1473.620000 1.100000 ;
      RECT 1466.240000 0.000000 1469.480000 1.100000 ;
      RECT 1462.100000 0.000000 1465.340000 1.100000 ;
      RECT 1458.420000 0.000000 1461.200000 1.100000 ;
      RECT 1454.280000 0.000000 1457.520000 1.100000 ;
      RECT 1450.140000 0.000000 1453.380000 1.100000 ;
      RECT 1446.000000 0.000000 1449.240000 1.100000 ;
      RECT 1441.860000 0.000000 1445.100000 1.100000 ;
      RECT 1437.720000 0.000000 1440.960000 1.100000 ;
      RECT 1433.580000 0.000000 1436.820000 1.100000 ;
      RECT 1429.440000 0.000000 1432.680000 1.100000 ;
      RECT 1425.300000 0.000000 1428.540000 1.100000 ;
      RECT 1421.160000 0.000000 1424.400000 1.100000 ;
      RECT 1417.020000 0.000000 1420.260000 1.100000 ;
      RECT 1412.880000 0.000000 1416.120000 1.100000 ;
      RECT 1408.740000 0.000000 1411.980000 1.100000 ;
      RECT 1404.600000 0.000000 1407.840000 1.100000 ;
      RECT 1400.460000 0.000000 1403.700000 1.100000 ;
      RECT 1396.320000 0.000000 1399.560000 1.100000 ;
      RECT 1392.180000 0.000000 1395.420000 1.100000 ;
      RECT 1388.040000 0.000000 1391.280000 1.100000 ;
      RECT 1383.900000 0.000000 1387.140000 1.100000 ;
      RECT 1380.220000 0.000000 1383.000000 1.100000 ;
      RECT 1376.080000 0.000000 1379.320000 1.100000 ;
      RECT 1371.940000 0.000000 1375.180000 1.100000 ;
      RECT 1367.800000 0.000000 1371.040000 1.100000 ;
      RECT 1363.660000 0.000000 1366.900000 1.100000 ;
      RECT 1359.520000 0.000000 1362.760000 1.100000 ;
      RECT 1355.380000 0.000000 1358.620000 1.100000 ;
      RECT 1351.240000 0.000000 1354.480000 1.100000 ;
      RECT 1347.100000 0.000000 1350.340000 1.100000 ;
      RECT 1342.960000 0.000000 1346.200000 1.100000 ;
      RECT 1338.820000 0.000000 1342.060000 1.100000 ;
      RECT 1334.680000 0.000000 1337.920000 1.100000 ;
      RECT 1330.540000 0.000000 1333.780000 1.100000 ;
      RECT 1326.400000 0.000000 1329.640000 1.100000 ;
      RECT 1322.260000 0.000000 1325.500000 1.100000 ;
      RECT 1318.120000 0.000000 1321.360000 1.100000 ;
      RECT 1313.980000 0.000000 1317.220000 1.100000 ;
      RECT 1309.840000 0.000000 1313.080000 1.100000 ;
      RECT 1305.700000 0.000000 1308.940000 1.100000 ;
      RECT 1301.560000 0.000000 1304.800000 1.100000 ;
      RECT 1297.880000 0.000000 1300.660000 1.100000 ;
      RECT 1293.740000 0.000000 1296.980000 1.100000 ;
      RECT 1289.600000 0.000000 1292.840000 1.100000 ;
      RECT 1285.460000 0.000000 1288.700000 1.100000 ;
      RECT 1281.320000 0.000000 1284.560000 1.100000 ;
      RECT 1277.180000 0.000000 1280.420000 1.100000 ;
      RECT 1273.040000 0.000000 1276.280000 1.100000 ;
      RECT 1268.900000 0.000000 1272.140000 1.100000 ;
      RECT 1264.760000 0.000000 1268.000000 1.100000 ;
      RECT 1260.620000 0.000000 1263.860000 1.100000 ;
      RECT 1256.480000 0.000000 1259.720000 1.100000 ;
      RECT 1252.340000 0.000000 1255.580000 1.100000 ;
      RECT 1248.200000 0.000000 1251.440000 1.100000 ;
      RECT 1244.060000 0.000000 1247.300000 1.100000 ;
      RECT 1239.920000 0.000000 1243.160000 1.100000 ;
      RECT 1235.780000 0.000000 1239.020000 1.100000 ;
      RECT 1231.640000 0.000000 1234.880000 1.100000 ;
      RECT 1227.500000 0.000000 1230.740000 1.100000 ;
      RECT 1223.360000 0.000000 1226.600000 1.100000 ;
      RECT 1219.220000 0.000000 1222.460000 1.100000 ;
      RECT 1215.540000 0.000000 1218.320000 1.100000 ;
      RECT 1211.400000 0.000000 1214.640000 1.100000 ;
      RECT 1207.260000 0.000000 1210.500000 1.100000 ;
      RECT 1203.120000 0.000000 1206.360000 1.100000 ;
      RECT 1198.980000 0.000000 1202.220000 1.100000 ;
      RECT 1194.840000 0.000000 1198.080000 1.100000 ;
      RECT 1190.700000 0.000000 1193.940000 1.100000 ;
      RECT 1186.560000 0.000000 1189.800000 1.100000 ;
      RECT 1182.420000 0.000000 1185.660000 1.100000 ;
      RECT 1178.280000 0.000000 1181.520000 1.100000 ;
      RECT 1174.140000 0.000000 1177.380000 1.100000 ;
      RECT 1170.000000 0.000000 1173.240000 1.100000 ;
      RECT 1165.860000 0.000000 1169.100000 1.100000 ;
      RECT 1161.720000 0.000000 1164.960000 1.100000 ;
      RECT 1157.580000 0.000000 1160.820000 1.100000 ;
      RECT 1153.440000 0.000000 1156.680000 1.100000 ;
      RECT 1149.300000 0.000000 1152.540000 1.100000 ;
      RECT 1145.160000 0.000000 1148.400000 1.100000 ;
      RECT 1141.020000 0.000000 1144.260000 1.100000 ;
      RECT 1137.340000 0.000000 1140.120000 1.100000 ;
      RECT 1133.200000 0.000000 1136.440000 1.100000 ;
      RECT 1129.060000 0.000000 1132.300000 1.100000 ;
      RECT 1124.920000 0.000000 1128.160000 1.100000 ;
      RECT 1120.780000 0.000000 1124.020000 1.100000 ;
      RECT 1116.640000 0.000000 1119.880000 1.100000 ;
      RECT 1112.500000 0.000000 1115.740000 1.100000 ;
      RECT 1108.360000 0.000000 1111.600000 1.100000 ;
      RECT 1104.220000 0.000000 1107.460000 1.100000 ;
      RECT 1100.080000 0.000000 1103.320000 1.100000 ;
      RECT 1095.940000 0.000000 1099.180000 1.100000 ;
      RECT 1091.800000 0.000000 1095.040000 1.100000 ;
      RECT 1087.660000 0.000000 1090.900000 1.100000 ;
      RECT 1083.520000 0.000000 1086.760000 1.100000 ;
      RECT 1079.380000 0.000000 1082.620000 1.100000 ;
      RECT 1075.240000 0.000000 1078.480000 1.100000 ;
      RECT 1071.100000 0.000000 1074.340000 1.100000 ;
      RECT 1066.960000 0.000000 1070.200000 1.100000 ;
      RECT 1062.820000 0.000000 1066.060000 1.100000 ;
      RECT 1058.680000 0.000000 1061.920000 1.100000 ;
      RECT 1055.000000 0.000000 1057.780000 1.100000 ;
      RECT 1050.860000 0.000000 1054.100000 1.100000 ;
      RECT 1046.720000 0.000000 1049.960000 1.100000 ;
      RECT 1042.580000 0.000000 1045.820000 1.100000 ;
      RECT 1038.440000 0.000000 1041.680000 1.100000 ;
      RECT 1034.300000 0.000000 1037.540000 1.100000 ;
      RECT 1030.160000 0.000000 1033.400000 1.100000 ;
      RECT 1026.020000 0.000000 1029.260000 1.100000 ;
      RECT 1021.880000 0.000000 1025.120000 1.100000 ;
      RECT 1017.740000 0.000000 1020.980000 1.100000 ;
      RECT 1013.600000 0.000000 1016.840000 1.100000 ;
      RECT 1009.460000 0.000000 1012.700000 1.100000 ;
      RECT 1005.320000 0.000000 1008.560000 1.100000 ;
      RECT 1001.180000 0.000000 1004.420000 1.100000 ;
      RECT 997.040000 0.000000 1000.280000 1.100000 ;
      RECT 992.900000 0.000000 996.140000 1.100000 ;
      RECT 988.760000 0.000000 992.000000 1.100000 ;
      RECT 984.620000 0.000000 987.860000 1.100000 ;
      RECT 980.480000 0.000000 983.720000 1.100000 ;
      RECT 976.340000 0.000000 979.580000 1.100000 ;
      RECT 972.660000 0.000000 975.440000 1.100000 ;
      RECT 968.520000 0.000000 971.760000 1.100000 ;
      RECT 964.380000 0.000000 967.620000 1.100000 ;
      RECT 960.240000 0.000000 963.480000 1.100000 ;
      RECT 956.100000 0.000000 959.340000 1.100000 ;
      RECT 951.960000 0.000000 955.200000 1.100000 ;
      RECT 947.820000 0.000000 951.060000 1.100000 ;
      RECT 943.680000 0.000000 946.920000 1.100000 ;
      RECT 939.540000 0.000000 942.780000 1.100000 ;
      RECT 935.400000 0.000000 938.640000 1.100000 ;
      RECT 931.260000 0.000000 934.500000 1.100000 ;
      RECT 927.120000 0.000000 930.360000 1.100000 ;
      RECT 922.980000 0.000000 926.220000 1.100000 ;
      RECT 918.840000 0.000000 922.080000 1.100000 ;
      RECT 914.700000 0.000000 917.940000 1.100000 ;
      RECT 910.560000 0.000000 913.800000 1.100000 ;
      RECT 906.420000 0.000000 909.660000 1.100000 ;
      RECT 902.280000 0.000000 905.520000 1.100000 ;
      RECT 898.140000 0.000000 901.380000 1.100000 ;
      RECT 894.000000 0.000000 897.240000 1.100000 ;
      RECT 890.320000 0.000000 893.100000 1.100000 ;
      RECT 886.180000 0.000000 889.420000 1.100000 ;
      RECT 882.040000 0.000000 885.280000 1.100000 ;
      RECT 877.900000 0.000000 881.140000 1.100000 ;
      RECT 873.760000 0.000000 877.000000 1.100000 ;
      RECT 869.620000 0.000000 872.860000 1.100000 ;
      RECT 865.480000 0.000000 868.720000 1.100000 ;
      RECT 861.340000 0.000000 864.580000 1.100000 ;
      RECT 857.200000 0.000000 860.440000 1.100000 ;
      RECT 853.060000 0.000000 856.300000 1.100000 ;
      RECT 848.920000 0.000000 852.160000 1.100000 ;
      RECT 844.780000 0.000000 848.020000 1.100000 ;
      RECT 840.640000 0.000000 843.880000 1.100000 ;
      RECT 836.500000 0.000000 839.740000 1.100000 ;
      RECT 832.360000 0.000000 835.600000 1.100000 ;
      RECT 828.220000 0.000000 831.460000 1.100000 ;
      RECT 824.080000 0.000000 827.320000 1.100000 ;
      RECT 819.940000 0.000000 823.180000 1.100000 ;
      RECT 815.800000 0.000000 819.040000 1.100000 ;
      RECT 812.120000 0.000000 814.900000 1.100000 ;
      RECT 807.980000 0.000000 811.220000 1.100000 ;
      RECT 803.840000 0.000000 807.080000 1.100000 ;
      RECT 799.700000 0.000000 802.940000 1.100000 ;
      RECT 795.560000 0.000000 798.800000 1.100000 ;
      RECT 791.420000 0.000000 794.660000 1.100000 ;
      RECT 787.280000 0.000000 790.520000 1.100000 ;
      RECT 783.140000 0.000000 786.380000 1.100000 ;
      RECT 779.000000 0.000000 782.240000 1.100000 ;
      RECT 774.860000 0.000000 778.100000 1.100000 ;
      RECT 770.720000 0.000000 773.960000 1.100000 ;
      RECT 766.580000 0.000000 769.820000 1.100000 ;
      RECT 762.440000 0.000000 765.680000 1.100000 ;
      RECT 758.300000 0.000000 761.540000 1.100000 ;
      RECT 754.160000 0.000000 757.400000 1.100000 ;
      RECT 750.020000 0.000000 753.260000 1.100000 ;
      RECT 745.880000 0.000000 749.120000 1.100000 ;
      RECT 741.740000 0.000000 744.980000 1.100000 ;
      RECT 737.600000 0.000000 740.840000 1.100000 ;
      RECT 733.460000 0.000000 736.700000 1.100000 ;
      RECT 729.780000 0.000000 732.560000 1.100000 ;
      RECT 725.640000 0.000000 728.880000 1.100000 ;
      RECT 721.500000 0.000000 724.740000 1.100000 ;
      RECT 717.360000 0.000000 720.600000 1.100000 ;
      RECT 713.220000 0.000000 716.460000 1.100000 ;
      RECT 709.080000 0.000000 712.320000 1.100000 ;
      RECT 704.940000 0.000000 708.180000 1.100000 ;
      RECT 700.800000 0.000000 704.040000 1.100000 ;
      RECT 696.660000 0.000000 699.900000 1.100000 ;
      RECT 692.520000 0.000000 695.760000 1.100000 ;
      RECT 688.380000 0.000000 691.620000 1.100000 ;
      RECT 684.240000 0.000000 687.480000 1.100000 ;
      RECT 680.100000 0.000000 683.340000 1.100000 ;
      RECT 675.960000 0.000000 679.200000 1.100000 ;
      RECT 671.820000 0.000000 675.060000 1.100000 ;
      RECT 667.680000 0.000000 670.920000 1.100000 ;
      RECT 663.540000 0.000000 666.780000 1.100000 ;
      RECT 659.400000 0.000000 662.640000 1.100000 ;
      RECT 655.260000 0.000000 658.500000 1.100000 ;
      RECT 651.120000 0.000000 654.360000 1.100000 ;
      RECT 647.440000 0.000000 650.220000 1.100000 ;
      RECT 643.300000 0.000000 646.540000 1.100000 ;
      RECT 639.160000 0.000000 642.400000 1.100000 ;
      RECT 635.020000 0.000000 638.260000 1.100000 ;
      RECT 630.880000 0.000000 634.120000 1.100000 ;
      RECT 626.740000 0.000000 629.980000 1.100000 ;
      RECT 622.600000 0.000000 625.840000 1.100000 ;
      RECT 618.460000 0.000000 621.700000 1.100000 ;
      RECT 614.320000 0.000000 617.560000 1.100000 ;
      RECT 610.180000 0.000000 613.420000 1.100000 ;
      RECT 606.040000 0.000000 609.280000 1.100000 ;
      RECT 601.900000 0.000000 605.140000 1.100000 ;
      RECT 597.760000 0.000000 601.000000 1.100000 ;
      RECT 593.620000 0.000000 596.860000 1.100000 ;
      RECT 589.480000 0.000000 592.720000 1.100000 ;
      RECT 585.340000 0.000000 588.580000 1.100000 ;
      RECT 581.200000 0.000000 584.440000 1.100000 ;
      RECT 577.060000 0.000000 580.300000 1.100000 ;
      RECT 572.920000 0.000000 576.160000 1.100000 ;
      RECT 569.240000 0.000000 572.020000 1.100000 ;
      RECT 565.100000 0.000000 568.340000 1.100000 ;
      RECT 560.960000 0.000000 564.200000 1.100000 ;
      RECT 556.820000 0.000000 560.060000 1.100000 ;
      RECT 552.680000 0.000000 555.920000 1.100000 ;
      RECT 548.540000 0.000000 551.780000 1.100000 ;
      RECT 544.400000 0.000000 547.640000 1.100000 ;
      RECT 540.260000 0.000000 543.500000 1.100000 ;
      RECT 536.120000 0.000000 539.360000 1.100000 ;
      RECT 531.980000 0.000000 535.220000 1.100000 ;
      RECT 527.840000 0.000000 531.080000 1.100000 ;
      RECT 523.700000 0.000000 526.940000 1.100000 ;
      RECT 519.560000 0.000000 522.800000 1.100000 ;
      RECT 515.420000 0.000000 518.660000 1.100000 ;
      RECT 511.280000 0.000000 514.520000 1.100000 ;
      RECT 507.140000 0.000000 510.380000 1.100000 ;
      RECT 503.000000 0.000000 506.240000 1.100000 ;
      RECT 498.860000 0.000000 502.100000 1.100000 ;
      RECT 494.720000 0.000000 497.960000 1.100000 ;
      RECT 490.580000 0.000000 493.820000 1.100000 ;
      RECT 486.900000 0.000000 489.680000 1.100000 ;
      RECT 482.760000 0.000000 486.000000 1.100000 ;
      RECT 478.620000 0.000000 481.860000 1.100000 ;
      RECT 474.480000 0.000000 477.720000 1.100000 ;
      RECT 470.340000 0.000000 473.580000 1.100000 ;
      RECT 466.200000 0.000000 469.440000 1.100000 ;
      RECT 462.060000 0.000000 465.300000 1.100000 ;
      RECT 457.920000 0.000000 461.160000 1.100000 ;
      RECT 453.780000 0.000000 457.020000 1.100000 ;
      RECT 449.640000 0.000000 452.880000 1.100000 ;
      RECT 445.500000 0.000000 448.740000 1.100000 ;
      RECT 441.360000 0.000000 444.600000 1.100000 ;
      RECT 437.220000 0.000000 440.460000 1.100000 ;
      RECT 433.080000 0.000000 436.320000 1.100000 ;
      RECT 428.940000 0.000000 432.180000 1.100000 ;
      RECT 424.800000 0.000000 428.040000 1.100000 ;
      RECT 420.660000 0.000000 423.900000 1.100000 ;
      RECT 416.520000 0.000000 419.760000 1.100000 ;
      RECT 412.380000 0.000000 415.620000 1.100000 ;
      RECT 408.240000 0.000000 411.480000 1.100000 ;
      RECT 404.560000 0.000000 407.340000 1.100000 ;
      RECT 400.420000 0.000000 403.660000 1.100000 ;
      RECT 396.280000 0.000000 399.520000 1.100000 ;
      RECT 392.140000 0.000000 395.380000 1.100000 ;
      RECT 388.000000 0.000000 391.240000 1.100000 ;
      RECT 383.860000 0.000000 387.100000 1.100000 ;
      RECT 379.720000 0.000000 382.960000 1.100000 ;
      RECT 375.580000 0.000000 378.820000 1.100000 ;
      RECT 371.440000 0.000000 374.680000 1.100000 ;
      RECT 367.300000 0.000000 370.540000 1.100000 ;
      RECT 363.160000 0.000000 366.400000 1.100000 ;
      RECT 359.020000 0.000000 362.260000 1.100000 ;
      RECT 354.880000 0.000000 358.120000 1.100000 ;
      RECT 350.740000 0.000000 353.980000 1.100000 ;
      RECT 346.600000 0.000000 349.840000 1.100000 ;
      RECT 342.460000 0.000000 345.700000 1.100000 ;
      RECT 338.320000 0.000000 341.560000 1.100000 ;
      RECT 334.180000 0.000000 337.420000 1.100000 ;
      RECT 330.040000 0.000000 333.280000 1.100000 ;
      RECT 325.900000 0.000000 329.140000 1.100000 ;
      RECT 322.220000 0.000000 325.000000 1.100000 ;
      RECT 318.080000 0.000000 321.320000 1.100000 ;
      RECT 313.940000 0.000000 317.180000 1.100000 ;
      RECT 309.800000 0.000000 313.040000 1.100000 ;
      RECT 305.660000 0.000000 308.900000 1.100000 ;
      RECT 301.520000 0.000000 304.760000 1.100000 ;
      RECT 297.380000 0.000000 300.620000 1.100000 ;
      RECT 293.240000 0.000000 296.480000 1.100000 ;
      RECT 289.100000 0.000000 292.340000 1.100000 ;
      RECT 284.960000 0.000000 288.200000 1.100000 ;
      RECT 280.820000 0.000000 284.060000 1.100000 ;
      RECT 276.680000 0.000000 279.920000 1.100000 ;
      RECT 272.540000 0.000000 275.780000 1.100000 ;
      RECT 268.400000 0.000000 271.640000 1.100000 ;
      RECT 264.260000 0.000000 267.500000 1.100000 ;
      RECT 260.120000 0.000000 263.360000 1.100000 ;
      RECT 255.980000 0.000000 259.220000 1.100000 ;
      RECT 251.840000 0.000000 255.080000 1.100000 ;
      RECT 247.700000 0.000000 250.940000 1.100000 ;
      RECT 244.020000 0.000000 246.800000 1.100000 ;
      RECT 239.880000 0.000000 243.120000 1.100000 ;
      RECT 235.740000 0.000000 238.980000 1.100000 ;
      RECT 231.600000 0.000000 234.840000 1.100000 ;
      RECT 227.460000 0.000000 230.700000 1.100000 ;
      RECT 223.320000 0.000000 226.560000 1.100000 ;
      RECT 219.180000 0.000000 222.420000 1.100000 ;
      RECT 215.040000 0.000000 218.280000 1.100000 ;
      RECT 210.900000 0.000000 214.140000 1.100000 ;
      RECT 206.760000 0.000000 210.000000 1.100000 ;
      RECT 202.620000 0.000000 205.860000 1.100000 ;
      RECT 198.480000 0.000000 201.720000 1.100000 ;
      RECT 194.340000 0.000000 197.580000 1.100000 ;
      RECT 190.200000 0.000000 193.440000 1.100000 ;
      RECT 186.060000 0.000000 189.300000 1.100000 ;
      RECT 181.920000 0.000000 185.160000 1.100000 ;
      RECT 177.780000 0.000000 181.020000 1.100000 ;
      RECT 173.640000 0.000000 176.880000 1.100000 ;
      RECT 169.500000 0.000000 172.740000 1.100000 ;
      RECT 165.360000 0.000000 168.600000 1.100000 ;
      RECT 161.680000 0.000000 164.460000 1.100000 ;
      RECT 157.540000 0.000000 160.780000 1.100000 ;
      RECT 153.400000 0.000000 156.640000 1.100000 ;
      RECT 149.260000 0.000000 152.500000 1.100000 ;
      RECT 145.120000 0.000000 148.360000 1.100000 ;
      RECT 140.980000 0.000000 144.220000 1.100000 ;
      RECT 136.840000 0.000000 140.080000 1.100000 ;
      RECT 132.700000 0.000000 135.940000 1.100000 ;
      RECT 128.560000 0.000000 131.800000 1.100000 ;
      RECT 124.420000 0.000000 127.660000 1.100000 ;
      RECT 120.280000 0.000000 123.520000 1.100000 ;
      RECT 116.140000 0.000000 119.380000 1.100000 ;
      RECT 112.000000 0.000000 115.240000 1.100000 ;
      RECT 107.860000 0.000000 111.100000 1.100000 ;
      RECT 103.720000 0.000000 106.960000 1.100000 ;
      RECT 99.580000 0.000000 102.820000 1.100000 ;
      RECT 95.440000 0.000000 98.680000 1.100000 ;
      RECT 91.300000 0.000000 94.540000 1.100000 ;
      RECT 87.160000 0.000000 90.400000 1.100000 ;
      RECT 83.020000 0.000000 86.260000 1.100000 ;
      RECT 79.340000 0.000000 82.120000 1.100000 ;
      RECT 75.200000 0.000000 78.440000 1.100000 ;
      RECT 71.060000 0.000000 74.300000 1.100000 ;
      RECT 66.920000 0.000000 70.160000 1.100000 ;
      RECT 62.780000 0.000000 66.020000 1.100000 ;
      RECT 58.640000 0.000000 61.880000 1.100000 ;
      RECT 54.500000 0.000000 57.740000 1.100000 ;
      RECT 50.360000 0.000000 53.600000 1.100000 ;
      RECT 46.220000 0.000000 49.460000 1.100000 ;
      RECT 42.080000 0.000000 45.320000 1.100000 ;
      RECT 37.940000 0.000000 41.180000 1.100000 ;
      RECT 33.800000 0.000000 37.040000 1.100000 ;
      RECT 29.660000 0.000000 32.900000 1.100000 ;
      RECT 25.520000 0.000000 28.760000 1.100000 ;
      RECT 21.380000 0.000000 24.620000 1.100000 ;
      RECT 17.240000 0.000000 20.480000 1.100000 ;
      RECT 13.100000 0.000000 16.340000 1.100000 ;
      RECT 8.960000 0.000000 12.200000 1.100000 ;
      RECT 4.820000 0.000000 8.060000 1.100000 ;
      RECT 2.060000 0.000000 3.920000 1.100000 ;
      RECT 0.000000 0.000000 1.160000 1.100000 ;
    LAYER met4 ;
      RECT 0.000000 1927.020000 2029.980000 1929.840000 ;
      RECT 0.000000 1923.820000 2026.660000 1927.020000 ;
      RECT 2025.660000 4.660000 2026.660000 1923.820000 ;
      RECT 6.520000 4.660000 2023.460000 1923.820000 ;
      RECT 0.000000 4.660000 4.320000 1923.820000 ;
      RECT 2028.860000 1.460000 2029.980000 1927.020000 ;
      RECT 0.000000 1.460000 2026.660000 4.660000 ;
      RECT 0.000000 0.000000 2029.980000 1.460000 ;
    LAYER met5 ;
      RECT 0.000000 0.000000 2029.980000 1929.840000 ;
  END
END azadi_soc_top_caravel

END LIBRARY
