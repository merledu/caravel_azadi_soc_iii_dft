magic
tech sky130A
magscale 1 2
timestamp 1654179656
<< metal1 >>
rect 1394 448536 1400 448588
rect 1452 448576 1458 448588
rect 57606 448576 57612 448588
rect 1452 448548 57612 448576
rect 1452 448536 1458 448548
rect 57606 448536 57612 448548
rect 57664 448536 57670 448588
rect 314286 59780 314292 59832
rect 314344 59820 314350 59832
rect 315390 59820 315396 59832
rect 314344 59792 315396 59820
rect 314344 59780 314350 59792
rect 315390 59780 315396 59792
rect 315448 59780 315454 59832
rect 357526 59780 357532 59832
rect 357584 59820 357590 59832
rect 359458 59820 359464 59832
rect 357584 59792 359464 59820
rect 357584 59780 357590 59792
rect 359458 59780 359464 59792
rect 359516 59780 359522 59832
rect 422386 59780 422392 59832
rect 422444 59820 422450 59832
rect 424134 59820 424140 59832
rect 422444 59792 424140 59820
rect 422444 59780 422450 59792
rect 424134 59780 424140 59792
rect 424192 59780 424198 59832
rect 63402 59712 63408 59764
rect 63460 59752 63466 59764
rect 64230 59752 64236 59764
rect 63460 59724 64236 59752
rect 63460 59712 63466 59724
rect 64230 59712 64236 59724
rect 64288 59712 64294 59764
rect 67542 59712 67548 59764
rect 67600 59752 67606 59764
rect 68462 59752 68468 59764
rect 67600 59724 68468 59752
rect 67600 59712 67606 59724
rect 68462 59712 68468 59724
rect 68520 59712 68526 59764
rect 68922 59712 68928 59764
rect 68980 59752 68986 59764
rect 70118 59752 70124 59764
rect 68980 59724 70124 59752
rect 68980 59712 68986 59724
rect 70118 59712 70124 59724
rect 70176 59712 70182 59764
rect 72694 59712 72700 59764
rect 72752 59752 72758 59764
rect 74626 59752 74632 59764
rect 72752 59724 74632 59752
rect 72752 59712 72758 59724
rect 74626 59712 74632 59724
rect 74684 59712 74690 59764
rect 81066 59712 81072 59764
rect 81124 59752 81130 59764
rect 83458 59752 83464 59764
rect 81124 59724 83464 59752
rect 81124 59712 81130 59724
rect 83458 59712 83464 59724
rect 83516 59712 83522 59764
rect 86218 59712 86224 59764
rect 86276 59752 86282 59764
rect 88426 59752 88432 59764
rect 86276 59724 88432 59752
rect 86276 59712 86282 59724
rect 88426 59712 88432 59724
rect 88484 59712 88490 59764
rect 88978 59712 88984 59764
rect 89036 59752 89042 59764
rect 91738 59752 91744 59764
rect 89036 59724 91744 59752
rect 89036 59712 89042 59724
rect 91738 59712 91744 59724
rect 91796 59712 91802 59764
rect 96062 59712 96068 59764
rect 96120 59752 96126 59764
rect 98362 59752 98368 59764
rect 96120 59724 98368 59752
rect 96120 59712 96126 59724
rect 98362 59712 98368 59724
rect 98420 59712 98426 59764
rect 98638 59712 98644 59764
rect 98696 59752 98702 59764
rect 100846 59752 100852 59764
rect 98696 59724 100852 59752
rect 98696 59712 98702 59724
rect 100846 59712 100852 59724
rect 100904 59712 100910 59764
rect 113082 59712 113088 59764
rect 113140 59752 113146 59764
rect 115014 59752 115020 59764
rect 113140 59724 115020 59752
rect 113140 59712 113146 59724
rect 115014 59712 115020 59724
rect 115072 59712 115078 59764
rect 122742 59712 122748 59764
rect 122800 59752 122806 59764
rect 123294 59752 123300 59764
rect 122800 59724 123300 59752
rect 122800 59712 122806 59724
rect 123294 59712 123300 59724
rect 123352 59712 123358 59764
rect 125134 59712 125140 59764
rect 125192 59752 125198 59764
rect 127526 59752 127532 59764
rect 125192 59724 127532 59752
rect 125192 59712 125198 59724
rect 127526 59712 127532 59724
rect 127584 59712 127590 59764
rect 134518 59712 134524 59764
rect 134576 59752 134582 59764
rect 136634 59752 136640 59764
rect 134576 59724 136640 59752
rect 134576 59712 134582 59724
rect 136634 59712 136640 59724
rect 136692 59712 136698 59764
rect 140222 59712 140228 59764
rect 140280 59752 140286 59764
rect 142430 59752 142436 59764
rect 140280 59724 142436 59752
rect 140280 59712 140286 59724
rect 142430 59712 142436 59724
rect 142488 59712 142494 59764
rect 148502 59712 148508 59764
rect 148560 59752 148566 59764
rect 149422 59752 149428 59764
rect 148560 59724 149428 59752
rect 148560 59712 148566 59724
rect 149422 59712 149428 59724
rect 149480 59712 149486 59764
rect 151722 59712 151728 59764
rect 151780 59752 151786 59764
rect 152458 59752 152464 59764
rect 151780 59724 152464 59752
rect 151780 59712 151786 59724
rect 152458 59712 152464 59724
rect 152516 59712 152522 59764
rect 154298 59712 154304 59764
rect 154356 59752 154362 59764
rect 156598 59752 156604 59764
rect 154356 59724 156604 59752
rect 154356 59712 154362 59724
rect 156598 59712 156604 59724
rect 156656 59712 156662 59764
rect 158530 59712 158536 59764
rect 158588 59752 158594 59764
rect 160738 59752 160744 59764
rect 158588 59724 160744 59752
rect 158588 59712 158594 59724
rect 160738 59712 160744 59724
rect 160796 59712 160802 59764
rect 165246 59712 165252 59764
rect 165304 59752 165310 59764
rect 167454 59752 167460 59764
rect 165304 59724 167460 59752
rect 165304 59712 165310 59724
rect 167454 59712 167460 59724
rect 167512 59712 167518 59764
rect 173618 59712 173624 59764
rect 173676 59752 173682 59764
rect 175734 59752 175740 59764
rect 173676 59724 175740 59752
rect 173676 59712 173682 59724
rect 175734 59712 175740 59724
rect 175792 59712 175798 59764
rect 180610 59712 180616 59764
rect 180668 59752 180674 59764
rect 182358 59752 182364 59764
rect 180668 59724 182364 59752
rect 180668 59712 180674 59724
rect 182358 59712 182364 59724
rect 182416 59712 182422 59764
rect 184566 59712 184572 59764
rect 184624 59752 184630 59764
rect 185670 59752 185676 59764
rect 184624 59724 185676 59752
rect 184624 59712 184630 59724
rect 185670 59712 185676 59724
rect 185728 59712 185734 59764
rect 188706 59712 188712 59764
rect 188764 59752 188770 59764
rect 189902 59752 189908 59764
rect 188764 59724 189908 59752
rect 188764 59712 188770 59724
rect 189902 59712 189908 59724
rect 189960 59712 189966 59764
rect 202690 59712 202696 59764
rect 202748 59752 202754 59764
rect 204806 59752 204812 59764
rect 202748 59724 204812 59752
rect 202748 59712 202754 59724
rect 204806 59712 204812 59724
rect 204864 59712 204870 59764
rect 209406 59712 209412 59764
rect 209464 59752 209470 59764
rect 209866 59752 209872 59764
rect 209464 59724 209872 59752
rect 209464 59712 209470 59724
rect 209866 59712 209872 59724
rect 209924 59712 209930 59764
rect 210786 59712 210792 59764
rect 210844 59752 210850 59764
rect 213178 59752 213184 59764
rect 210844 59724 213184 59752
rect 210844 59712 210850 59724
rect 213178 59712 213184 59724
rect 213236 59712 213242 59764
rect 216582 59712 216588 59764
rect 216640 59752 216646 59764
rect 218146 59752 218152 59764
rect 216640 59724 218152 59752
rect 216640 59712 216646 59724
rect 218146 59712 218152 59724
rect 218204 59712 218210 59764
rect 219250 59712 219256 59764
rect 219308 59752 219314 59764
rect 221458 59752 221464 59764
rect 219308 59724 221464 59752
rect 219308 59712 219314 59724
rect 221458 59712 221464 59724
rect 221516 59712 221522 59764
rect 238570 59712 238576 59764
rect 238628 59752 238634 59764
rect 240594 59752 240600 59764
rect 238628 59724 240600 59752
rect 238628 59712 238634 59724
rect 240594 59712 240600 59724
rect 240652 59712 240658 59764
rect 242710 59712 242716 59764
rect 242768 59752 242774 59764
rect 244734 59752 244740 59764
rect 242768 59724 244740 59752
rect 242768 59712 242774 59724
rect 244734 59712 244740 59724
rect 244792 59712 244798 59764
rect 248322 59712 248328 59764
rect 248380 59752 248386 59764
rect 249702 59752 249708 59764
rect 248380 59724 249708 59752
rect 248380 59712 248386 59724
rect 249702 59712 249708 59724
rect 249760 59712 249766 59764
rect 251818 59712 251824 59764
rect 251876 59752 251882 59764
rect 253198 59752 253204 59764
rect 251876 59724 253204 59752
rect 251876 59712 251882 59724
rect 253198 59712 253204 59724
rect 253256 59712 253262 59764
rect 267734 59712 267740 59764
rect 267792 59752 267798 59764
rect 269206 59752 269212 59764
rect 267792 59724 269212 59752
rect 267792 59712 267798 59724
rect 269206 59712 269212 59724
rect 269264 59712 269270 59764
rect 272702 59712 272708 59764
rect 272760 59752 272766 59764
rect 274726 59752 274732 59764
rect 272760 59724 274732 59752
rect 272760 59712 272766 59724
rect 274726 59712 274732 59724
rect 274784 59712 274790 59764
rect 276842 59712 276848 59764
rect 276900 59752 276906 59764
rect 278774 59752 278780 59764
rect 276900 59724 278780 59752
rect 276900 59712 276906 59724
rect 278774 59712 278780 59724
rect 278832 59712 278838 59764
rect 286778 59712 286784 59764
rect 286836 59752 286842 59764
rect 288434 59752 288440 59764
rect 286836 59724 288440 59752
rect 286836 59712 286842 59724
rect 288434 59712 288440 59724
rect 288492 59712 288498 59764
rect 291838 59712 291844 59764
rect 291896 59752 291902 59764
rect 294138 59752 294144 59764
rect 291896 59724 294144 59752
rect 291896 59712 291902 59724
rect 294138 59712 294144 59724
rect 294196 59712 294202 59764
rect 300118 59712 300124 59764
rect 300176 59752 300182 59764
rect 303062 59752 303068 59764
rect 300176 59724 303068 59752
rect 300176 59712 300182 59724
rect 303062 59712 303068 59724
rect 303120 59712 303126 59764
rect 303430 59712 303436 59764
rect 303488 59752 303494 59764
rect 305730 59752 305736 59764
rect 303488 59724 305736 59752
rect 303488 59712 303494 59724
rect 305730 59712 305736 59724
rect 305788 59712 305794 59764
rect 310698 59712 310704 59764
rect 310756 59752 310762 59764
rect 312538 59752 312544 59764
rect 310756 59724 312544 59752
rect 310756 59712 310762 59724
rect 312538 59712 312544 59724
rect 312596 59712 312602 59764
rect 318426 59712 318432 59764
rect 318484 59752 318490 59764
rect 320910 59752 320916 59764
rect 318484 59724 320916 59752
rect 318484 59712 318490 59724
rect 320910 59712 320916 59724
rect 320968 59712 320974 59764
rect 326706 59712 326712 59764
rect 326764 59752 326770 59764
rect 329098 59752 329104 59764
rect 326764 59724 329104 59752
rect 326764 59712 326770 59724
rect 329098 59712 329104 59724
rect 329156 59712 329162 59764
rect 330846 59712 330852 59764
rect 330904 59752 330910 59764
rect 331674 59752 331680 59764
rect 330904 59724 331680 59752
rect 330904 59712 330910 59724
rect 331674 59712 331680 59724
rect 331732 59712 331738 59764
rect 337562 59712 337568 59764
rect 337620 59752 337626 59764
rect 340322 59752 340328 59764
rect 337620 59724 340328 59752
rect 337620 59712 337626 59724
rect 340322 59712 340328 59724
rect 340380 59712 340386 59764
rect 345014 59712 345020 59764
rect 345072 59752 345078 59764
rect 347038 59752 347044 59764
rect 345072 59724 347044 59752
rect 345072 59712 345078 59724
rect 347038 59712 347044 59724
rect 347096 59712 347102 59764
rect 356698 59712 356704 59764
rect 356756 59752 356762 59764
rect 359642 59752 359648 59764
rect 356756 59724 359648 59752
rect 356756 59712 356762 59724
rect 359642 59712 359648 59724
rect 359700 59712 359706 59764
rect 360838 59712 360844 59764
rect 360896 59752 360902 59764
rect 363598 59752 363604 59764
rect 360896 59724 363604 59752
rect 360896 59712 360902 59724
rect 363598 59712 363604 59724
rect 363656 59712 363662 59764
rect 373810 59712 373816 59764
rect 373868 59752 373874 59764
rect 375466 59752 375472 59764
rect 373868 59724 375472 59752
rect 373868 59712 373874 59724
rect 375466 59712 375472 59724
rect 375524 59712 375530 59764
rect 379974 59712 379980 59764
rect 380032 59752 380038 59764
rect 380986 59752 380992 59764
rect 380032 59724 380992 59752
rect 380032 59712 380038 59724
rect 380986 59712 380992 59724
rect 381044 59712 381050 59764
rect 406562 59712 406568 59764
rect 406620 59752 406626 59764
rect 408494 59752 408500 59764
rect 406620 59724 408500 59752
rect 406620 59712 406626 59724
rect 408494 59712 408500 59724
rect 408552 59712 408558 59764
rect 409046 59712 409052 59764
rect 409104 59752 409110 59764
rect 410150 59752 410156 59764
rect 409104 59724 410156 59752
rect 409104 59712 409110 59724
rect 410150 59712 410156 59724
rect 410208 59712 410214 59764
rect 417602 59712 417608 59764
rect 417660 59752 417666 59764
rect 419626 59752 419632 59764
rect 417660 59724 419632 59752
rect 417660 59712 417666 59724
rect 419626 59712 419632 59724
rect 419684 59712 419690 59764
rect 422110 59712 422116 59764
rect 422168 59752 422174 59764
rect 423950 59752 423956 59764
rect 422168 59724 423956 59752
rect 422168 59712 422174 59724
rect 423950 59712 423956 59724
rect 424008 59712 424014 59764
rect 425698 59712 425704 59764
rect 425756 59752 425762 59764
rect 427998 59752 428004 59764
rect 425756 59724 428004 59752
rect 425756 59712 425762 59724
rect 427998 59712 428004 59724
rect 428056 59712 428062 59764
rect 429838 59712 429844 59764
rect 429896 59752 429902 59764
rect 432322 59752 432328 59764
rect 429896 59724 432328 59752
rect 429896 59712 429902 59724
rect 432322 59712 432328 59724
rect 432380 59712 432386 59764
rect 435818 59712 435824 59764
rect 435876 59752 435882 59764
rect 438302 59752 438308 59764
rect 435876 59724 438308 59752
rect 435876 59712 435882 59724
rect 438302 59712 438308 59724
rect 438360 59712 438366 59764
rect 442350 59712 442356 59764
rect 442408 59752 442414 59764
rect 445202 59752 445208 59764
rect 442408 59724 445208 59752
rect 442408 59712 442414 59724
rect 445202 59712 445208 59724
rect 445260 59712 445266 59764
rect 445662 59712 445668 59764
rect 445720 59752 445726 59764
rect 447778 59752 447784 59764
rect 445720 59724 447784 59752
rect 445720 59712 445726 59724
rect 447778 59712 447784 59724
rect 447836 59712 447842 59764
rect 456518 59712 456524 59764
rect 456576 59752 456582 59764
rect 458818 59752 458824 59764
rect 456576 59724 458824 59752
rect 456576 59712 456582 59724
rect 458818 59712 458824 59724
rect 458876 59712 458882 59764
rect 461486 59712 461492 59764
rect 461544 59752 461550 59764
rect 462958 59752 462964 59764
rect 461544 59724 462964 59752
rect 461544 59712 461550 59724
rect 462958 59712 462964 59724
rect 463016 59712 463022 59764
rect 158346 59644 158352 59696
rect 158404 59684 158410 59696
rect 159910 59684 159916 59696
rect 158404 59656 159916 59684
rect 158404 59644 158410 59656
rect 159910 59644 159916 59656
rect 159968 59644 159974 59696
rect 257338 59644 257344 59696
rect 257396 59684 257402 59696
rect 258074 59684 258080 59696
rect 257396 59656 258080 59684
rect 257396 59644 257402 59656
rect 258074 59644 258080 59656
rect 258132 59644 258138 59696
rect 301774 59644 301780 59696
rect 301832 59684 301838 59696
rect 304442 59684 304448 59696
rect 301832 59656 304448 59684
rect 301832 59644 301838 59656
rect 304442 59644 304448 59656
rect 304500 59644 304506 59696
rect 319254 59644 319260 59696
rect 319312 59684 319318 59696
rect 320174 59684 320180 59696
rect 319312 59656 320180 59684
rect 319312 59644 319318 59656
rect 320174 59644 320180 59656
rect 320232 59644 320238 59696
rect 320818 59644 320824 59696
rect 320876 59684 320882 59696
rect 322934 59684 322940 59696
rect 320876 59656 322940 59684
rect 320876 59644 320882 59656
rect 322934 59644 322940 59656
rect 322992 59644 322998 59696
rect 325050 59644 325056 59696
rect 325108 59684 325114 59696
rect 327718 59684 327724 59696
rect 325108 59656 327724 59684
rect 325108 59644 325114 59656
rect 327718 59644 327724 59656
rect 327776 59644 327782 59696
rect 330938 59644 330944 59696
rect 330996 59684 331002 59696
rect 333330 59684 333336 59696
rect 330996 59656 333336 59684
rect 330996 59644 331002 59656
rect 333330 59644 333336 59656
rect 333388 59644 333394 59696
rect 438210 59644 438216 59696
rect 438268 59684 438274 59696
rect 440878 59684 440884 59696
rect 438268 59656 440884 59684
rect 438268 59644 438274 59656
rect 440878 59644 440884 59656
rect 440936 59644 440942 59696
rect 454770 59644 454776 59696
rect 454828 59684 454834 59696
rect 457438 59684 457444 59696
rect 454828 59656 457444 59684
rect 454828 59644 454834 59656
rect 457438 59644 457444 59656
rect 457496 59644 457502 59696
rect 57238 59576 57244 59628
rect 57296 59616 57302 59628
rect 62666 59616 62672 59628
rect 57296 59588 62672 59616
rect 57296 59576 57302 59588
rect 62666 59576 62672 59588
rect 62724 59576 62730 59628
rect 75730 59576 75736 59628
rect 75788 59616 75794 59628
rect 77570 59616 77576 59628
rect 75788 59588 77576 59616
rect 75788 59576 75794 59588
rect 77570 59576 77576 59588
rect 77628 59576 77634 59628
rect 94498 59576 94504 59628
rect 94556 59616 94562 59628
rect 96706 59616 96712 59628
rect 94556 59588 96712 59616
rect 94556 59576 94562 59588
rect 96706 59576 96712 59588
rect 96764 59576 96770 59628
rect 102778 59576 102784 59628
rect 102836 59616 102842 59628
rect 105078 59616 105084 59628
rect 102836 59588 105084 59616
rect 102836 59576 102842 59588
rect 105078 59576 105084 59588
rect 105136 59576 105142 59628
rect 108298 59576 108304 59628
rect 108356 59616 108362 59628
rect 110874 59616 110880 59628
rect 108356 59588 110880 59616
rect 108356 59576 108362 59588
rect 110874 59576 110880 59588
rect 110932 59576 110938 59628
rect 117958 59576 117964 59628
rect 118016 59616 118022 59628
rect 119982 59616 119988 59628
rect 118016 59588 119988 59616
rect 118016 59576 118022 59588
rect 119982 59576 119988 59588
rect 120040 59576 120046 59628
rect 128998 59576 129004 59628
rect 129056 59616 129062 59628
rect 131666 59616 131672 59628
rect 129056 59588 131672 59616
rect 129056 59576 129062 59588
rect 131666 59576 131672 59588
rect 131724 59576 131730 59628
rect 131758 59576 131764 59628
rect 131816 59616 131822 59628
rect 134150 59616 134156 59628
rect 131816 59588 134156 59616
rect 131816 59576 131822 59588
rect 134150 59576 134156 59588
rect 134208 59576 134214 59628
rect 146202 59576 146208 59628
rect 146260 59616 146266 59628
rect 147490 59616 147496 59628
rect 146260 59588 147496 59616
rect 146260 59576 146266 59588
rect 147490 59576 147496 59588
rect 147548 59576 147554 59628
rect 179322 59576 179328 59628
rect 179380 59616 179386 59628
rect 180702 59616 180708 59628
rect 179380 59588 180708 59616
rect 179380 59576 179386 59588
rect 180702 59576 180708 59588
rect 180760 59576 180766 59628
rect 198550 59576 198556 59628
rect 198608 59616 198614 59628
rect 200666 59616 200672 59628
rect 198608 59588 200672 59616
rect 198608 59576 198614 59588
rect 200666 59576 200672 59588
rect 200724 59576 200730 59628
rect 227622 59576 227628 59628
rect 227680 59616 227686 59628
rect 228910 59616 228916 59628
rect 227680 59588 228916 59616
rect 227680 59576 227686 59588
rect 228910 59576 228916 59588
rect 228968 59576 228974 59628
rect 255958 59576 255964 59628
rect 256016 59616 256022 59628
rect 257246 59616 257252 59628
rect 256016 59588 257252 59616
rect 256016 59576 256022 59588
rect 257246 59576 257252 59588
rect 257304 59576 257310 59628
rect 258718 59576 258724 59628
rect 258776 59616 258782 59628
rect 260558 59616 260564 59628
rect 258776 59588 260564 59616
rect 258776 59576 258782 59588
rect 260558 59576 260564 59588
rect 260616 59576 260622 59628
rect 293494 59576 293500 59628
rect 293552 59616 293558 59628
rect 295518 59616 295524 59628
rect 293552 59588 295524 59616
rect 293552 59576 293558 59588
rect 295518 59576 295524 59588
rect 295576 59576 295582 59628
rect 296806 59576 296812 59628
rect 296864 59616 296870 59628
rect 298738 59616 298744 59628
rect 296864 59588 298744 59616
rect 296864 59576 296870 59588
rect 298738 59576 298744 59588
rect 298796 59576 298802 59628
rect 305914 59576 305920 59628
rect 305972 59616 305978 59628
rect 307018 59616 307024 59628
rect 305972 59588 307024 59616
rect 305972 59576 305978 59588
rect 307018 59576 307024 59588
rect 307076 59576 307082 59628
rect 316586 59576 316592 59628
rect 316644 59616 316650 59628
rect 318058 59616 318064 59628
rect 316644 59588 318064 59616
rect 316644 59576 316650 59588
rect 318058 59576 318064 59588
rect 318116 59576 318122 59628
rect 342346 59576 342352 59628
rect 342404 59616 342410 59628
rect 344462 59616 344468 59628
rect 342404 59588 344468 59616
rect 342404 59576 342410 59588
rect 344462 59576 344468 59588
rect 344520 59576 344526 59628
rect 353386 59576 353392 59628
rect 353444 59616 353450 59628
rect 354674 59616 354680 59628
rect 353444 59588 354680 59616
rect 353444 59576 353450 59588
rect 354674 59576 354680 59588
rect 354732 59576 354738 59628
rect 360102 59576 360108 59628
rect 360160 59616 360166 59628
rect 361022 59616 361028 59628
rect 360160 59588 361028 59616
rect 360160 59576 360166 59588
rect 361022 59576 361028 59588
rect 361080 59576 361086 59628
rect 369026 59576 369032 59628
rect 369084 59616 369090 59628
rect 369946 59616 369952 59628
rect 369084 59588 369952 59616
rect 369084 59576 369090 59588
rect 369946 59576 369952 59588
rect 370004 59576 370010 59628
rect 384114 59576 384120 59628
rect 384172 59616 384178 59628
rect 385402 59616 385408 59628
rect 384172 59588 385408 59616
rect 384172 59576 384178 59588
rect 385402 59576 385408 59588
rect 385460 59576 385466 59628
rect 393314 59576 393320 59628
rect 393372 59616 393378 59628
rect 394786 59616 394792 59628
rect 393372 59588 394792 59616
rect 393372 59576 393378 59588
rect 394786 59576 394792 59588
rect 394844 59576 394850 59628
rect 431770 59576 431776 59628
rect 431828 59616 431834 59628
rect 433702 59616 433708 59628
rect 431828 59588 433708 59616
rect 431828 59576 431834 59588
rect 433702 59576 433708 59588
rect 433760 59576 433766 59628
rect 450630 59576 450636 59628
rect 450688 59616 450694 59628
rect 451918 59616 451924 59628
rect 450688 59588 451924 59616
rect 450688 59576 450694 59588
rect 451918 59576 451924 59588
rect 451976 59576 451982 59628
rect 458174 59576 458180 59628
rect 458232 59616 458238 59628
rect 460198 59616 460204 59628
rect 458232 59588 460204 59616
rect 458232 59576 458238 59588
rect 460198 59576 460204 59588
rect 460256 59576 460262 59628
rect 146938 59508 146944 59560
rect 146996 59548 147002 59560
rect 149146 59548 149152 59560
rect 146996 59520 149152 59548
rect 146996 59508 147002 59520
rect 149146 59508 149152 59520
rect 149204 59508 149210 59560
rect 446398 59508 446404 59560
rect 446456 59548 446462 59560
rect 448514 59548 448520 59560
rect 446456 59520 448520 59548
rect 446456 59508 446462 59520
rect 448514 59508 448520 59520
rect 448572 59508 448578 59560
rect 115382 59440 115388 59492
rect 115440 59480 115446 59492
rect 117498 59480 117504 59492
rect 115440 59452 117504 59480
rect 115440 59440 115446 59452
rect 117498 59440 117504 59452
rect 117556 59440 117562 59492
rect 157058 59440 157064 59492
rect 157116 59480 157122 59492
rect 157334 59480 157340 59492
rect 157116 59452 157340 59480
rect 157116 59440 157122 59452
rect 157334 59440 157340 59452
rect 157392 59440 157398 59492
rect 176286 59440 176292 59492
rect 176344 59480 176350 59492
rect 178218 59480 178224 59492
rect 176344 59452 178224 59480
rect 176344 59440 176350 59452
rect 178218 59440 178224 59452
rect 178276 59440 178282 59492
rect 205266 59440 205272 59492
rect 205324 59480 205330 59492
rect 207290 59480 207296 59492
rect 205324 59452 207296 59480
rect 205324 59440 205330 59452
rect 207290 59440 207296 59452
rect 207348 59440 207354 59492
rect 215110 59440 215116 59492
rect 215168 59480 215174 59492
rect 215938 59480 215944 59492
rect 215168 59452 215944 59480
rect 215168 59440 215174 59452
rect 215938 59440 215944 59452
rect 215996 59440 216002 59492
rect 258994 59440 259000 59492
rect 259052 59480 259058 59492
rect 260558 59480 260564 59492
rect 259052 59452 260564 59480
rect 259052 59440 259058 59452
rect 260558 59440 260564 59452
rect 260616 59440 260622 59492
rect 282638 59440 282644 59492
rect 282696 59480 282702 59492
rect 284570 59480 284576 59492
rect 282696 59452 284576 59480
rect 282696 59440 282702 59452
rect 284570 59440 284576 59452
rect 284628 59440 284634 59492
rect 306742 59440 306748 59492
rect 306800 59480 306806 59492
rect 307754 59480 307760 59492
rect 306800 59452 307760 59480
rect 306800 59440 306806 59452
rect 307754 59440 307760 59452
rect 307812 59440 307818 59492
rect 321738 59440 321744 59492
rect 321796 59480 321802 59492
rect 323578 59480 323584 59492
rect 321796 59452 323584 59480
rect 321796 59440 321802 59452
rect 323578 59440 323584 59452
rect 323636 59440 323642 59492
rect 331766 59440 331772 59492
rect 331824 59480 331830 59492
rect 333238 59480 333244 59492
rect 331824 59452 333244 59480
rect 331824 59440 331830 59452
rect 333238 59440 333244 59452
rect 333296 59440 333302 59492
rect 333422 59440 333428 59492
rect 333480 59480 333486 59492
rect 336090 59480 336096 59492
rect 333480 59452 336096 59480
rect 333480 59440 333486 59452
rect 336090 59440 336096 59452
rect 336148 59440 336154 59492
rect 347498 59440 347504 59492
rect 347556 59480 347562 59492
rect 349982 59480 349988 59492
rect 347556 59452 349988 59480
rect 347556 59440 347562 59452
rect 349982 59440 349988 59452
rect 350040 59440 350046 59492
rect 362494 59440 362500 59492
rect 362552 59480 362558 59492
rect 364426 59480 364432 59492
rect 362552 59452 364432 59480
rect 362552 59440 362558 59452
rect 364426 59440 364432 59452
rect 364484 59440 364490 59492
rect 364794 59440 364800 59492
rect 364852 59480 364858 59492
rect 365714 59480 365720 59492
rect 364852 59452 365720 59480
rect 364852 59440 364858 59452
rect 365714 59440 365720 59452
rect 365772 59440 365778 59492
rect 366634 59440 366640 59492
rect 366692 59480 366698 59492
rect 368566 59480 368572 59492
rect 366692 59452 368572 59480
rect 366692 59440 366698 59452
rect 368566 59440 368572 59452
rect 368624 59440 368630 59492
rect 385770 59440 385776 59492
rect 385828 59480 385834 59492
rect 388162 59480 388168 59492
rect 385828 59452 388168 59480
rect 385828 59440 385834 59452
rect 388162 59440 388168 59452
rect 388220 59440 388226 59492
rect 419074 59440 419080 59492
rect 419132 59480 419138 59492
rect 421282 59480 421288 59492
rect 419132 59452 421288 59480
rect 419132 59440 419138 59452
rect 421282 59440 421288 59452
rect 421340 59440 421346 59492
rect 448146 59440 448152 59492
rect 448204 59480 448210 59492
rect 450722 59480 450728 59492
rect 448204 59452 450728 59480
rect 448204 59440 448210 59452
rect 450722 59440 450728 59452
rect 450780 59440 450786 59492
rect 452286 59440 452292 59492
rect 452344 59480 452350 59492
rect 454862 59480 454868 59492
rect 452344 59452 454868 59480
rect 452344 59440 452350 59452
rect 454862 59440 454868 59452
rect 454920 59440 454926 59492
rect 463142 59440 463148 59492
rect 463200 59480 463206 59492
rect 465902 59480 465908 59492
rect 463200 59452 465908 59480
rect 463200 59440 463206 59452
rect 465902 59440 465908 59452
rect 465960 59440 465966 59492
rect 3418 59372 3424 59424
rect 3476 59412 3482 59424
rect 57974 59412 57980 59424
rect 3476 59384 57980 59412
rect 3476 59372 3482 59384
rect 57974 59372 57980 59384
rect 58032 59372 58038 59424
rect 169478 59372 169484 59424
rect 169536 59412 169542 59424
rect 171594 59412 171600 59424
rect 169536 59384 171600 59412
rect 169536 59372 169542 59384
rect 171594 59372 171600 59384
rect 171652 59372 171658 59424
rect 194410 59372 194416 59424
rect 194468 59412 194474 59424
rect 196526 59412 196532 59424
rect 194468 59384 196532 59412
rect 194468 59372 194474 59384
rect 196526 59372 196532 59384
rect 196584 59372 196590 59424
rect 246666 59372 246672 59424
rect 246724 59412 246730 59424
rect 248874 59412 248880 59424
rect 246724 59384 248880 59412
rect 246724 59372 246730 59384
rect 248874 59372 248880 59384
rect 248932 59372 248938 59424
rect 135990 59304 135996 59356
rect 136048 59344 136054 59356
rect 137554 59344 137560 59356
rect 136048 59316 137560 59344
rect 136048 59304 136054 59316
rect 137554 59304 137560 59316
rect 137612 59304 137618 59356
rect 156966 59304 156972 59356
rect 157024 59344 157030 59356
rect 160094 59344 160100 59356
rect 157024 59316 160100 59344
rect 157024 59304 157030 59316
rect 160094 59304 160100 59316
rect 160152 59304 160158 59356
rect 451274 59304 451280 59356
rect 451332 59344 451338 59356
rect 453482 59344 453488 59356
rect 451332 59316 453488 59344
rect 451332 59304 451338 59316
rect 453482 59304 453488 59316
rect 453540 59304 453546 59356
rect 461486 59304 461492 59356
rect 461544 59344 461550 59356
rect 463142 59344 463148 59356
rect 461544 59316 463148 59344
rect 461544 59304 461550 59316
rect 463142 59304 463148 59316
rect 463200 59304 463206 59356
rect 350626 58964 350632 59016
rect 350684 59004 350690 59016
rect 352282 59004 352288 59016
rect 350684 58976 352288 59004
rect 350684 58964 350690 58976
rect 352282 58964 352288 58976
rect 352340 58964 352346 59016
rect 174538 58828 174544 58880
rect 174596 58868 174602 58880
rect 234614 58868 234620 58880
rect 174596 58840 234620 58868
rect 174596 58828 174602 58840
rect 234614 58828 234620 58840
rect 234672 58828 234678 58880
rect 235994 58828 236000 58880
rect 236052 58868 236058 58880
rect 280062 58868 280068 58880
rect 236052 58840 280068 58868
rect 236052 58828 236058 58840
rect 280062 58828 280068 58840
rect 280120 58828 280126 58880
rect 305638 58828 305644 58880
rect 305696 58868 305702 58880
rect 401502 58868 401508 58880
rect 305696 58840 401508 58868
rect 305696 58828 305702 58840
rect 401502 58828 401508 58840
rect 401560 58828 401566 58880
rect 186314 58760 186320 58812
rect 186372 58800 186378 58812
rect 268194 58800 268200 58812
rect 186372 58772 268200 58800
rect 186372 58760 186378 58772
rect 268194 58760 268200 58772
rect 268252 58760 268258 58812
rect 305822 58760 305828 58812
rect 305880 58800 305886 58812
rect 342254 58800 342260 58812
rect 305880 58772 342260 58800
rect 305880 58760 305886 58772
rect 342254 58760 342260 58772
rect 342312 58760 342318 58812
rect 351730 58760 351736 58812
rect 351788 58800 351794 58812
rect 538214 58800 538220 58812
rect 351788 58772 538220 58800
rect 351788 58760 351794 58772
rect 538214 58760 538220 58772
rect 538272 58760 538278 58812
rect 40034 58692 40040 58744
rect 40092 58732 40098 58744
rect 67542 58732 67548 58744
rect 40092 58704 67548 58732
rect 40092 58692 40098 58704
rect 67542 58692 67548 58704
rect 67600 58692 67606 58744
rect 81342 58692 81348 58744
rect 81400 58732 81406 58744
rect 89714 58732 89720 58744
rect 81400 58704 89720 58732
rect 81400 58692 81406 58704
rect 89714 58692 89720 58704
rect 89772 58692 89778 58744
rect 125594 58692 125600 58744
rect 125652 58732 125658 58744
rect 146202 58732 146208 58744
rect 125652 58704 146208 58732
rect 125652 58692 125658 58704
rect 146202 58692 146208 58704
rect 146260 58692 146266 58744
rect 194594 58692 194600 58744
rect 194652 58732 194658 58744
rect 376662 58732 376668 58744
rect 194652 58704 376668 58732
rect 194652 58692 194658 58704
rect 376662 58692 376668 58704
rect 376720 58692 376726 58744
rect 6914 58624 6920 58676
rect 6972 58664 6978 58676
rect 60642 58664 60648 58676
rect 6972 58636 60648 58664
rect 6972 58624 6978 58636
rect 60642 58624 60648 58636
rect 60700 58624 60706 58676
rect 88334 58624 88340 58676
rect 88392 58664 88398 58676
rect 131850 58664 131856 58676
rect 88392 58636 131856 58664
rect 88392 58624 88398 58636
rect 131850 58624 131856 58636
rect 131908 58624 131914 58676
rect 232774 58624 232780 58676
rect 232832 58664 232838 58676
rect 483014 58664 483020 58676
rect 232832 58636 483020 58664
rect 232832 58624 232838 58636
rect 483014 58624 483020 58636
rect 483072 58624 483078 58676
rect 142798 58488 142804 58540
rect 142856 58528 142862 58540
rect 144270 58528 144276 58540
rect 142856 58500 144276 58528
rect 142856 58488 142862 58500
rect 144270 58488 144276 58500
rect 144328 58488 144334 58540
rect 417602 58488 417608 58540
rect 417660 58528 417666 58540
rect 418430 58528 418436 58540
rect 417660 58500 418436 58528
rect 417660 58488 417666 58500
rect 418430 58488 418436 58500
rect 418488 58488 418494 58540
rect 222194 57468 222200 57520
rect 222252 57508 222258 57520
rect 277394 57508 277400 57520
rect 222252 57480 277400 57508
rect 222252 57468 222258 57480
rect 277394 57468 277400 57480
rect 277452 57468 277458 57520
rect 273254 57400 273260 57452
rect 273312 57440 273318 57452
rect 394694 57440 394700 57452
rect 273312 57412 394700 57440
rect 273312 57400 273318 57412
rect 394694 57400 394700 57412
rect 394752 57400 394758 57452
rect 165614 57332 165620 57384
rect 165672 57372 165678 57384
rect 262122 57372 262128 57384
rect 165672 57344 262128 57372
rect 165672 57332 165678 57344
rect 262122 57332 262128 57344
rect 262180 57332 262186 57384
rect 307754 57332 307760 57384
rect 307812 57372 307818 57384
rect 346394 57372 346400 57384
rect 307812 57344 346400 57372
rect 307812 57332 307818 57344
rect 346394 57332 346400 57344
rect 346452 57332 346458 57384
rect 354674 57332 354680 57384
rect 354732 57372 354738 57384
rect 545114 57372 545120 57384
rect 354732 57344 545120 57372
rect 354732 57332 354738 57344
rect 545114 57332 545120 57344
rect 545172 57332 545178 57384
rect 46934 57264 46940 57316
rect 46992 57304 46998 57316
rect 68922 57304 68928 57316
rect 46992 57276 68928 57304
rect 46992 57264 46998 57276
rect 68922 57264 68928 57276
rect 68980 57264 68986 57316
rect 88058 57264 88064 57316
rect 88116 57304 88122 57316
rect 118694 57304 118700 57316
rect 88116 57276 118700 57304
rect 88116 57264 88122 57276
rect 118694 57264 118700 57276
rect 118752 57264 118758 57316
rect 162854 57264 162860 57316
rect 162912 57304 162918 57316
rect 369486 57304 369492 57316
rect 162912 57276 369492 57304
rect 162912 57264 162918 57276
rect 369486 57264 369492 57276
rect 369544 57264 369550 57316
rect 32398 57196 32404 57248
rect 32456 57236 32462 57248
rect 91922 57236 91928 57248
rect 32456 57208 91928 57236
rect 32456 57196 32462 57208
rect 91922 57196 91928 57208
rect 91980 57196 91986 57248
rect 235258 57196 235264 57248
rect 235316 57236 235322 57248
rect 494054 57236 494060 57248
rect 235316 57208 494060 57236
rect 235316 57196 235322 57208
rect 494054 57196 494060 57208
rect 494112 57196 494118 57248
rect 218054 56040 218060 56092
rect 218112 56080 218118 56092
rect 278774 56080 278780 56092
rect 218112 56052 278780 56080
rect 218112 56040 218118 56052
rect 278774 56040 278780 56052
rect 278832 56040 278838 56092
rect 314654 56040 314660 56092
rect 314712 56080 314718 56092
rect 371234 56080 371240 56092
rect 314712 56052 371240 56080
rect 314712 56040 314718 56052
rect 371234 56040 371240 56052
rect 371292 56040 371298 56092
rect 168374 55972 168380 56024
rect 168432 56012 168438 56024
rect 262030 56012 262036 56024
rect 168432 55984 262036 56012
rect 168432 55972 168438 55984
rect 262030 55972 262036 55984
rect 262088 55972 262094 56024
rect 267734 55972 267740 56024
rect 267792 56012 267798 56024
rect 287054 56012 287060 56024
rect 267792 55984 287060 56012
rect 267792 55972 267798 55984
rect 287054 55972 287060 55984
rect 287112 55972 287118 56024
rect 320174 55972 320180 56024
rect 320232 56012 320238 56024
rect 398834 56012 398840 56024
rect 320232 55984 398840 56012
rect 320232 55972 320238 55984
rect 398834 55972 398840 55984
rect 398892 55972 398898 56024
rect 251174 55904 251180 55956
rect 251232 55944 251238 55956
rect 389450 55944 389456 55956
rect 251232 55916 389456 55944
rect 251232 55904 251238 55916
rect 389450 55904 389456 55916
rect 389508 55904 389514 55956
rect 448514 55904 448520 55956
rect 448572 55944 448578 55956
rect 489914 55944 489920 55956
rect 448572 55916 489920 55944
rect 448572 55904 448578 55916
rect 489914 55904 489920 55916
rect 489972 55904 489978 55956
rect 20714 55836 20720 55888
rect 20772 55876 20778 55888
rect 63402 55876 63408 55888
rect 20772 55848 63408 55876
rect 20772 55836 20778 55848
rect 63402 55836 63408 55848
rect 63460 55836 63466 55888
rect 87506 55836 87512 55888
rect 87564 55876 87570 55888
rect 121454 55876 121460 55888
rect 87564 55848 121460 55876
rect 87564 55836 87570 55848
rect 121454 55836 121460 55848
rect 121512 55836 121518 55888
rect 236914 55836 236920 55888
rect 236972 55876 236978 55888
rect 500954 55876 500960 55888
rect 236972 55848 500960 55876
rect 236972 55836 236978 55848
rect 500954 55836 500960 55848
rect 501012 55836 501018 55888
rect 190454 54680 190460 54732
rect 190512 54720 190518 54732
rect 271966 54720 271972 54732
rect 190512 54692 271972 54720
rect 190512 54680 190518 54692
rect 271966 54680 271972 54692
rect 272024 54680 272030 54732
rect 353938 54680 353944 54732
rect 353996 54720 354002 54732
rect 412818 54720 412824 54732
rect 353996 54692 412824 54720
rect 353996 54680 354002 54692
rect 412818 54680 412824 54692
rect 412876 54680 412882 54732
rect 198734 54612 198740 54664
rect 198792 54652 198798 54664
rect 379698 54652 379704 54664
rect 198792 54624 379704 54652
rect 198792 54612 198798 54624
rect 379698 54612 379704 54624
rect 379756 54612 379762 54664
rect 28994 54544 29000 54596
rect 29052 54584 29058 54596
rect 64322 54584 64328 54596
rect 29052 54556 64328 54584
rect 29052 54544 29058 54556
rect 64322 54544 64328 54556
rect 64380 54544 64386 54596
rect 226150 54544 226156 54596
rect 226208 54584 226214 54596
rect 465166 54584 465172 54596
rect 226208 54556 465172 54584
rect 226208 54544 226214 54556
rect 465166 54544 465172 54556
rect 465224 54544 465230 54596
rect 52454 54476 52460 54528
rect 52512 54516 52518 54528
rect 96062 54516 96068 54528
rect 52512 54488 96068 54516
rect 52512 54476 52518 54488
rect 96062 54476 96068 54488
rect 96120 54476 96126 54528
rect 106274 54476 106280 54528
rect 106332 54516 106338 54528
rect 136542 54516 136548 54528
rect 106332 54488 136548 54516
rect 106332 54476 106338 54488
rect 136542 54476 136548 54488
rect 136600 54476 136606 54528
rect 237282 54476 237288 54528
rect 237340 54516 237346 54528
rect 511994 54516 512000 54528
rect 237340 54488 512000 54516
rect 237340 54476 237346 54488
rect 511994 54476 512000 54488
rect 512052 54476 512058 54528
rect 129734 53252 129740 53304
rect 129792 53292 129798 53304
rect 253382 53292 253388 53304
rect 129792 53264 253388 53292
rect 129792 53252 129798 53264
rect 253382 53252 253388 53264
rect 253440 53252 253446 53304
rect 320818 53252 320824 53304
rect 320876 53292 320882 53304
rect 408494 53292 408500 53304
rect 320876 53264 408500 53292
rect 320876 53252 320882 53264
rect 408494 53252 408500 53264
rect 408552 53252 408558 53304
rect 170398 53184 170404 53236
rect 170456 53224 170462 53236
rect 372706 53224 372712 53236
rect 170456 53196 372712 53224
rect 170456 53184 170462 53196
rect 372706 53184 372712 53196
rect 372764 53184 372770 53236
rect 222010 53116 222016 53168
rect 222068 53156 222074 53168
rect 451274 53156 451280 53168
rect 222068 53128 451280 53156
rect 222068 53116 222074 53128
rect 451274 53116 451280 53128
rect 451332 53116 451338 53168
rect 451918 53116 451924 53168
rect 451976 53156 451982 53168
rect 503714 53156 503720 53168
rect 451976 53128 503720 53156
rect 451976 53116 451982 53128
rect 503714 53116 503720 53128
rect 503772 53116 503778 53168
rect 33134 53048 33140 53100
rect 33192 53088 33198 53100
rect 64138 53088 64144 53100
rect 33192 53060 64144 53088
rect 33192 53048 33198 53060
rect 64138 53048 64144 53060
rect 64196 53048 64202 53100
rect 69014 53048 69020 53100
rect 69072 53088 69078 53100
rect 100202 53088 100208 53100
rect 69072 53060 100208 53088
rect 69072 53048 69078 53060
rect 100202 53048 100208 53060
rect 100260 53048 100266 53100
rect 239950 53048 239956 53100
rect 240008 53088 240014 53100
rect 514754 53088 514760 53100
rect 240008 53060 514760 53088
rect 240008 53048 240014 53060
rect 514754 53048 514760 53060
rect 514812 53048 514818 53100
rect 240134 51892 240140 51944
rect 240192 51932 240198 51944
rect 282914 51932 282920 51944
rect 240192 51904 282920 51932
rect 240192 51892 240198 51904
rect 282914 51892 282920 51904
rect 282972 51892 282978 51944
rect 315298 51892 315304 51944
rect 315356 51932 315362 51944
rect 373994 51932 374000 51944
rect 315356 51904 374000 51932
rect 315356 51892 315362 51904
rect 373994 51892 374000 51904
rect 374052 51892 374058 51944
rect 136634 51824 136640 51876
rect 136692 51864 136698 51876
rect 254762 51864 254768 51876
rect 136692 51836 254768 51864
rect 136692 51824 136698 51836
rect 254762 51824 254768 51836
rect 254820 51824 254826 51876
rect 291194 51824 291200 51876
rect 291252 51864 291258 51876
rect 401594 51864 401600 51876
rect 291252 51836 401600 51864
rect 291252 51824 291258 51836
rect 401594 51824 401600 51836
rect 401652 51824 401658 51876
rect 190270 51756 190276 51808
rect 190328 51796 190334 51808
rect 316034 51796 316040 51808
rect 190328 51768 316040 51796
rect 190328 51756 190334 51768
rect 316034 51756 316040 51768
rect 316092 51756 316098 51808
rect 322934 51756 322940 51808
rect 322992 51796 322998 51808
rect 407114 51796 407120 51808
rect 322992 51768 407120 51796
rect 322992 51756 322998 51768
rect 407114 51756 407120 51768
rect 407172 51756 407178 51808
rect 44174 51688 44180 51740
rect 44232 51728 44238 51740
rect 66898 51728 66904 51740
rect 44232 51700 66904 51728
rect 44232 51688 44238 51700
rect 66898 51688 66904 51700
rect 66956 51688 66962 51740
rect 244182 51688 244188 51740
rect 244240 51728 244246 51740
rect 543734 51728 543740 51740
rect 244240 51700 543740 51728
rect 244240 51688 244246 51700
rect 543734 51688 543740 51700
rect 543792 51688 543798 51740
rect 183554 50532 183560 50584
rect 183612 50572 183618 50584
rect 270678 50572 270684 50584
rect 183612 50544 270684 50572
rect 183612 50532 183618 50544
rect 270678 50532 270684 50544
rect 270736 50532 270742 50584
rect 330570 50532 330576 50584
rect 330628 50572 330634 50584
rect 409966 50572 409972 50584
rect 330628 50544 409972 50572
rect 330628 50532 330634 50544
rect 409966 50532 409972 50544
rect 410024 50532 410030 50584
rect 169754 50464 169760 50516
rect 169812 50504 169818 50516
rect 372614 50504 372620 50516
rect 169812 50476 372620 50504
rect 169812 50464 169818 50476
rect 372614 50464 372620 50476
rect 372672 50464 372678 50516
rect 222102 50396 222108 50448
rect 222160 50436 222166 50448
rect 448514 50436 448520 50448
rect 222160 50408 448520 50436
rect 222160 50396 222166 50408
rect 448514 50396 448520 50408
rect 448572 50396 448578 50448
rect 48314 50328 48320 50380
rect 48372 50368 48378 50380
rect 95878 50368 95884 50380
rect 48372 50340 95884 50368
rect 48372 50328 48378 50340
rect 95878 50328 95884 50340
rect 95936 50328 95942 50380
rect 245470 50328 245476 50380
rect 245528 50368 245534 50380
rect 547874 50368 547880 50380
rect 245528 50340 547880 50368
rect 245528 50328 245534 50340
rect 547874 50328 547880 50340
rect 547932 50328 547938 50380
rect 172514 49172 172520 49224
rect 172572 49212 172578 49224
rect 268010 49212 268016 49224
rect 172572 49184 268016 49212
rect 172572 49172 172578 49184
rect 268010 49172 268016 49184
rect 268068 49172 268074 49224
rect 338758 49172 338764 49224
rect 338816 49212 338822 49224
rect 412726 49212 412732 49224
rect 338816 49184 412732 49212
rect 338816 49172 338822 49184
rect 412726 49172 412732 49184
rect 412784 49172 412790 49224
rect 186958 49104 186964 49156
rect 187016 49144 187022 49156
rect 376754 49144 376760 49156
rect 187016 49116 376760 49144
rect 187016 49104 187022 49116
rect 376754 49104 376760 49116
rect 376812 49104 376818 49156
rect 219250 49036 219256 49088
rect 219308 49076 219314 49088
rect 440326 49076 440332 49088
rect 219308 49048 440332 49076
rect 219308 49036 219314 49048
rect 440326 49036 440332 49048
rect 440384 49036 440390 49088
rect 14458 48968 14464 49020
rect 14516 49008 14522 49020
rect 87782 49008 87788 49020
rect 14516 48980 87788 49008
rect 14516 48968 14522 48980
rect 87782 48968 87788 48980
rect 87840 48968 87846 49020
rect 246850 48968 246856 49020
rect 246908 49008 246914 49020
rect 554774 49008 554780 49020
rect 246908 48980 554780 49008
rect 246908 48968 246914 48980
rect 554774 48968 554780 48980
rect 554832 48968 554838 49020
rect 176654 47744 176660 47796
rect 176712 47784 176718 47796
rect 267826 47784 267832 47796
rect 176712 47756 267832 47784
rect 176712 47744 176718 47756
rect 267826 47744 267832 47756
rect 267884 47744 267890 47796
rect 337470 47744 337476 47796
rect 337528 47784 337534 47796
rect 470594 47784 470600 47796
rect 337528 47756 470600 47784
rect 337528 47744 337534 47756
rect 470594 47744 470600 47756
rect 470652 47744 470658 47796
rect 214558 47676 214564 47728
rect 214616 47716 214622 47728
rect 383746 47716 383752 47728
rect 214616 47688 383752 47716
rect 214616 47676 214622 47688
rect 383746 47676 383752 47688
rect 383804 47676 383810 47728
rect 215110 47608 215116 47660
rect 215168 47648 215174 47660
rect 423674 47648 423680 47660
rect 215168 47620 423680 47648
rect 215168 47608 215174 47620
rect 423674 47608 423680 47620
rect 423732 47608 423738 47660
rect 17954 47540 17960 47592
rect 18012 47580 18018 47592
rect 89162 47580 89168 47592
rect 18012 47552 89168 47580
rect 18012 47540 18018 47552
rect 89162 47540 89168 47552
rect 89220 47540 89226 47592
rect 248322 47540 248328 47592
rect 248380 47580 248386 47592
rect 561674 47580 561680 47592
rect 248380 47552 561680 47580
rect 248380 47540 248386 47552
rect 561674 47540 561680 47552
rect 561732 47540 561738 47592
rect 193214 46384 193220 46436
rect 193272 46424 193278 46436
rect 271874 46424 271880 46436
rect 193272 46396 271880 46424
rect 193272 46384 193278 46396
rect 271874 46384 271880 46396
rect 271932 46384 271938 46436
rect 336090 46384 336096 46436
rect 336148 46424 336154 46436
rect 459554 46424 459560 46436
rect 336148 46396 459560 46424
rect 336148 46384 336154 46396
rect 459554 46384 459560 46396
rect 459612 46384 459618 46436
rect 206830 46316 206836 46368
rect 206888 46356 206894 46368
rect 387794 46356 387800 46368
rect 206888 46328 387800 46356
rect 206888 46316 206894 46328
rect 387794 46316 387800 46328
rect 387852 46316 387858 46368
rect 138014 46248 138020 46300
rect 138072 46288 138078 46300
rect 365714 46288 365720 46300
rect 138072 46260 365720 46288
rect 138072 46248 138078 46260
rect 365714 46248 365720 46260
rect 365772 46248 365778 46300
rect 27614 46180 27620 46232
rect 27672 46220 27678 46232
rect 90358 46220 90364 46232
rect 27672 46192 90364 46220
rect 27672 46180 27678 46192
rect 90358 46180 90364 46192
rect 90416 46180 90422 46232
rect 249610 46180 249616 46232
rect 249668 46220 249674 46232
rect 564526 46220 564532 46232
rect 249668 46192 564532 46220
rect 249668 46180 249674 46192
rect 564526 46180 564532 46192
rect 564584 46180 564590 46232
rect 316862 45024 316868 45076
rect 316920 45064 316926 45076
rect 378134 45064 378140 45076
rect 316920 45036 378140 45064
rect 316920 45024 316926 45036
rect 378134 45024 378140 45036
rect 378192 45024 378198 45076
rect 201494 44956 201500 45008
rect 201552 44996 201558 45008
rect 274726 44996 274732 45008
rect 201552 44968 274732 44996
rect 201552 44956 201558 44968
rect 274726 44956 274732 44968
rect 274784 44956 274790 45008
rect 333422 44956 333428 45008
rect 333480 44996 333486 45008
rect 448606 44996 448612 45008
rect 333480 44968 448612 44996
rect 333480 44956 333486 44968
rect 448606 44956 448612 44968
rect 448664 44956 448670 45008
rect 194318 44888 194324 44940
rect 194376 44928 194382 44940
rect 333974 44928 333980 44940
rect 194376 44900 333980 44928
rect 194376 44888 194382 44900
rect 333974 44888 333980 44900
rect 334032 44888 334038 44940
rect 352558 44888 352564 44940
rect 352616 44928 352622 44940
rect 414106 44928 414112 44940
rect 352616 44900 414112 44928
rect 352616 44888 352622 44900
rect 414106 44888 414112 44900
rect 414164 44888 414170 44940
rect 34514 44820 34520 44872
rect 34572 44860 34578 44872
rect 91738 44860 91744 44872
rect 34572 44832 91744 44860
rect 34572 44820 34578 44832
rect 91738 44820 91744 44832
rect 91796 44820 91802 44872
rect 158530 44820 158536 44872
rect 158588 44860 158594 44872
rect 182174 44860 182180 44872
rect 158588 44832 182180 44860
rect 158588 44820 158594 44832
rect 182174 44820 182180 44832
rect 182232 44820 182238 44872
rect 250990 44820 250996 44872
rect 251048 44860 251054 44872
rect 572714 44860 572720 44872
rect 251048 44832 572720 44860
rect 251048 44820 251054 44832
rect 572714 44820 572720 44832
rect 572772 44820 572778 44872
rect 177850 43596 177856 43648
rect 177908 43636 177914 43648
rect 263594 43636 263600 43648
rect 177908 43608 263600 43636
rect 177908 43596 177914 43608
rect 263594 43596 263600 43608
rect 263652 43596 263658 43648
rect 322934 43596 322940 43648
rect 322992 43636 322998 43648
rect 408770 43636 408776 43648
rect 322992 43608 408776 43636
rect 322992 43596 322998 43608
rect 408770 43596 408776 43608
rect 408828 43596 408834 43648
rect 194502 43528 194508 43580
rect 194560 43568 194566 43580
rect 331214 43568 331220 43580
rect 194560 43540 331220 43568
rect 194560 43528 194566 43540
rect 331214 43528 331220 43540
rect 331272 43528 331278 43580
rect 348602 43528 348608 43580
rect 348660 43568 348666 43580
rect 516134 43568 516140 43580
rect 348660 43540 516140 43568
rect 348660 43528 348666 43540
rect 516134 43528 516140 43540
rect 516192 43528 516198 43580
rect 205634 43460 205640 43512
rect 205692 43500 205698 43512
rect 380986 43500 380992 43512
rect 205692 43472 380992 43500
rect 205692 43460 205698 43472
rect 380986 43460 380992 43472
rect 381044 43460 381050 43512
rect 9674 43392 9680 43444
rect 9732 43432 9738 43444
rect 113818 43432 113824 43444
rect 9732 43404 113824 43432
rect 9732 43392 9738 43404
rect 113818 43392 113824 43404
rect 113876 43392 113882 43444
rect 217870 43392 217876 43444
rect 217928 43432 217934 43444
rect 430574 43432 430580 43444
rect 217928 43404 430580 43432
rect 217928 43392 217934 43404
rect 430574 43392 430580 43404
rect 430632 43392 430638 43444
rect 259454 42236 259460 42288
rect 259512 42276 259518 42288
rect 393406 42276 393412 42288
rect 259512 42248 393412 42276
rect 259512 42236 259518 42248
rect 393406 42236 393412 42248
rect 393464 42236 393470 42288
rect 201310 42168 201316 42220
rect 201368 42208 201374 42220
rect 362954 42208 362960 42220
rect 201368 42180 362960 42208
rect 201368 42168 201374 42180
rect 362954 42168 362960 42180
rect 363012 42168 363018 42220
rect 186130 42100 186136 42152
rect 186188 42140 186194 42152
rect 295334 42140 295340 42152
rect 186188 42112 295340 42140
rect 186188 42100 186194 42112
rect 295334 42100 295340 42112
rect 295392 42100 295398 42152
rect 352834 42100 352840 42152
rect 352892 42140 352898 42152
rect 534074 42140 534080 42152
rect 352892 42112 534080 42140
rect 352892 42100 352898 42112
rect 534074 42100 534080 42112
rect 534132 42100 534138 42152
rect 49694 42032 49700 42084
rect 49752 42072 49758 42084
rect 122098 42072 122104 42084
rect 49752 42044 122104 42072
rect 49752 42032 49758 42044
rect 122098 42032 122104 42044
rect 122156 42032 122162 42084
rect 224770 42032 224776 42084
rect 224828 42072 224834 42084
rect 462314 42072 462320 42084
rect 224828 42044 462320 42072
rect 224828 42032 224834 42044
rect 462314 42032 462320 42044
rect 462372 42032 462378 42084
rect 158714 40876 158720 40928
rect 158772 40916 158778 40928
rect 258902 40916 258908 40928
rect 158772 40888 258908 40916
rect 158772 40876 158778 40888
rect 258902 40876 258908 40888
rect 258960 40876 258966 40928
rect 319622 40876 319628 40928
rect 319680 40916 319686 40928
rect 389174 40916 389180 40928
rect 319680 40888 389180 40916
rect 319680 40876 319686 40888
rect 389174 40876 389180 40888
rect 389232 40876 389238 40928
rect 244274 40808 244280 40860
rect 244332 40848 244338 40860
rect 390554 40848 390560 40860
rect 244332 40820 390560 40848
rect 244332 40808 244338 40820
rect 390554 40808 390560 40820
rect 390612 40808 390618 40860
rect 190086 40740 190092 40792
rect 190144 40780 190150 40792
rect 313274 40780 313280 40792
rect 190144 40752 313280 40780
rect 190144 40740 190150 40752
rect 313274 40740 313280 40752
rect 313332 40740 313338 40792
rect 344462 40740 344468 40792
rect 344520 40780 344526 40792
rect 495434 40780 495440 40792
rect 344520 40752 495440 40780
rect 344520 40740 344526 40752
rect 495434 40740 495440 40752
rect 495492 40740 495498 40792
rect 205450 40672 205456 40724
rect 205508 40712 205514 40724
rect 376754 40712 376760 40724
rect 205508 40684 376760 40712
rect 205508 40672 205514 40684
rect 376754 40672 376760 40684
rect 376812 40672 376818 40724
rect 456058 40672 456064 40724
rect 456116 40712 456122 40724
rect 521654 40712 521660 40724
rect 456116 40684 521660 40712
rect 456116 40672 456122 40684
rect 521654 40672 521660 40684
rect 521712 40672 521718 40724
rect 326338 39516 326344 39568
rect 326396 39556 326402 39568
rect 420914 39556 420920 39568
rect 326396 39528 420920 39556
rect 326396 39516 326402 39528
rect 420914 39516 420920 39528
rect 420972 39516 420978 39568
rect 188890 39448 188896 39500
rect 188948 39488 188954 39500
rect 309134 39488 309140 39500
rect 188948 39460 309140 39488
rect 188948 39448 188954 39460
rect 309134 39448 309140 39460
rect 309192 39448 309198 39500
rect 309778 39448 309784 39500
rect 309836 39488 309842 39500
rect 405826 39488 405832 39500
rect 309836 39460 405832 39488
rect 309836 39448 309842 39460
rect 405826 39448 405832 39460
rect 405884 39448 405890 39500
rect 204162 39380 204168 39432
rect 204220 39420 204226 39432
rect 374086 39420 374092 39432
rect 204220 39392 374092 39420
rect 204220 39380 204226 39392
rect 374086 39380 374092 39392
rect 374144 39380 374150 39432
rect 449158 39380 449164 39432
rect 449216 39420 449222 39432
rect 492674 39420 492680 39432
rect 449216 39392 492680 39420
rect 449216 39380 449222 39392
rect 492674 39380 492680 39392
rect 492732 39380 492738 39432
rect 227622 39312 227628 39364
rect 227680 39352 227686 39364
rect 473354 39352 473360 39364
rect 227680 39324 473360 39352
rect 227680 39312 227686 39324
rect 473354 39312 473360 39324
rect 473412 39312 473418 39364
rect 278038 38088 278044 38140
rect 278096 38128 278102 38140
rect 397546 38128 397552 38140
rect 278096 38100 397552 38128
rect 278096 38088 278102 38100
rect 397546 38088 397552 38100
rect 397604 38088 397610 38140
rect 202690 38020 202696 38072
rect 202748 38060 202754 38072
rect 369854 38060 369860 38072
rect 202748 38032 369860 38060
rect 202748 38020 202754 38032
rect 369854 38020 369860 38032
rect 369912 38020 369918 38072
rect 188706 37952 188712 38004
rect 188764 37992 188770 38004
rect 306374 37992 306380 38004
rect 188764 37964 306380 37992
rect 188764 37952 188770 37964
rect 306374 37952 306380 37964
rect 306432 37952 306438 38004
rect 354030 37952 354036 38004
rect 354088 37992 354094 38004
rect 540974 37992 540980 38004
rect 354088 37964 540980 37992
rect 354088 37952 354094 37964
rect 540974 37952 540980 37964
rect 541032 37952 541038 38004
rect 225966 37884 225972 37936
rect 226024 37924 226030 37936
rect 469214 37924 469220 37936
rect 226024 37896 469220 37924
rect 226024 37884 226030 37896
rect 469214 37884 469220 37896
rect 469272 37884 469278 37936
rect 266354 36728 266360 36780
rect 266412 36768 266418 36780
rect 396166 36768 396172 36780
rect 266412 36740 396172 36768
rect 266412 36728 266418 36740
rect 396166 36728 396172 36740
rect 396224 36728 396230 36780
rect 202506 36660 202512 36712
rect 202564 36700 202570 36712
rect 365714 36700 365720 36712
rect 202564 36672 365720 36700
rect 202564 36660 202570 36672
rect 365714 36660 365720 36672
rect 365772 36660 365778 36712
rect 187602 36592 187608 36644
rect 187660 36632 187666 36644
rect 302234 36632 302240 36644
rect 187660 36604 302240 36632
rect 187660 36592 187666 36604
rect 302234 36592 302240 36604
rect 302292 36592 302298 36644
rect 352650 36592 352656 36644
rect 352708 36632 352714 36644
rect 531314 36632 531320 36644
rect 352708 36604 531320 36632
rect 352708 36592 352714 36604
rect 531314 36592 531320 36604
rect 531372 36592 531378 36644
rect 223482 36524 223488 36576
rect 223540 36564 223546 36576
rect 455414 36564 455420 36576
rect 223540 36536 455420 36564
rect 223540 36524 223546 36536
rect 455414 36524 455420 36536
rect 455472 36524 455478 36576
rect 262214 35368 262220 35420
rect 262272 35408 262278 35420
rect 394694 35408 394700 35420
rect 262272 35380 394700 35408
rect 262272 35368 262278 35380
rect 394694 35368 394700 35380
rect 394752 35368 394758 35420
rect 201126 35300 201132 35352
rect 201184 35340 201190 35352
rect 358814 35340 358820 35352
rect 201184 35312 358820 35340
rect 201184 35300 201190 35312
rect 358814 35300 358820 35312
rect 358872 35300 358878 35352
rect 185946 35232 185952 35284
rect 186004 35272 186010 35284
rect 299474 35272 299480 35284
rect 186004 35244 299480 35272
rect 186004 35232 186010 35244
rect 299474 35232 299480 35244
rect 299532 35232 299538 35284
rect 351178 35232 351184 35284
rect 351236 35272 351242 35284
rect 527174 35272 527180 35284
rect 351236 35244 527180 35272
rect 351236 35232 351242 35244
rect 527174 35232 527180 35244
rect 527232 35232 527238 35284
rect 220722 35164 220728 35216
rect 220780 35204 220786 35216
rect 444374 35204 444380 35216
rect 220780 35176 444380 35204
rect 220780 35164 220786 35176
rect 444374 35164 444380 35176
rect 444432 35164 444438 35216
rect 184750 33940 184756 33992
rect 184808 33980 184814 33992
rect 292574 33980 292580 33992
rect 184808 33952 292580 33980
rect 184808 33940 184814 33952
rect 292574 33940 292580 33952
rect 292632 33940 292638 33992
rect 336090 33940 336096 33992
rect 336148 33980 336154 33992
rect 411254 33980 411260 33992
rect 336148 33952 411260 33980
rect 336148 33940 336154 33952
rect 411254 33940 411260 33952
rect 411312 33940 411318 33992
rect 216674 33872 216680 33924
rect 216732 33912 216738 33924
rect 383930 33912 383936 33924
rect 216732 33884 383936 33912
rect 216732 33872 216738 33884
rect 383930 33872 383936 33884
rect 383988 33872 383994 33924
rect 197170 33804 197176 33856
rect 197228 33844 197234 33856
rect 340874 33844 340880 33856
rect 197228 33816 340880 33844
rect 197228 33804 197234 33816
rect 340874 33804 340880 33816
rect 340932 33804 340938 33856
rect 349982 33804 349988 33856
rect 350040 33844 350046 33856
rect 520274 33844 520280 33856
rect 350040 33816 520280 33844
rect 350040 33804 350046 33816
rect 520274 33804 520280 33816
rect 520332 33804 520338 33856
rect 92474 33736 92480 33788
rect 92532 33776 92538 33788
rect 131758 33776 131764 33788
rect 92532 33748 131764 33776
rect 92532 33736 92538 33748
rect 131758 33736 131764 33748
rect 131816 33736 131822 33788
rect 219066 33736 219072 33788
rect 219124 33776 219130 33788
rect 437474 33776 437480 33788
rect 219124 33748 437480 33776
rect 219124 33736 219130 33748
rect 437474 33736 437480 33748
rect 437532 33736 437538 33788
rect 177666 32580 177672 32632
rect 177724 32620 177730 32632
rect 259546 32620 259552 32632
rect 177724 32592 259552 32620
rect 177724 32580 177730 32592
rect 259546 32580 259552 32592
rect 259604 32580 259610 32632
rect 320910 32580 320916 32632
rect 320968 32620 320974 32632
rect 396074 32620 396080 32632
rect 320968 32592 396080 32620
rect 320968 32580 320974 32592
rect 396074 32580 396080 32592
rect 396132 32580 396138 32632
rect 193030 32512 193036 32564
rect 193088 32552 193094 32564
rect 324314 32552 324320 32564
rect 193088 32524 324320 32552
rect 193088 32512 193094 32524
rect 324314 32512 324320 32524
rect 324372 32512 324378 32564
rect 344278 32512 344284 32564
rect 344336 32552 344342 32564
rect 498194 32552 498200 32564
rect 344336 32524 498200 32552
rect 344336 32512 344342 32524
rect 498194 32512 498200 32524
rect 498252 32512 498258 32564
rect 214926 32444 214932 32496
rect 214984 32484 214990 32496
rect 419534 32484 419540 32496
rect 214984 32456 419540 32484
rect 214984 32444 214990 32456
rect 419534 32444 419540 32456
rect 419592 32444 419598 32496
rect 70394 32376 70400 32428
rect 70452 32416 70458 32428
rect 127802 32416 127808 32428
rect 70452 32388 127808 32416
rect 70452 32376 70458 32388
rect 127802 32376 127808 32388
rect 127860 32376 127866 32428
rect 142154 32376 142160 32428
rect 142212 32416 142218 32428
rect 367094 32416 367100 32428
rect 142212 32388 367100 32416
rect 142212 32376 142218 32388
rect 367094 32376 367100 32388
rect 367152 32376 367158 32428
rect 457622 32376 457628 32428
rect 457680 32416 457686 32428
rect 528554 32416 528560 32428
rect 457680 32388 528560 32416
rect 457680 32376 457686 32388
rect 528554 32376 528560 32388
rect 528612 32376 528618 32428
rect 147674 31220 147680 31272
rect 147732 31260 147738 31272
rect 257522 31260 257528 31272
rect 147732 31232 257528 31260
rect 147732 31220 147738 31232
rect 257522 31220 257528 31232
rect 257580 31220 257586 31272
rect 343634 31220 343640 31272
rect 343692 31260 343698 31272
rect 414290 31260 414296 31272
rect 343692 31232 414296 31260
rect 343692 31220 343698 31232
rect 414290 31220 414296 31232
rect 414348 31220 414354 31272
rect 201586 31152 201592 31204
rect 201644 31192 201650 31204
rect 380894 31192 380900 31204
rect 201644 31164 380900 31192
rect 201644 31152 201650 31164
rect 380894 31152 380900 31164
rect 380952 31152 380958 31204
rect 217686 31084 217692 31136
rect 217744 31124 217750 31136
rect 433334 31124 433340 31136
rect 217744 31096 433340 31124
rect 217744 31084 217750 31096
rect 433334 31084 433340 31096
rect 433392 31084 433398 31136
rect 63494 31016 63500 31068
rect 63552 31056 63558 31068
rect 125042 31056 125048 31068
rect 63552 31028 125048 31056
rect 63552 31016 63558 31028
rect 125042 31016 125048 31028
rect 125100 31016 125106 31068
rect 175182 31016 175188 31068
rect 175240 31056 175246 31068
rect 249794 31056 249800 31068
rect 175240 31028 249800 31056
rect 175240 31016 175246 31028
rect 249794 31016 249800 31028
rect 249852 31016 249858 31068
rect 251082 31016 251088 31068
rect 251140 31056 251146 31068
rect 575474 31056 575480 31068
rect 251140 31028 575480 31056
rect 251140 31016 251146 31028
rect 575474 31016 575480 31028
rect 575532 31016 575538 31068
rect 309870 29860 309876 29912
rect 309928 29900 309934 29912
rect 349154 29900 349160 29912
rect 309928 29872 349160 29900
rect 309928 29860 309934 29872
rect 349154 29860 349160 29872
rect 349212 29860 349218 29912
rect 229094 29792 229100 29844
rect 229152 29832 229158 29844
rect 280154 29832 280160 29844
rect 229152 29804 280160 29832
rect 229152 29792 229158 29804
rect 280154 29792 280160 29804
rect 280212 29792 280218 29844
rect 319438 29792 319444 29844
rect 319496 29832 319502 29844
rect 391934 29832 391940 29844
rect 319496 29804 391940 29832
rect 319496 29792 319502 29804
rect 391934 29792 391940 29804
rect 391992 29792 391998 29844
rect 140774 29724 140780 29776
rect 140832 29764 140838 29776
rect 254578 29764 254584 29776
rect 140832 29736 254584 29764
rect 140832 29724 140838 29736
rect 254578 29724 254584 29736
rect 254636 29724 254642 29776
rect 269114 29724 269120 29776
rect 269172 29764 269178 29776
rect 396350 29764 396356 29776
rect 269172 29736 396356 29764
rect 269172 29724 269178 29736
rect 396350 29724 396356 29736
rect 396408 29724 396414 29776
rect 191742 29656 191748 29708
rect 191800 29696 191806 29708
rect 320174 29696 320180 29708
rect 191800 29668 320180 29696
rect 191800 29656 191806 29668
rect 320174 29656 320180 29668
rect 320232 29656 320238 29708
rect 358170 29656 358176 29708
rect 358228 29696 358234 29708
rect 416866 29696 416872 29708
rect 358228 29668 416872 29696
rect 358228 29656 358234 29668
rect 416866 29656 416872 29668
rect 416924 29656 416930 29708
rect 60734 29588 60740 29640
rect 60792 29628 60798 29640
rect 124858 29628 124864 29640
rect 60792 29600 124864 29628
rect 60792 29588 60798 29600
rect 124858 29588 124864 29600
rect 124916 29588 124922 29640
rect 249426 29588 249432 29640
rect 249484 29628 249490 29640
rect 568574 29628 568580 29640
rect 249484 29600 568580 29628
rect 249484 29588 249490 29600
rect 568574 29588 568580 29600
rect 568632 29588 568638 29640
rect 311894 28432 311900 28484
rect 311952 28472 311958 28484
rect 405734 28472 405740 28484
rect 311952 28444 405740 28472
rect 311952 28432 311958 28444
rect 405734 28432 405740 28444
rect 405792 28432 405798 28484
rect 216582 28364 216588 28416
rect 216640 28404 216646 28416
rect 426434 28404 426440 28416
rect 216640 28376 426440 28404
rect 216640 28364 216646 28376
rect 426434 28364 426440 28376
rect 426492 28364 426498 28416
rect 126974 28296 126980 28348
rect 127032 28336 127038 28348
rect 363046 28336 363052 28348
rect 127032 28308 363052 28336
rect 127032 28296 127038 28308
rect 363046 28296 363052 28308
rect 363104 28296 363110 28348
rect 56594 28228 56600 28280
rect 56652 28268 56658 28280
rect 123662 28268 123668 28280
rect 56652 28240 123668 28268
rect 56652 28228 56658 28240
rect 123662 28228 123668 28240
rect 123720 28228 123726 28280
rect 173618 28228 173624 28280
rect 173676 28268 173682 28280
rect 245654 28268 245660 28280
rect 173676 28240 245660 28268
rect 173676 28228 173682 28240
rect 245654 28228 245660 28240
rect 245712 28228 245718 28280
rect 246666 28228 246672 28280
rect 246724 28268 246730 28280
rect 557534 28268 557540 28280
rect 246724 28240 557540 28268
rect 246724 28228 246730 28240
rect 557534 28228 557540 28240
rect 557592 28228 557598 28280
rect 338850 27072 338856 27124
rect 338908 27112 338914 27124
rect 473446 27112 473452 27124
rect 338908 27084 473452 27112
rect 338908 27072 338914 27084
rect 473446 27072 473452 27084
rect 473504 27072 473510 27124
rect 191834 27004 191840 27056
rect 191892 27044 191898 27056
rect 378226 27044 378232 27056
rect 191892 27016 378232 27044
rect 191892 27004 191898 27016
rect 378226 27004 378232 27016
rect 378284 27004 378290 27056
rect 212442 26936 212448 26988
rect 212500 26976 212506 26988
rect 408494 26976 408500 26988
rect 212500 26948 408500 26976
rect 212500 26936 212506 26948
rect 408494 26936 408500 26948
rect 408552 26936 408558 26988
rect 52546 26868 52552 26920
rect 52604 26908 52610 26920
rect 123478 26908 123484 26920
rect 52604 26880 123484 26908
rect 52604 26868 52610 26880
rect 123478 26868 123484 26880
rect 123536 26868 123542 26920
rect 173802 26868 173808 26920
rect 173860 26908 173866 26920
rect 242894 26908 242900 26920
rect 173860 26880 242900 26908
rect 173860 26868 173866 26880
rect 242894 26868 242900 26880
rect 242952 26868 242958 26920
rect 245286 26868 245292 26920
rect 245344 26908 245350 26920
rect 550634 26908 550640 26920
rect 245344 26880 550640 26908
rect 245344 26868 245350 26880
rect 550634 26868 550640 26880
rect 550692 26868 550698 26920
rect 172422 25712 172428 25764
rect 172480 25752 172486 25764
rect 238754 25752 238760 25764
rect 172480 25724 238760 25752
rect 172480 25712 172486 25724
rect 238754 25712 238760 25724
rect 238812 25712 238818 25764
rect 337378 25712 337384 25764
rect 337436 25752 337442 25764
rect 466454 25752 466460 25764
rect 337436 25724 466460 25752
rect 337436 25712 337442 25724
rect 466454 25712 466460 25724
rect 466512 25712 466518 25764
rect 210970 25644 210976 25696
rect 211028 25684 211034 25696
rect 401594 25684 401600 25696
rect 211028 25656 401600 25684
rect 211028 25644 211034 25656
rect 401594 25644 401600 25656
rect 401652 25644 401658 25696
rect 131114 25576 131120 25628
rect 131172 25616 131178 25628
rect 364426 25616 364432 25628
rect 131172 25588 364432 25616
rect 131172 25576 131178 25588
rect 364426 25576 364432 25588
rect 364484 25576 364490 25628
rect 44266 25508 44272 25560
rect 44324 25548 44330 25560
rect 94498 25548 94504 25560
rect 44324 25520 94504 25548
rect 44324 25508 44330 25520
rect 94498 25508 94504 25520
rect 94556 25508 94562 25560
rect 238570 25508 238576 25560
rect 238628 25548 238634 25560
rect 523034 25548 523040 25560
rect 238628 25520 523040 25548
rect 238628 25508 238634 25520
rect 523034 25508 523040 25520
rect 523092 25508 523098 25560
rect 318058 24284 318064 24336
rect 318116 24324 318122 24336
rect 385034 24324 385040 24336
rect 318116 24296 385040 24324
rect 318116 24284 318122 24296
rect 385034 24284 385040 24296
rect 385092 24284 385098 24336
rect 127066 24216 127072 24268
rect 127124 24256 127130 24268
rect 251818 24256 251824 24268
rect 127124 24228 251824 24256
rect 127124 24216 127130 24228
rect 251818 24216 251824 24228
rect 251876 24216 251882 24268
rect 335998 24216 336004 24268
rect 336056 24256 336062 24268
rect 463694 24256 463700 24268
rect 336056 24228 463700 24256
rect 336056 24216 336062 24228
rect 463694 24216 463700 24228
rect 463752 24216 463758 24268
rect 195882 24148 195888 24200
rect 195940 24188 195946 24200
rect 338114 24188 338120 24200
rect 195940 24160 338120 24188
rect 195940 24148 195946 24160
rect 338114 24148 338120 24160
rect 338172 24148 338178 24200
rect 22094 24080 22100 24132
rect 22152 24120 22158 24132
rect 88978 24120 88984 24132
rect 22152 24092 88984 24120
rect 22152 24080 22158 24092
rect 88978 24080 88984 24092
rect 89036 24080 89042 24132
rect 235902 24080 235908 24132
rect 235960 24120 235966 24132
rect 507854 24120 507860 24132
rect 235960 24092 507860 24120
rect 235960 24080 235966 24092
rect 507854 24080 507860 24092
rect 507912 24080 507918 24132
rect 316678 22924 316684 22976
rect 316736 22964 316742 22976
rect 382274 22964 382280 22976
rect 316736 22936 382280 22964
rect 316736 22924 316742 22936
rect 382274 22924 382280 22936
rect 382332 22924 382338 22976
rect 133874 22856 133880 22908
rect 133932 22896 133938 22908
rect 253198 22896 253204 22908
rect 133932 22868 253204 22896
rect 133932 22856 133938 22868
rect 253198 22856 253204 22868
rect 253256 22856 253262 22908
rect 329834 22856 329840 22908
rect 329892 22896 329898 22908
rect 410150 22896 410156 22908
rect 329892 22868 410156 22896
rect 329892 22856 329898 22868
rect 410150 22856 410156 22868
rect 410208 22856 410214 22908
rect 192846 22788 192852 22840
rect 192904 22828 192910 22840
rect 327074 22828 327080 22840
rect 192904 22800 327080 22828
rect 192904 22788 192910 22800
rect 327074 22788 327080 22800
rect 327132 22788 327138 22840
rect 332042 22788 332048 22840
rect 332100 22828 332106 22840
rect 445754 22828 445760 22840
rect 332100 22800 445760 22828
rect 332100 22788 332106 22800
rect 445754 22788 445760 22800
rect 445812 22788 445818 22840
rect 77294 22720 77300 22772
rect 77352 22760 77358 22772
rect 102962 22760 102968 22772
rect 77352 22732 102968 22760
rect 77352 22720 77358 22732
rect 102962 22720 102968 22732
rect 103020 22720 103026 22772
rect 234246 22720 234252 22772
rect 234304 22760 234310 22772
rect 505094 22760 505100 22772
rect 234304 22732 505100 22760
rect 234304 22720 234310 22732
rect 505094 22720 505100 22732
rect 505152 22720 505158 22772
rect 280154 21564 280160 21616
rect 280212 21604 280218 21616
rect 398926 21604 398932 21616
rect 280212 21576 398932 21604
rect 280212 21564 280218 21576
rect 398926 21564 398932 21576
rect 398984 21564 398990 21616
rect 151814 21496 151820 21548
rect 151872 21536 151878 21548
rect 257338 21536 257344 21548
rect 151872 21508 257344 21536
rect 151872 21496 151878 21508
rect 257338 21496 257344 21508
rect 257396 21496 257402 21548
rect 334618 21496 334624 21548
rect 334676 21536 334682 21548
rect 456886 21536 456892 21548
rect 334676 21508 456892 21536
rect 334676 21496 334682 21508
rect 456886 21496 456892 21508
rect 456944 21496 456950 21548
rect 208302 21428 208308 21480
rect 208360 21468 208366 21480
rect 390554 21468 390560 21480
rect 208360 21440 390560 21468
rect 208360 21428 208366 21440
rect 390554 21428 390560 21440
rect 390612 21428 390618 21480
rect 84194 21360 84200 21412
rect 84252 21400 84258 21412
rect 104342 21400 104348 21412
rect 84252 21372 104348 21400
rect 84252 21360 84258 21372
rect 104342 21360 104348 21372
rect 104400 21360 104406 21412
rect 168098 21360 168104 21412
rect 168156 21400 168162 21412
rect 220814 21400 220820 21412
rect 168156 21372 220820 21400
rect 168156 21360 168162 21372
rect 220814 21360 220820 21372
rect 220872 21360 220878 21412
rect 232958 21360 232964 21412
rect 233016 21400 233022 21412
rect 498286 21400 498292 21412
rect 233016 21372 498292 21400
rect 233016 21360 233022 21372
rect 498286 21360 498292 21372
rect 498344 21360 498350 21412
rect 293954 20136 293960 20188
rect 294012 20176 294018 20188
rect 401778 20176 401784 20188
rect 294012 20148 401784 20176
rect 294012 20136 294018 20148
rect 401778 20136 401784 20148
rect 401836 20136 401842 20188
rect 143534 20068 143540 20120
rect 143592 20108 143598 20120
rect 255958 20108 255964 20120
rect 143592 20080 255964 20108
rect 143592 20068 143598 20080
rect 255958 20068 255964 20080
rect 256016 20068 256022 20120
rect 260834 20068 260840 20120
rect 260892 20108 260898 20120
rect 288434 20108 288440 20120
rect 260892 20080 288440 20108
rect 260892 20068 260898 20080
rect 288434 20068 288440 20080
rect 288492 20068 288498 20120
rect 333238 20068 333244 20120
rect 333296 20108 333302 20120
rect 452654 20108 452660 20120
rect 333296 20080 452660 20108
rect 333296 20068 333302 20080
rect 452654 20068 452660 20080
rect 452712 20068 452718 20120
rect 206646 20000 206652 20052
rect 206704 20040 206710 20052
rect 383654 20040 383660 20052
rect 206704 20012 383660 20040
rect 206704 20000 206710 20012
rect 383654 20000 383660 20012
rect 383712 20000 383718 20052
rect 461762 20000 461768 20052
rect 461820 20040 461826 20052
rect 542354 20040 542360 20052
rect 461820 20012 542360 20040
rect 461820 20000 461826 20012
rect 542354 20000 542360 20012
rect 542412 20000 542418 20052
rect 80054 19932 80060 19984
rect 80112 19972 80118 19984
rect 102778 19972 102784 19984
rect 80112 19944 102784 19972
rect 80112 19932 80118 19944
rect 102778 19932 102784 19944
rect 102836 19932 102842 19984
rect 168282 19932 168288 19984
rect 168340 19972 168346 19984
rect 218146 19972 218152 19984
rect 168340 19944 218152 19972
rect 168340 19932 168346 19944
rect 218146 19932 218152 19944
rect 218204 19932 218210 19984
rect 231762 19932 231768 19984
rect 231820 19972 231826 19984
rect 490006 19972 490012 19984
rect 231820 19944 490012 19972
rect 231820 19932 231826 19944
rect 490006 19932 490012 19944
rect 490064 19932 490070 19984
rect 357434 18844 357440 18896
rect 357492 18884 357498 18896
rect 417050 18884 417056 18896
rect 357492 18856 417056 18884
rect 357492 18844 357498 18856
rect 417050 18844 417056 18856
rect 417108 18844 417114 18896
rect 247034 18776 247040 18828
rect 247092 18816 247098 18828
rect 284386 18816 284392 18828
rect 247092 18788 284392 18816
rect 247092 18776 247098 18788
rect 284386 18776 284392 18788
rect 284444 18776 284450 18828
rect 322198 18776 322204 18828
rect 322256 18816 322262 18828
rect 403066 18816 403072 18828
rect 322256 18788 403072 18816
rect 322256 18776 322262 18788
rect 403066 18776 403072 18788
rect 403124 18776 403130 18828
rect 205266 18708 205272 18760
rect 205324 18748 205330 18760
rect 380894 18748 380900 18760
rect 205324 18720 380900 18748
rect 205324 18708 205330 18720
rect 380894 18708 380900 18720
rect 380952 18708 380958 18760
rect 66254 18640 66260 18692
rect 66312 18680 66318 18692
rect 100018 18680 100024 18692
rect 66312 18652 100024 18680
rect 66312 18640 66318 18652
rect 100018 18640 100024 18652
rect 100076 18640 100082 18692
rect 135254 18640 135260 18692
rect 135312 18680 135318 18692
rect 364334 18680 364340 18692
rect 135312 18652 364340 18680
rect 135312 18640 135318 18652
rect 364334 18640 364340 18652
rect 364392 18640 364398 18692
rect 460198 18640 460204 18692
rect 460256 18680 460262 18692
rect 539594 18680 539600 18692
rect 460256 18652 539600 18680
rect 460256 18640 460262 18652
rect 539594 18640 539600 18652
rect 539652 18640 539658 18692
rect 99374 18572 99380 18624
rect 99432 18612 99438 18624
rect 133322 18612 133328 18624
rect 99432 18584 133328 18612
rect 99432 18572 99438 18584
rect 133322 18572 133328 18584
rect 133380 18572 133386 18624
rect 164050 18572 164056 18624
rect 164108 18612 164114 18624
rect 202874 18612 202880 18624
rect 164108 18584 202880 18612
rect 164108 18572 164114 18584
rect 202874 18572 202880 18584
rect 202932 18572 202938 18624
rect 230198 18572 230204 18624
rect 230256 18612 230262 18624
rect 487154 18612 487160 18624
rect 230256 18584 487160 18612
rect 230256 18572 230262 18584
rect 487154 18572 487160 18584
rect 487212 18572 487218 18624
rect 200022 17416 200028 17468
rect 200080 17456 200086 17468
rect 356054 17456 356060 17468
rect 200080 17428 356060 17456
rect 200080 17416 200086 17428
rect 356054 17416 356060 17428
rect 356112 17416 356118 17468
rect 209774 17348 209780 17400
rect 209832 17388 209838 17400
rect 382366 17388 382372 17400
rect 209832 17360 382372 17388
rect 209832 17348 209838 17360
rect 382366 17348 382372 17360
rect 382424 17348 382430 17400
rect 60826 17280 60832 17332
rect 60884 17320 60890 17332
rect 71222 17320 71228 17332
rect 60884 17292 71228 17320
rect 60884 17280 60890 17292
rect 71222 17280 71228 17292
rect 71280 17280 71286 17332
rect 242986 17280 242992 17332
rect 243044 17320 243050 17332
rect 284570 17320 284576 17332
rect 243044 17292 284576 17320
rect 243044 17280 243050 17292
rect 284570 17280 284576 17292
rect 284628 17280 284634 17332
rect 305730 17280 305736 17332
rect 305788 17320 305794 17332
rect 332594 17320 332600 17332
rect 305788 17292 332600 17320
rect 305788 17280 305794 17292
rect 332594 17280 332600 17292
rect 332652 17280 332658 17332
rect 349798 17280 349804 17332
rect 349856 17320 349862 17332
rect 523126 17320 523132 17332
rect 349856 17292 523132 17320
rect 349856 17280 349862 17292
rect 523126 17280 523132 17292
rect 523184 17280 523190 17332
rect 16574 17212 16580 17264
rect 16632 17252 16638 17264
rect 61378 17252 61384 17264
rect 16632 17224 61384 17252
rect 16632 17212 16638 17224
rect 61378 17212 61384 17224
rect 61436 17212 61442 17264
rect 79870 17212 79876 17264
rect 79928 17252 79934 17264
rect 93854 17252 93860 17264
rect 79928 17224 93860 17252
rect 79928 17212 79934 17224
rect 93854 17212 93860 17224
rect 93912 17212 93918 17264
rect 102134 17212 102140 17264
rect 102192 17252 102198 17264
rect 108482 17252 108488 17264
rect 102192 17224 108488 17252
rect 102192 17212 102198 17224
rect 108482 17212 108488 17224
rect 108540 17212 108546 17264
rect 163866 17212 163872 17264
rect 163924 17252 163930 17264
rect 200114 17252 200120 17264
rect 163924 17224 200120 17252
rect 163924 17212 163930 17224
rect 200114 17212 200120 17224
rect 200172 17212 200178 17264
rect 228818 17212 228824 17264
rect 228876 17252 228882 17264
rect 480254 17252 480260 17264
rect 228876 17224 480260 17252
rect 228876 17212 228882 17224
rect 480254 17212 480260 17224
rect 480312 17212 480318 17264
rect 340966 16124 340972 16176
rect 341024 16164 341030 16176
rect 412910 16164 412916 16176
rect 341024 16136 412916 16164
rect 341024 16124 341030 16136
rect 412910 16124 412916 16136
rect 412968 16124 412974 16176
rect 272426 16056 272432 16108
rect 272484 16096 272490 16108
rect 291378 16096 291384 16108
rect 272484 16068 291384 16096
rect 272484 16056 272490 16068
rect 291378 16056 291384 16068
rect 291436 16056 291442 16108
rect 316218 16056 316224 16108
rect 316276 16096 316282 16108
rect 407206 16096 407212 16108
rect 316276 16068 407212 16096
rect 316276 16056 316282 16068
rect 407206 16056 407212 16068
rect 407264 16056 407270 16108
rect 162762 15988 162768 16040
rect 162820 16028 162826 16040
rect 196802 16028 196808 16040
rect 162820 16000 196808 16028
rect 162820 15988 162826 16000
rect 196802 15988 196808 16000
rect 196860 15988 196866 16040
rect 233418 15988 233424 16040
rect 233476 16028 233482 16040
rect 281534 16028 281540 16040
rect 233476 16000 281540 16028
rect 233476 15988 233482 16000
rect 281534 15988 281540 16000
rect 281592 15988 281598 16040
rect 305546 15988 305552 16040
rect 305604 16028 305610 16040
rect 404538 16028 404544 16040
rect 305604 16000 404544 16028
rect 305604 15988 305610 16000
rect 404538 15988 404544 16000
rect 404596 15988 404602 16040
rect 98178 15920 98184 15972
rect 98236 15960 98242 15972
rect 107102 15960 107108 15972
rect 98236 15932 107108 15960
rect 98236 15920 98242 15932
rect 107102 15920 107108 15932
rect 107160 15920 107166 15972
rect 184566 15920 184572 15972
rect 184624 15960 184630 15972
rect 288526 15960 288532 15972
rect 184624 15932 288532 15960
rect 184624 15920 184630 15932
rect 288526 15920 288532 15932
rect 288584 15920 288590 15972
rect 298094 15920 298100 15972
rect 298152 15960 298158 15972
rect 402974 15960 402980 15972
rect 298152 15932 402980 15960
rect 298152 15920 298158 15932
rect 402974 15920 402980 15932
rect 403032 15920 403038 15972
rect 446582 15920 446588 15972
rect 446640 15960 446646 15972
rect 482370 15960 482376 15972
rect 446640 15932 482376 15960
rect 446640 15920 446646 15932
rect 482370 15920 482376 15932
rect 482428 15920 482434 15972
rect 59354 15852 59360 15904
rect 59412 15892 59418 15904
rect 98822 15892 98828 15904
rect 59412 15864 98828 15892
rect 59412 15852 59418 15864
rect 98822 15852 98828 15864
rect 98880 15852 98886 15904
rect 180242 15852 180248 15904
rect 180300 15892 180306 15904
rect 269206 15892 269212 15904
rect 180300 15864 269212 15892
rect 180300 15852 180306 15864
rect 269206 15852 269212 15864
rect 269264 15852 269270 15904
rect 287146 15852 287152 15904
rect 287204 15892 287210 15904
rect 400306 15892 400312 15904
rect 287204 15864 400312 15892
rect 287204 15852 287210 15864
rect 400306 15852 400312 15864
rect 400364 15852 400370 15904
rect 459002 15852 459008 15904
rect 459060 15892 459066 15904
rect 536098 15892 536104 15904
rect 459060 15864 536104 15892
rect 459060 15852 459066 15864
rect 536098 15852 536104 15864
rect 536156 15852 536162 15904
rect 289814 15172 289820 15224
rect 289872 15212 289878 15224
rect 295518 15212 295524 15224
rect 289872 15184 295524 15212
rect 289872 15172 289878 15184
rect 295518 15172 295524 15184
rect 295576 15172 295582 15224
rect 255866 14968 255872 15020
rect 255924 15008 255930 15020
rect 393590 15008 393596 15020
rect 255924 14980 393596 15008
rect 255924 14968 255930 14980
rect 393590 14968 393596 14980
rect 393648 14968 393654 15020
rect 248414 14900 248420 14952
rect 248472 14940 248478 14952
rect 392118 14940 392124 14952
rect 248472 14912 392124 14940
rect 248472 14900 248478 14912
rect 392118 14900 392124 14912
rect 392176 14900 392182 14952
rect 241698 14832 241704 14884
rect 241756 14872 241762 14884
rect 389542 14872 389548 14884
rect 241756 14844 389548 14872
rect 241756 14832 241762 14844
rect 389542 14832 389548 14844
rect 389600 14832 389606 14884
rect 237650 14764 237656 14816
rect 237708 14804 237714 14816
rect 389358 14804 389364 14816
rect 237708 14776 389364 14804
rect 237708 14764 237714 14776
rect 389358 14764 389364 14776
rect 389416 14764 389422 14816
rect 234706 14696 234712 14748
rect 234764 14736 234770 14748
rect 387978 14736 387984 14748
rect 234764 14708 387984 14736
rect 234764 14696 234770 14708
rect 387978 14696 387984 14708
rect 388036 14696 388042 14748
rect 231026 14628 231032 14680
rect 231084 14668 231090 14680
rect 388162 14668 388168 14680
rect 231084 14640 388168 14668
rect 231084 14628 231090 14640
rect 388162 14628 388168 14640
rect 388220 14628 388226 14680
rect 227530 14560 227536 14612
rect 227588 14600 227594 14612
rect 386414 14600 386420 14612
rect 227588 14572 386420 14600
rect 227588 14560 227594 14572
rect 386414 14560 386420 14572
rect 386472 14560 386478 14612
rect 223574 14492 223580 14544
rect 223632 14532 223638 14544
rect 385402 14532 385408 14544
rect 223632 14504 385408 14532
rect 223632 14492 223638 14504
rect 385402 14492 385408 14504
rect 385460 14492 385466 14544
rect 84010 14424 84016 14476
rect 84068 14464 84074 14476
rect 114738 14464 114744 14476
rect 84068 14436 114744 14464
rect 84068 14424 84074 14436
rect 114738 14424 114744 14436
rect 114796 14424 114802 14476
rect 161290 14424 161296 14476
rect 161348 14464 161354 14476
rect 193306 14464 193312 14476
rect 161348 14436 193312 14464
rect 161348 14424 161354 14436
rect 193306 14424 193312 14436
rect 193364 14424 193370 14476
rect 219986 14424 219992 14476
rect 220044 14464 220050 14476
rect 385218 14464 385224 14476
rect 220044 14436 385224 14464
rect 220044 14424 220050 14436
rect 385218 14424 385224 14436
rect 385276 14424 385282 14476
rect 450722 14424 450728 14476
rect 450780 14464 450786 14476
rect 497090 14464 497096 14476
rect 450780 14436 497096 14464
rect 450780 14424 450786 14436
rect 497090 14424 497096 14436
rect 497148 14424 497154 14476
rect 155402 13336 155408 13388
rect 155460 13376 155466 13388
rect 258718 13376 258724 13388
rect 155460 13348 258724 13376
rect 155460 13336 155466 13348
rect 258718 13336 258724 13348
rect 258776 13336 258782 13388
rect 340322 13336 340328 13388
rect 340380 13376 340386 13388
rect 478138 13376 478144 13388
rect 340380 13348 478144 13376
rect 340380 13336 340386 13348
rect 478138 13336 478144 13348
rect 478196 13336 478202 13388
rect 188522 13268 188528 13320
rect 188580 13308 188586 13320
rect 376938 13308 376944 13320
rect 188580 13280 376944 13308
rect 188580 13268 188586 13280
rect 376938 13268 376944 13280
rect 376996 13268 377002 13320
rect 180978 13200 180984 13252
rect 181036 13240 181042 13252
rect 375650 13240 375656 13252
rect 181036 13212 375656 13240
rect 181036 13200 181042 13212
rect 375650 13200 375656 13212
rect 375708 13200 375714 13252
rect 177850 13132 177856 13184
rect 177908 13172 177914 13184
rect 375466 13172 375472 13184
rect 177908 13144 375472 13172
rect 177908 13132 177914 13144
rect 375466 13132 375472 13144
rect 375524 13132 375530 13184
rect 26234 13064 26240 13116
rect 26292 13104 26298 13116
rect 62758 13104 62764 13116
rect 26292 13076 62764 13104
rect 26292 13064 26298 13076
rect 62758 13064 62764 13076
rect 62816 13064 62822 13116
rect 82722 13064 82728 13116
rect 82780 13104 82786 13116
rect 108114 13104 108120 13116
rect 82780 13076 108120 13104
rect 82780 13064 82786 13076
rect 108114 13064 108120 13076
rect 108172 13064 108178 13116
rect 173894 13064 173900 13116
rect 173952 13104 173958 13116
rect 374178 13104 374184 13116
rect 173952 13076 374184 13104
rect 173952 13064 173958 13076
rect 374178 13064 374184 13076
rect 374236 13064 374242 13116
rect 376018 13064 376024 13116
rect 376076 13104 376082 13116
rect 418246 13104 418252 13116
rect 376076 13076 418252 13104
rect 376076 13064 376082 13076
rect 418246 13064 418252 13076
rect 418304 13064 418310 13116
rect 454862 13064 454868 13116
rect 454920 13104 454926 13116
rect 514846 13104 514852 13116
rect 454920 13076 514852 13104
rect 454920 13064 454926 13076
rect 514846 13064 514852 13076
rect 514904 13064 514910 13116
rect 300302 12384 300308 12436
rect 300360 12424 300366 12436
rect 307938 12424 307944 12436
rect 300360 12396 307944 12424
rect 300360 12384 300366 12396
rect 307938 12384 307944 12396
rect 307996 12384 308002 12436
rect 323578 12248 323584 12300
rect 323636 12288 323642 12300
rect 410794 12288 410800 12300
rect 323636 12260 410800 12288
rect 323636 12248 323642 12260
rect 410794 12248 410800 12260
rect 410852 12248 410858 12300
rect 153010 12180 153016 12232
rect 153068 12220 153074 12232
rect 157794 12220 157800 12232
rect 153068 12192 157800 12220
rect 153068 12180 153074 12192
rect 157794 12180 157800 12192
rect 157852 12180 157858 12232
rect 325142 12180 325148 12232
rect 325200 12220 325206 12232
rect 414290 12220 414296 12232
rect 325200 12192 414296 12220
rect 325200 12180 325206 12192
rect 414290 12180 414296 12192
rect 414348 12180 414354 12232
rect 324958 12112 324964 12164
rect 325016 12152 325022 12164
rect 417418 12152 417424 12164
rect 325016 12124 417424 12152
rect 325016 12112 325022 12124
rect 417418 12112 417424 12124
rect 417476 12112 417482 12164
rect 226334 12044 226340 12096
rect 226392 12084 226398 12096
rect 280338 12084 280344 12096
rect 226392 12056 280344 12084
rect 226392 12044 226398 12056
rect 280338 12044 280344 12056
rect 280396 12044 280402 12096
rect 327718 12044 327724 12096
rect 327776 12084 327782 12096
rect 423766 12084 423772 12096
rect 327776 12056 423772 12084
rect 327776 12044 327782 12056
rect 423766 12044 423772 12056
rect 423824 12044 423830 12096
rect 215294 11976 215300 12028
rect 215352 12016 215358 12028
rect 277394 12016 277400 12028
rect 215352 11988 277400 12016
rect 215352 11976 215358 11988
rect 277394 11976 277400 11988
rect 277452 11976 277458 12028
rect 327902 11976 327908 12028
rect 327960 12016 327966 12028
rect 427906 12016 427912 12028
rect 327960 11988 427912 12016
rect 327960 11976 327966 11988
rect 427906 11976 427912 11988
rect 427964 11976 427970 12028
rect 211706 11908 211712 11960
rect 211764 11948 211770 11960
rect 276290 11948 276296 11960
rect 211764 11920 276296 11948
rect 211764 11908 211770 11920
rect 276290 11908 276296 11920
rect 276348 11908 276354 11960
rect 329098 11908 329104 11960
rect 329156 11948 329162 11960
rect 432046 11948 432052 11960
rect 329156 11920 432052 11948
rect 329156 11908 329162 11920
rect 432046 11908 432052 11920
rect 432104 11908 432110 11960
rect 208578 11840 208584 11892
rect 208636 11880 208642 11892
rect 276106 11880 276112 11892
rect 208636 11852 276112 11880
rect 208636 11840 208642 11852
rect 276106 11840 276112 11852
rect 276164 11840 276170 11892
rect 329282 11840 329288 11892
rect 329340 11880 329346 11892
rect 434714 11880 434720 11892
rect 329340 11852 434720 11880
rect 329340 11840 329346 11852
rect 434714 11840 434720 11852
rect 434772 11840 434778 11892
rect 81250 11772 81256 11824
rect 81308 11812 81314 11824
rect 100754 11812 100760 11824
rect 81308 11784 100760 11812
rect 81308 11772 81314 11784
rect 100754 11772 100760 11784
rect 100812 11772 100818 11824
rect 129182 11812 129188 11824
rect 122806 11784 129188 11812
rect 11882 11704 11888 11756
rect 11940 11744 11946 11756
rect 57238 11744 57244 11756
rect 11940 11716 57244 11744
rect 11940 11704 11946 11716
rect 57238 11704 57244 11716
rect 57296 11704 57302 11756
rect 78122 11704 78128 11756
rect 78180 11744 78186 11756
rect 122806 11744 122834 11784
rect 129182 11772 129188 11784
rect 129240 11772 129246 11824
rect 205082 11772 205088 11824
rect 205140 11812 205146 11824
rect 274910 11812 274916 11824
rect 205140 11784 274916 11812
rect 205140 11772 205146 11784
rect 274910 11772 274916 11784
rect 274968 11772 274974 11824
rect 283098 11772 283104 11824
rect 283156 11812 283162 11824
rect 294138 11812 294144 11824
rect 283156 11784 294144 11812
rect 283156 11772 283162 11784
rect 294138 11772 294144 11784
rect 294196 11772 294202 11824
rect 330478 11772 330484 11824
rect 330536 11812 330542 11824
rect 439130 11812 439136 11824
rect 330536 11784 439136 11812
rect 330536 11772 330542 11784
rect 439130 11772 439136 11784
rect 439188 11772 439194 11824
rect 78180 11716 122834 11744
rect 78180 11704 78186 11716
rect 126974 11704 126980 11756
rect 127032 11744 127038 11756
rect 128170 11744 128176 11756
rect 127032 11716 128176 11744
rect 127032 11704 127038 11716
rect 128170 11704 128176 11716
rect 128228 11704 128234 11756
rect 158346 11704 158352 11756
rect 158404 11744 158410 11756
rect 178586 11744 178592 11756
rect 158404 11716 178592 11744
rect 158404 11704 158410 11716
rect 178586 11704 178592 11716
rect 178644 11704 178650 11756
rect 197906 11704 197912 11756
rect 197964 11744 197970 11756
rect 273346 11744 273352 11756
rect 197964 11716 273352 11744
rect 197964 11704 197970 11716
rect 273346 11704 273352 11716
rect 273404 11704 273410 11756
rect 279050 11704 279056 11756
rect 279108 11744 279114 11756
rect 292666 11744 292672 11756
rect 279108 11716 292672 11744
rect 279108 11704 279114 11716
rect 292666 11704 292672 11716
rect 292724 11704 292730 11756
rect 331858 11704 331864 11756
rect 331916 11744 331922 11756
rect 442166 11744 442172 11756
rect 331916 11716 442172 11744
rect 331916 11704 331922 11716
rect 442166 11704 442172 11716
rect 442224 11704 442230 11756
rect 447778 11704 447784 11756
rect 447836 11744 447842 11756
rect 486418 11744 486424 11756
rect 447836 11716 486424 11744
rect 447836 11704 447842 11716
rect 486418 11704 486424 11716
rect 486476 11704 486482 11756
rect 218054 11636 218060 11688
rect 218112 11676 218118 11688
rect 219250 11676 219256 11688
rect 218112 11648 219256 11676
rect 218112 11636 218118 11648
rect 219250 11636 219256 11648
rect 219308 11636 219314 11688
rect 234614 11636 234620 11688
rect 234672 11676 234678 11688
rect 235810 11676 235816 11688
rect 234672 11648 235816 11676
rect 234672 11636 234678 11648
rect 235810 11636 235816 11648
rect 235868 11636 235874 11688
rect 251266 10480 251272 10532
rect 251324 10520 251330 10532
rect 285674 10520 285680 10532
rect 251324 10492 285680 10520
rect 251324 10480 251330 10492
rect 285674 10480 285680 10492
rect 285732 10480 285738 10532
rect 313918 10480 313924 10532
rect 313976 10520 313982 10532
rect 367186 10520 367192 10532
rect 313976 10492 367192 10520
rect 313976 10480 313982 10492
rect 367186 10480 367192 10492
rect 367244 10480 367250 10532
rect 162026 10412 162032 10464
rect 162084 10452 162090 10464
rect 260098 10452 260104 10464
rect 162084 10424 260104 10452
rect 162084 10412 162090 10424
rect 260098 10412 260104 10424
rect 260156 10412 260162 10464
rect 284294 10412 284300 10464
rect 284352 10452 284358 10464
rect 400490 10452 400496 10464
rect 284352 10424 400496 10452
rect 284352 10412 284358 10424
rect 400490 10412 400496 10424
rect 400548 10412 400554 10464
rect 459186 10452 459192 10464
rect 447106 10424 459192 10452
rect 58434 10344 58440 10396
rect 58492 10384 58498 10396
rect 71038 10384 71044 10396
rect 58492 10356 71044 10384
rect 58492 10344 58498 10356
rect 71038 10344 71044 10356
rect 71096 10344 71102 10396
rect 77110 10344 77116 10396
rect 77168 10384 77174 10396
rect 86126 10384 86132 10396
rect 77168 10356 86132 10384
rect 77168 10344 77174 10356
rect 86126 10344 86132 10356
rect 86184 10344 86190 10396
rect 224586 10344 224592 10396
rect 224644 10384 224650 10396
rect 447106 10384 447134 10424
rect 459186 10412 459192 10424
rect 459244 10412 459250 10464
rect 224644 10356 447134 10384
rect 224644 10344 224650 10356
rect 458818 10344 458824 10396
rect 458876 10384 458882 10396
rect 532050 10384 532056 10396
rect 458876 10356 532056 10384
rect 458876 10344 458882 10356
rect 532050 10344 532056 10356
rect 532108 10344 532114 10396
rect 4798 10276 4804 10328
rect 4856 10316 4862 10328
rect 58618 10316 58624 10328
rect 4856 10288 58624 10316
rect 4856 10276 4862 10288
rect 58618 10276 58624 10288
rect 58676 10276 58682 10328
rect 84102 10276 84108 10328
rect 84160 10316 84166 10328
rect 110414 10316 110420 10328
rect 84160 10288 110420 10316
rect 84160 10276 84166 10288
rect 110414 10276 110420 10288
rect 110472 10276 110478 10328
rect 229002 10276 229008 10328
rect 229060 10316 229066 10328
rect 476482 10316 476488 10328
rect 229060 10288 476488 10316
rect 229060 10276 229066 10288
rect 476482 10276 476488 10288
rect 476540 10276 476546 10328
rect 76926 9596 76932 9648
rect 76984 9636 76990 9648
rect 83274 9636 83280 9648
rect 76984 9608 83280 9636
rect 76984 9596 76990 9608
rect 83274 9596 83280 9608
rect 83332 9596 83338 9648
rect 72602 9256 72608 9308
rect 72660 9296 72666 9308
rect 73798 9296 73804 9308
rect 72660 9268 73804 9296
rect 72660 9256 72666 9268
rect 73798 9256 73804 9268
rect 73856 9256 73862 9308
rect 209590 9188 209596 9240
rect 209648 9228 209654 9240
rect 395338 9228 395344 9240
rect 209648 9200 395344 9228
rect 209648 9188 209654 9200
rect 395338 9188 395344 9200
rect 395396 9188 395402 9240
rect 209406 9120 209412 9172
rect 209464 9160 209470 9172
rect 398926 9160 398932 9172
rect 209464 9132 398932 9160
rect 209464 9120 209470 9132
rect 398926 9120 398932 9132
rect 398984 9120 398990 9172
rect 453298 9120 453304 9172
rect 453356 9160 453362 9172
rect 507670 9160 507676 9172
rect 453356 9132 507676 9160
rect 453356 9120 453362 9132
rect 507670 9120 507676 9132
rect 507728 9120 507734 9172
rect 210786 9052 210792 9104
rect 210844 9092 210850 9104
rect 406010 9092 406016 9104
rect 210844 9064 406016 9092
rect 210844 9052 210850 9064
rect 406010 9052 406016 9064
rect 406068 9052 406074 9104
rect 453482 9052 453488 9104
rect 453540 9092 453546 9104
rect 511258 9092 511264 9104
rect 453540 9064 511264 9092
rect 453540 9052 453546 9064
rect 511258 9052 511264 9064
rect 511316 9052 511322 9104
rect 81066 8984 81072 9036
rect 81124 9024 81130 9036
rect 104526 9024 104532 9036
rect 81124 8996 104532 9024
rect 81124 8984 81130 8996
rect 104526 8984 104532 8996
rect 104584 8984 104590 9036
rect 157058 8984 157064 9036
rect 157116 9024 157122 9036
rect 175458 9024 175464 9036
rect 157116 8996 175464 9024
rect 157116 8984 157122 8996
rect 175458 8984 175464 8996
rect 175516 8984 175522 9036
rect 213546 8984 213552 9036
rect 213604 9024 213610 9036
rect 413094 9024 413100 9036
rect 213604 8996 413100 9024
rect 213604 8984 213610 8996
rect 413094 8984 413100 8996
rect 413152 8984 413158 9036
rect 454678 8984 454684 9036
rect 454736 9024 454742 9036
rect 518342 9024 518348 9036
rect 454736 8996 518348 9024
rect 454736 8984 454742 8996
rect 518342 8984 518348 8996
rect 518400 8984 518406 9036
rect 51350 8916 51356 8968
rect 51408 8956 51414 8968
rect 68278 8956 68284 8968
rect 51408 8928 68284 8956
rect 51408 8916 51414 8928
rect 68278 8916 68284 8928
rect 68336 8916 68342 8968
rect 96246 8916 96252 8968
rect 96304 8956 96310 8968
rect 133138 8956 133144 8968
rect 96304 8928 133144 8956
rect 96304 8916 96310 8928
rect 133138 8916 133144 8928
rect 133196 8916 133202 8968
rect 161106 8916 161112 8968
rect 161164 8956 161170 8968
rect 189718 8956 189724 8968
rect 161164 8928 189724 8956
rect 161164 8916 161170 8928
rect 189718 8916 189724 8928
rect 189776 8916 189782 8968
rect 213730 8916 213736 8968
rect 213788 8956 213794 8968
rect 416682 8956 416688 8968
rect 213788 8928 416688 8956
rect 213788 8916 213794 8928
rect 416682 8916 416688 8928
rect 416740 8916 416746 8968
rect 457438 8916 457444 8968
rect 457496 8956 457502 8968
rect 525426 8956 525432 8968
rect 457496 8928 525432 8956
rect 457496 8916 457502 8928
rect 525426 8916 525432 8928
rect 525484 8916 525490 8968
rect 75730 8236 75736 8288
rect 75788 8276 75794 8288
rect 79318 8276 79324 8288
rect 75788 8248 79324 8276
rect 75788 8236 75794 8248
rect 79318 8236 79324 8248
rect 79376 8236 79382 8288
rect 356698 8236 356704 8288
rect 356756 8276 356762 8288
rect 361482 8276 361488 8288
rect 356756 8248 361488 8276
rect 356756 8236 356762 8248
rect 361482 8236 361488 8248
rect 361540 8236 361546 8288
rect 312722 8168 312728 8220
rect 312780 8208 312786 8220
rect 364610 8208 364616 8220
rect 312780 8180 364616 8208
rect 312780 8168 312786 8180
rect 364610 8168 364616 8180
rect 364668 8168 364674 8220
rect 450538 8168 450544 8220
rect 450596 8208 450602 8220
rect 500586 8208 500592 8220
rect 450596 8180 500592 8208
rect 450596 8168 450602 8180
rect 500586 8168 500592 8180
rect 500644 8168 500650 8220
rect 356882 8100 356888 8152
rect 356940 8140 356946 8152
rect 549070 8140 549076 8152
rect 356940 8112 549076 8140
rect 356940 8100 356946 8112
rect 549070 8100 549076 8112
rect 549128 8100 549134 8152
rect 358078 8032 358084 8084
rect 358136 8072 358142 8084
rect 358136 8044 361436 8072
rect 358136 8032 358142 8044
rect 359458 7964 359464 8016
rect 359516 8004 359522 8016
rect 361408 8004 361436 8044
rect 361482 8032 361488 8084
rect 361540 8072 361546 8084
rect 552658 8072 552664 8084
rect 361540 8044 552664 8072
rect 361540 8032 361546 8044
rect 552658 8032 552664 8044
rect 552716 8032 552722 8084
rect 556154 8004 556160 8016
rect 359516 7976 361344 8004
rect 361408 7976 556160 8004
rect 359516 7964 359522 7976
rect 311158 7896 311164 7948
rect 311216 7936 311222 7948
rect 354030 7936 354036 7948
rect 311216 7908 354036 7936
rect 311216 7896 311222 7908
rect 354030 7896 354036 7908
rect 354088 7896 354094 7948
rect 359642 7896 359648 7948
rect 359700 7936 359706 7948
rect 361206 7936 361212 7948
rect 359700 7908 361212 7936
rect 359700 7896 359706 7908
rect 361206 7896 361212 7908
rect 361264 7896 361270 7948
rect 311342 7828 311348 7880
rect 311400 7868 311406 7880
rect 357526 7868 357532 7880
rect 311400 7840 357532 7868
rect 311400 7828 311406 7840
rect 357526 7828 357532 7840
rect 357584 7828 357590 7880
rect 361022 7828 361028 7880
rect 361080 7868 361086 7880
rect 361316 7868 361344 7976
rect 556154 7964 556160 7976
rect 556212 7964 556218 8016
rect 361390 7896 361396 7948
rect 361448 7936 361454 7948
rect 559742 7936 559748 7948
rect 361448 7908 559748 7936
rect 361448 7896 361454 7908
rect 559742 7896 559748 7908
rect 559800 7896 559806 7948
rect 563238 7868 563244 7880
rect 361080 7840 361252 7868
rect 361316 7840 563244 7868
rect 361080 7828 361086 7840
rect 312538 7760 312544 7812
rect 312596 7800 312602 7812
rect 361114 7800 361120 7812
rect 312596 7772 361120 7800
rect 312596 7760 312602 7772
rect 361114 7760 361120 7772
rect 361172 7760 361178 7812
rect 361224 7800 361252 7840
rect 563238 7828 563244 7840
rect 563296 7828 563302 7880
rect 566826 7800 566832 7812
rect 361224 7772 566832 7800
rect 566826 7760 566832 7772
rect 566884 7760 566890 7812
rect 91554 7692 91560 7744
rect 91612 7732 91618 7744
rect 105538 7732 105544 7744
rect 91612 7704 105544 7732
rect 91612 7692 91618 7704
rect 105538 7692 105544 7704
rect 105596 7692 105602 7744
rect 171962 7732 171968 7744
rect 166966 7704 171968 7732
rect 79686 7624 79692 7676
rect 79744 7664 79750 7676
rect 97442 7664 97448 7676
rect 79744 7636 97448 7664
rect 79744 7624 79750 7636
rect 97442 7624 97448 7636
rect 97500 7624 97506 7676
rect 157242 7624 157248 7676
rect 157300 7664 157306 7676
rect 166966 7664 166994 7704
rect 171962 7692 171968 7704
rect 172020 7692 172026 7744
rect 196986 7692 196992 7744
rect 197044 7732 197050 7744
rect 345750 7732 345756 7744
rect 197044 7704 345756 7732
rect 197044 7692 197050 7704
rect 345750 7692 345756 7704
rect 345808 7692 345814 7744
rect 360838 7692 360844 7744
rect 360896 7732 360902 7744
rect 570322 7732 570328 7744
rect 360896 7704 570328 7732
rect 360896 7692 360902 7704
rect 570322 7692 570328 7704
rect 570380 7692 570386 7744
rect 157300 7636 166994 7664
rect 157300 7624 157306 7636
rect 168374 7624 168380 7676
rect 168432 7664 168438 7676
rect 169570 7664 169576 7676
rect 168432 7636 169576 7664
rect 168432 7624 168438 7636
rect 169570 7624 169576 7636
rect 169628 7624 169634 7676
rect 198366 7624 198372 7676
rect 198424 7664 198430 7676
rect 349246 7664 349252 7676
rect 198424 7636 349252 7664
rect 198424 7624 198430 7636
rect 349246 7624 349252 7636
rect 349304 7624 349310 7676
rect 362218 7624 362224 7676
rect 362276 7664 362282 7676
rect 573910 7664 573916 7676
rect 362276 7636 573916 7664
rect 362276 7624 362282 7636
rect 573910 7624 573916 7636
rect 573968 7624 573974 7676
rect 54938 7556 54944 7608
rect 54996 7596 55002 7608
rect 69658 7596 69664 7608
rect 54996 7568 69664 7596
rect 54996 7556 55002 7568
rect 69658 7556 69664 7568
rect 69716 7556 69722 7608
rect 73798 7556 73804 7608
rect 73856 7596 73862 7608
rect 101398 7596 101404 7608
rect 73856 7568 101404 7596
rect 73856 7556 73862 7568
rect 101398 7556 101404 7568
rect 101456 7556 101462 7608
rect 103330 7556 103336 7608
rect 103388 7596 103394 7608
rect 134518 7596 134524 7608
rect 103388 7568 134524 7596
rect 103388 7556 103394 7568
rect 134518 7556 134524 7568
rect 134576 7556 134582 7608
rect 160002 7556 160008 7608
rect 160060 7596 160066 7608
rect 186130 7596 186136 7608
rect 160060 7568 186136 7596
rect 160060 7556 160066 7568
rect 186130 7556 186136 7568
rect 186188 7556 186194 7608
rect 198550 7556 198556 7608
rect 198608 7596 198614 7608
rect 352834 7596 352840 7608
rect 198608 7568 352840 7596
rect 198608 7556 198614 7568
rect 352834 7556 352840 7568
rect 352892 7556 352898 7608
rect 363598 7556 363604 7608
rect 363656 7596 363662 7608
rect 577406 7596 577412 7608
rect 363656 7568 577412 7596
rect 363656 7556 363662 7568
rect 577406 7556 577412 7568
rect 577464 7556 577470 7608
rect 105722 7488 105728 7540
rect 105780 7528 105786 7540
rect 108298 7528 108304 7540
rect 105780 7500 108304 7528
rect 105780 7488 105786 7500
rect 108298 7488 108304 7500
rect 108356 7488 108362 7540
rect 448606 7488 448612 7540
rect 448664 7528 448670 7540
rect 449802 7528 449808 7540
rect 448664 7500 449808 7528
rect 448664 7488 448670 7500
rect 449802 7488 449808 7500
rect 449860 7488 449866 7540
rect 265342 6672 265348 6724
rect 265400 6712 265406 6724
rect 288618 6712 288624 6724
rect 265400 6684 288624 6712
rect 265400 6672 265406 6684
rect 288618 6672 288624 6684
rect 288676 6672 288682 6724
rect 176470 6604 176476 6656
rect 176528 6644 176534 6656
rect 253474 6644 253480 6656
rect 176528 6616 253480 6644
rect 176528 6604 176534 6616
rect 253474 6604 253480 6616
rect 253532 6604 253538 6656
rect 254670 6604 254676 6656
rect 254728 6644 254734 6656
rect 287238 6644 287244 6656
rect 254728 6616 287244 6644
rect 254728 6604 254734 6616
rect 287238 6604 287244 6616
rect 287296 6604 287302 6656
rect 300118 6604 300124 6656
rect 300176 6644 300182 6656
rect 311434 6644 311440 6656
rect 300176 6616 311440 6644
rect 300176 6604 300182 6616
rect 311434 6604 311440 6616
rect 311492 6604 311498 6656
rect 340138 6604 340144 6656
rect 340196 6644 340202 6656
rect 481726 6644 481732 6656
rect 340196 6616 481732 6644
rect 340196 6604 340202 6616
rect 481726 6604 481732 6616
rect 481784 6604 481790 6656
rect 82078 6536 82084 6588
rect 82136 6576 82142 6588
rect 128998 6576 129004 6588
rect 82136 6548 129004 6576
rect 82136 6536 82142 6548
rect 128998 6536 129004 6548
rect 129056 6536 129062 6588
rect 176286 6536 176292 6588
rect 176344 6576 176350 6588
rect 257062 6576 257068 6588
rect 176344 6548 257068 6576
rect 176344 6536 176350 6548
rect 257062 6536 257068 6548
rect 257120 6536 257126 6588
rect 258258 6536 258264 6588
rect 258316 6576 258322 6588
rect 287422 6576 287428 6588
rect 258316 6548 287428 6576
rect 258316 6536 258322 6548
rect 287422 6536 287428 6548
rect 287480 6536 287486 6588
rect 301498 6536 301504 6588
rect 301556 6576 301562 6588
rect 315022 6576 315028 6588
rect 301556 6548 315028 6576
rect 301556 6536 301562 6548
rect 315022 6536 315028 6548
rect 315080 6536 315086 6588
rect 341702 6536 341708 6588
rect 341760 6576 341766 6588
rect 485222 6576 485228 6588
rect 341760 6548 485228 6576
rect 341760 6536 341766 6548
rect 485222 6536 485228 6548
rect 485280 6536 485286 6588
rect 41874 6468 41880 6520
rect 41932 6508 41938 6520
rect 93118 6508 93124 6520
rect 41932 6480 93124 6508
rect 41932 6468 41938 6480
rect 93118 6468 93124 6480
rect 93176 6468 93182 6520
rect 179322 6468 179328 6520
rect 179380 6508 179386 6520
rect 267734 6508 267740 6520
rect 179380 6480 267740 6508
rect 179380 6468 179386 6480
rect 267734 6468 267740 6480
rect 267792 6468 267798 6520
rect 303062 6468 303068 6520
rect 303120 6508 303126 6520
rect 318518 6508 318524 6520
rect 303120 6480 318524 6508
rect 303120 6468 303126 6480
rect 318518 6468 318524 6480
rect 318576 6468 318582 6520
rect 341518 6468 341524 6520
rect 341576 6508 341582 6520
rect 488810 6508 488816 6520
rect 341576 6480 488816 6508
rect 341576 6468 341582 6480
rect 488810 6468 488816 6480
rect 488868 6468 488874 6520
rect 74994 6400 75000 6452
rect 75052 6440 75058 6452
rect 127618 6440 127624 6452
rect 75052 6412 127624 6440
rect 75052 6400 75058 6412
rect 127618 6400 127624 6412
rect 127676 6400 127682 6452
rect 180702 6400 180708 6452
rect 180760 6440 180766 6452
rect 271230 6440 271236 6452
rect 180760 6412 271236 6440
rect 180760 6400 180766 6412
rect 271230 6400 271236 6412
rect 271288 6400 271294 6452
rect 302878 6400 302884 6452
rect 302936 6440 302942 6452
rect 322106 6440 322112 6452
rect 302936 6412 322112 6440
rect 302936 6400 302942 6412
rect 322106 6400 322112 6412
rect 322164 6400 322170 6452
rect 342990 6400 342996 6452
rect 343048 6440 343054 6452
rect 492306 6440 492312 6452
rect 343048 6412 492312 6440
rect 343048 6400 343054 6412
rect 492306 6400 492312 6412
rect 492364 6400 492370 6452
rect 38378 6332 38384 6384
rect 38436 6372 38442 6384
rect 93302 6372 93308 6384
rect 38436 6344 93308 6372
rect 38436 6332 38442 6344
rect 93302 6332 93308 6344
rect 93360 6332 93366 6384
rect 180610 6332 180616 6384
rect 180668 6372 180674 6384
rect 274818 6372 274824 6384
rect 180668 6344 274824 6372
rect 180668 6332 180674 6344
rect 274818 6332 274824 6344
rect 274876 6332 274882 6384
rect 276014 6332 276020 6384
rect 276072 6372 276078 6384
rect 291562 6372 291568 6384
rect 276072 6344 291568 6372
rect 276072 6332 276078 6344
rect 291562 6332 291568 6344
rect 291620 6332 291626 6384
rect 304442 6332 304448 6384
rect 304500 6372 304506 6384
rect 325602 6372 325608 6384
rect 304500 6344 325608 6372
rect 304500 6332 304506 6344
rect 325602 6332 325608 6344
rect 325660 6332 325666 6384
rect 345658 6332 345664 6384
rect 345716 6372 345722 6384
rect 502978 6372 502984 6384
rect 345716 6344 502984 6372
rect 345716 6332 345722 6344
rect 502978 6332 502984 6344
rect 503036 6332 503042 6384
rect 67910 6264 67916 6316
rect 67968 6304 67974 6316
rect 126238 6304 126244 6316
rect 67968 6276 126244 6304
rect 67968 6264 67974 6276
rect 126238 6264 126244 6276
rect 126296 6264 126302 6316
rect 181806 6264 181812 6316
rect 181864 6304 181870 6316
rect 278314 6304 278320 6316
rect 181864 6276 278320 6304
rect 181864 6264 181870 6276
rect 278314 6264 278320 6276
rect 278372 6264 278378 6316
rect 304258 6264 304264 6316
rect 304316 6304 304322 6316
rect 329190 6304 329196 6316
rect 304316 6276 329196 6304
rect 304316 6264 304322 6276
rect 329190 6264 329196 6276
rect 329248 6264 329254 6316
rect 345842 6264 345848 6316
rect 345900 6304 345906 6316
rect 506474 6304 506480 6316
rect 345900 6276 506480 6304
rect 345900 6264 345906 6276
rect 506474 6264 506480 6276
rect 506532 6264 506538 6316
rect 19426 6196 19432 6248
rect 19484 6236 19490 6248
rect 115382 6236 115388 6248
rect 19484 6208 115388 6236
rect 19484 6196 19490 6208
rect 115382 6196 115388 6208
rect 115440 6196 115446 6248
rect 181990 6196 181996 6248
rect 182048 6236 182054 6248
rect 281902 6236 281908 6248
rect 182048 6208 281908 6236
rect 182048 6196 182054 6208
rect 281902 6196 281908 6208
rect 281960 6196 281966 6248
rect 307018 6196 307024 6248
rect 307076 6236 307082 6248
rect 336274 6236 336280 6248
rect 307076 6208 336280 6236
rect 307076 6196 307082 6208
rect 336274 6196 336280 6208
rect 336332 6196 336338 6248
rect 347038 6196 347044 6248
rect 347096 6236 347102 6248
rect 510062 6236 510068 6248
rect 347096 6208 510068 6236
rect 347096 6196 347102 6208
rect 510062 6196 510068 6208
rect 510120 6196 510126 6248
rect 14734 6128 14740 6180
rect 14792 6168 14798 6180
rect 115198 6168 115204 6180
rect 14792 6140 115204 6168
rect 14792 6128 14798 6140
rect 115198 6128 115204 6140
rect 115256 6128 115262 6180
rect 129366 6128 129372 6180
rect 129424 6168 129430 6180
rect 145558 6168 145564 6180
rect 129424 6140 145564 6168
rect 129424 6128 129430 6140
rect 145558 6128 145564 6140
rect 145616 6128 145622 6180
rect 155862 6128 155868 6180
rect 155920 6168 155926 6180
rect 168374 6168 168380 6180
rect 155920 6140 168380 6168
rect 155920 6128 155926 6140
rect 168374 6128 168380 6140
rect 168432 6128 168438 6180
rect 183462 6128 183468 6180
rect 183520 6168 183526 6180
rect 285398 6168 285404 6180
rect 183520 6140 285404 6168
rect 183520 6128 183526 6140
rect 285398 6128 285404 6140
rect 285456 6128 285462 6180
rect 286594 6128 286600 6180
rect 286652 6168 286658 6180
rect 294046 6168 294052 6180
rect 286652 6140 294052 6168
rect 286652 6128 286658 6140
rect 294046 6128 294052 6140
rect 294104 6128 294110 6180
rect 307202 6128 307208 6180
rect 307260 6168 307266 6180
rect 339862 6168 339868 6180
rect 307260 6140 339868 6168
rect 307260 6128 307266 6140
rect 339862 6128 339868 6140
rect 339920 6128 339926 6180
rect 348418 6128 348424 6180
rect 348476 6168 348482 6180
rect 513558 6168 513564 6180
rect 348476 6140 513564 6168
rect 348476 6128 348482 6140
rect 513558 6128 513564 6140
rect 513616 6128 513622 6180
rect 298738 5584 298744 5636
rect 298796 5624 298802 5636
rect 304350 5624 304356 5636
rect 298796 5596 304356 5624
rect 298796 5584 298802 5596
rect 304350 5584 304356 5596
rect 304408 5584 304414 5636
rect 293678 5516 293684 5568
rect 293736 5556 293742 5568
rect 295702 5556 295708 5568
rect 293736 5528 295708 5556
rect 293736 5516 293742 5528
rect 295702 5516 295708 5528
rect 295760 5516 295766 5568
rect 298922 5516 298928 5568
rect 298980 5556 298986 5568
rect 300762 5556 300768 5568
rect 298980 5528 300768 5556
rect 298980 5516 298986 5528
rect 300762 5516 300768 5528
rect 300820 5516 300826 5568
rect 165430 5244 165436 5296
rect 165488 5284 165494 5296
rect 165488 5256 173894 5284
rect 165488 5244 165494 5256
rect 173866 5148 173894 5256
rect 207382 5148 207388 5160
rect 173866 5120 207388 5148
rect 207382 5108 207388 5120
rect 207440 5108 207446 5160
rect 238386 5108 238392 5160
rect 238444 5148 238450 5160
rect 519538 5148 519544 5160
rect 238444 5120 519544 5148
rect 238444 5108 238450 5120
rect 519538 5108 519544 5120
rect 519596 5108 519602 5160
rect 63218 5040 63224 5092
rect 63276 5080 63282 5092
rect 98638 5080 98644 5092
rect 63276 5052 98644 5080
rect 63276 5040 63282 5052
rect 98638 5040 98644 5052
rect 98696 5040 98702 5092
rect 165246 5040 165252 5092
rect 165304 5080 165310 5092
rect 210970 5080 210976 5092
rect 165304 5052 210976 5080
rect 165304 5040 165310 5052
rect 210970 5040 210976 5052
rect 211028 5040 211034 5092
rect 240042 5040 240048 5092
rect 240100 5080 240106 5092
rect 526622 5080 526628 5092
rect 240100 5052 526628 5080
rect 240100 5040 240106 5052
rect 526622 5040 526628 5052
rect 526680 5040 526686 5092
rect 56042 4972 56048 5024
rect 56100 5012 56106 5024
rect 97258 5012 97264 5024
rect 56100 4984 97264 5012
rect 56100 4972 56106 4984
rect 97258 4972 97264 4984
rect 97316 4972 97322 5024
rect 111610 4972 111616 5024
rect 111668 5012 111674 5024
rect 116394 5012 116400 5024
rect 111668 4984 116400 5012
rect 111668 4972 111674 4984
rect 116394 4972 116400 4984
rect 116452 4972 116458 5024
rect 166902 4972 166908 5024
rect 166960 5012 166966 5024
rect 214466 5012 214472 5024
rect 166960 4984 214472 5012
rect 166960 4972 166966 4984
rect 214466 4972 214472 4984
rect 214524 4972 214530 5024
rect 241330 4972 241336 5024
rect 241388 5012 241394 5024
rect 530118 5012 530124 5024
rect 241388 4984 530124 5012
rect 241388 4972 241394 4984
rect 530118 4972 530124 4984
rect 530176 4972 530182 5024
rect 37182 4904 37188 4956
rect 37240 4944 37246 4956
rect 65518 4944 65524 4956
rect 37240 4916 65524 4944
rect 37240 4904 37246 4916
rect 65518 4904 65524 4916
rect 65576 4904 65582 4956
rect 85666 4904 85672 4956
rect 85724 4944 85730 4956
rect 130378 4944 130384 4956
rect 85724 4916 130384 4944
rect 85724 4904 85730 4916
rect 130378 4904 130384 4916
rect 130436 4904 130442 4956
rect 136450 4904 136456 4956
rect 136508 4944 136514 4956
rect 148502 4944 148508 4956
rect 136508 4916 148508 4944
rect 136508 4904 136514 4916
rect 148502 4904 148508 4916
rect 148560 4904 148566 4956
rect 169662 4904 169668 4956
rect 169720 4944 169726 4956
rect 225138 4944 225144 4956
rect 169720 4916 225144 4944
rect 169720 4904 169726 4916
rect 225138 4904 225144 4916
rect 225196 4904 225202 4956
rect 241146 4904 241152 4956
rect 241204 4944 241210 4956
rect 533706 4944 533712 4956
rect 241204 4916 533712 4944
rect 241204 4904 241210 4916
rect 533706 4904 533712 4916
rect 533764 4904 533770 4956
rect 8754 4836 8760 4888
rect 8812 4876 8818 4888
rect 87598 4876 87604 4888
rect 8812 4848 87604 4876
rect 8812 4836 8818 4848
rect 87598 4836 87604 4848
rect 87656 4836 87662 4888
rect 95142 4836 95148 4888
rect 95200 4876 95206 4888
rect 106918 4876 106924 4888
rect 95200 4848 106924 4876
rect 95200 4836 95206 4848
rect 106918 4836 106924 4848
rect 106976 4836 106982 4888
rect 112990 4836 112996 4888
rect 113048 4876 113054 4888
rect 119890 4876 119896 4888
rect 113048 4848 119896 4876
rect 113048 4836 113054 4848
rect 119890 4836 119896 4848
rect 119948 4836 119954 4888
rect 169386 4836 169392 4888
rect 169444 4876 169450 4888
rect 228726 4876 228732 4888
rect 169444 4848 228732 4876
rect 169444 4836 169450 4848
rect 228726 4836 228732 4848
rect 228784 4836 228790 4888
rect 242526 4836 242532 4888
rect 242584 4876 242590 4888
rect 537202 4876 537208 4888
rect 242584 4848 537208 4876
rect 242584 4836 242590 4848
rect 537202 4836 537208 4848
rect 537260 4836 537266 4888
rect 4062 4768 4068 4820
rect 4120 4808 4126 4820
rect 86218 4808 86224 4820
rect 4120 4780 86224 4808
rect 4120 4768 4126 4780
rect 86218 4768 86224 4780
rect 86276 4768 86282 4820
rect 87966 4768 87972 4820
rect 88024 4808 88030 4820
rect 104158 4808 104164 4820
rect 88024 4780 104164 4808
rect 88024 4768 88030 4780
rect 104158 4768 104164 4780
rect 104216 4768 104222 4820
rect 113082 4768 113088 4820
rect 113140 4808 113146 4820
rect 123478 4808 123484 4820
rect 113140 4780 123484 4808
rect 113140 4768 113146 4780
rect 123478 4768 123484 4780
rect 123536 4768 123542 4820
rect 132954 4768 132960 4820
rect 133012 4808 133018 4820
rect 146938 4808 146944 4820
rect 133012 4780 146944 4808
rect 133012 4768 133018 4780
rect 146938 4768 146944 4780
rect 146996 4768 147002 4820
rect 154298 4768 154304 4820
rect 154356 4808 154362 4820
rect 164878 4808 164884 4820
rect 154356 4780 164884 4808
rect 154356 4768 154362 4780
rect 164878 4768 164884 4780
rect 164936 4768 164942 4820
rect 171042 4768 171048 4820
rect 171100 4808 171106 4820
rect 232222 4808 232228 4820
rect 171100 4780 232228 4808
rect 171100 4768 171106 4780
rect 232222 4768 232228 4780
rect 232280 4768 232286 4820
rect 242710 4768 242716 4820
rect 242768 4808 242774 4820
rect 540790 4808 540796 4820
rect 242768 4780 540796 4808
rect 242768 4768 242774 4780
rect 540790 4768 540796 4780
rect 540848 4768 540854 4820
rect 65518 4224 65524 4276
rect 65576 4264 65582 4276
rect 72418 4264 72424 4276
rect 65576 4236 72424 4264
rect 65576 4224 65582 4236
rect 72418 4224 72424 4236
rect 72476 4224 72482 4276
rect 69106 4156 69112 4208
rect 69164 4196 69170 4208
rect 72510 4196 72516 4208
rect 69164 4168 72516 4196
rect 69164 4156 69170 4168
rect 72510 4156 72516 4168
rect 72568 4156 72574 4208
rect 111426 4156 111432 4208
rect 111484 4196 111490 4208
rect 112806 4196 112812 4208
rect 111484 4168 112812 4196
rect 111484 4156 111490 4168
rect 112806 4156 112812 4168
rect 112864 4156 112870 4208
rect 153102 4156 153108 4208
rect 153160 4196 153166 4208
rect 154206 4196 154212 4208
rect 153160 4168 154212 4196
rect 153160 4156 153166 4168
rect 154206 4156 154212 4168
rect 154264 4156 154270 4208
rect 43070 4088 43076 4140
rect 43128 4128 43134 4140
rect 120902 4128 120908 4140
rect 43128 4100 120908 4128
rect 43128 4088 43134 4100
rect 120902 4088 120908 4100
rect 120960 4088 120966 4140
rect 167178 4088 167184 4140
rect 167236 4128 167242 4140
rect 170398 4128 170404 4140
rect 167236 4100 170404 4128
rect 167236 4088 167242 4100
rect 170398 4088 170404 4100
rect 170456 4088 170462 4140
rect 277118 4088 277124 4140
rect 277176 4128 277182 4140
rect 278038 4128 278044 4140
rect 277176 4100 278044 4128
rect 277176 4088 277182 4100
rect 278038 4088 278044 4100
rect 278096 4088 278102 4140
rect 333882 4088 333888 4140
rect 333940 4128 333946 4140
rect 336090 4128 336096 4140
rect 333940 4100 336096 4128
rect 333940 4088 333946 4100
rect 336090 4088 336096 4100
rect 336148 4088 336154 4140
rect 404814 4088 404820 4140
rect 404872 4128 404878 4140
rect 428182 4128 428188 4140
rect 404872 4100 428188 4128
rect 404872 4088 404878 4100
rect 428182 4088 428188 4100
rect 428240 4088 428246 4140
rect 463142 4088 463148 4140
rect 463200 4128 463206 4140
rect 550266 4128 550272 4140
rect 463200 4100 550272 4128
rect 463200 4088 463206 4100
rect 550266 4088 550272 4100
rect 550324 4088 550330 4140
rect 39574 4020 39580 4072
rect 39632 4060 39638 4072
rect 119522 4060 119528 4072
rect 39632 4032 119528 4060
rect 39632 4020 39638 4032
rect 119522 4020 119528 4032
rect 119580 4020 119586 4072
rect 401318 4020 401324 4072
rect 401376 4060 401382 4072
rect 427998 4060 428004 4072
rect 401376 4032 428004 4060
rect 401376 4020 401382 4032
rect 427998 4020 428004 4032
rect 428056 4020 428062 4072
rect 462958 4020 462964 4072
rect 463016 4060 463022 4072
rect 553762 4060 553768 4072
rect 463016 4032 553768 4060
rect 463016 4020 463022 4032
rect 553762 4020 553768 4032
rect 553820 4020 553826 4072
rect 35986 3952 35992 4004
rect 36044 3992 36050 4004
rect 119338 3992 119344 4004
rect 36044 3964 119344 3992
rect 36044 3952 36050 3964
rect 119338 3952 119344 3964
rect 119396 3952 119402 4004
rect 362310 3952 362316 4004
rect 362368 3992 362374 4004
rect 376018 3992 376024 4004
rect 362368 3964 376024 3992
rect 362368 3952 362374 3964
rect 376018 3952 376024 3964
rect 376076 3952 376082 4004
rect 397730 3952 397736 4004
rect 397788 3992 397794 4004
rect 426526 3992 426532 4004
rect 397788 3964 426532 3992
rect 397788 3952 397794 3964
rect 426526 3952 426532 3964
rect 426584 3952 426590 4004
rect 429654 3952 429660 4004
rect 429712 3992 429718 4004
rect 433518 3992 433524 4004
rect 429712 3964 433524 3992
rect 429712 3952 429718 3964
rect 433518 3952 433524 3964
rect 433576 3952 433582 4004
rect 464338 3952 464344 4004
rect 464396 3992 464402 4004
rect 557350 3992 557356 4004
rect 464396 3964 557356 3992
rect 464396 3952 464402 3964
rect 557350 3952 557356 3964
rect 557408 3952 557414 4004
rect 32490 3884 32496 3936
rect 32548 3924 32554 3936
rect 117958 3924 117964 3936
rect 32548 3896 117964 3924
rect 32548 3884 32554 3896
rect 117958 3884 117964 3896
rect 118016 3884 118022 3936
rect 124674 3884 124680 3936
rect 124732 3924 124738 3936
rect 140038 3924 140044 3936
rect 124732 3896 140044 3924
rect 124732 3884 124738 3896
rect 140038 3884 140044 3896
rect 140096 3884 140102 3936
rect 394234 3884 394240 3936
rect 394292 3924 394298 3936
rect 425054 3924 425060 3936
rect 394292 3896 425060 3924
rect 394292 3884 394298 3896
rect 425054 3884 425060 3896
rect 425112 3884 425118 3936
rect 438118 3884 438124 3936
rect 438176 3924 438182 3936
rect 447410 3924 447416 3936
rect 438176 3896 447416 3924
rect 438176 3884 438182 3896
rect 447410 3884 447416 3896
rect 447468 3884 447474 3936
rect 465902 3884 465908 3936
rect 465960 3924 465966 3936
rect 560846 3924 560852 3936
rect 465960 3896 560852 3924
rect 465960 3884 465966 3896
rect 560846 3884 560852 3896
rect 560904 3884 560910 3936
rect 28902 3816 28908 3868
rect 28960 3856 28966 3868
rect 116762 3856 116768 3868
rect 28960 3828 116768 3856
rect 28960 3816 28966 3828
rect 116762 3816 116768 3828
rect 116820 3816 116826 3868
rect 121086 3816 121092 3868
rect 121144 3856 121150 3868
rect 138658 3856 138664 3868
rect 121144 3828 138664 3856
rect 121144 3816 121150 3828
rect 138658 3816 138664 3828
rect 138716 3816 138722 3868
rect 371418 3856 371424 3868
rect 365548 3828 371424 3856
rect 24210 3748 24216 3800
rect 24268 3788 24274 3800
rect 116578 3788 116584 3800
rect 24268 3760 116584 3788
rect 24268 3748 24274 3760
rect 116578 3748 116584 3760
rect 116636 3748 116642 3800
rect 117590 3748 117596 3800
rect 117648 3788 117654 3800
rect 137278 3788 137284 3800
rect 117648 3760 137284 3788
rect 117648 3748 117654 3760
rect 137278 3748 137284 3760
rect 137336 3748 137342 3800
rect 140038 3748 140044 3800
rect 140096 3788 140102 3800
rect 148318 3788 148324 3800
rect 140096 3760 148324 3788
rect 140096 3748 140102 3760
rect 148318 3748 148324 3760
rect 148376 3748 148382 3800
rect 193214 3748 193220 3800
rect 193272 3788 193278 3800
rect 194410 3788 194416 3800
rect 193272 3760 194416 3788
rect 193272 3748 193278 3760
rect 194410 3748 194416 3760
rect 194468 3748 194474 3800
rect 251174 3748 251180 3800
rect 251232 3788 251238 3800
rect 252370 3788 252376 3800
rect 251232 3760 252376 3788
rect 251232 3748 251238 3760
rect 252370 3748 252376 3760
rect 252428 3748 252434 3800
rect 365548 3788 365576 3828
rect 371418 3816 371424 3828
rect 371476 3816 371482 3868
rect 390646 3816 390652 3868
rect 390704 3856 390710 3868
rect 425146 3856 425152 3868
rect 390704 3828 425152 3856
rect 390704 3816 390710 3828
rect 425146 3816 425152 3828
rect 425204 3816 425210 3868
rect 439498 3816 439504 3868
rect 439556 3856 439562 3868
rect 450906 3856 450912 3868
rect 439556 3828 450912 3856
rect 439556 3816 439562 3828
rect 450906 3816 450912 3828
rect 450964 3816 450970 3868
rect 465718 3816 465724 3868
rect 465776 3856 465782 3868
rect 564434 3856 564440 3868
rect 465776 3828 564440 3856
rect 465776 3816 465782 3828
rect 564434 3816 564440 3828
rect 564492 3816 564498 3868
rect 354646 3760 365576 3788
rect 25314 3680 25320 3732
rect 25372 3720 25378 3732
rect 142798 3720 142804 3732
rect 25372 3692 142804 3720
rect 25372 3680 25378 3692
rect 142798 3680 142804 3692
rect 142856 3680 142862 3732
rect 160186 3680 160192 3732
rect 160244 3720 160250 3732
rect 354646 3720 354674 3760
rect 365806 3748 365812 3800
rect 365864 3788 365870 3800
rect 418430 3788 418436 3800
rect 365864 3760 418436 3788
rect 365864 3748 365870 3760
rect 418430 3748 418436 3760
rect 418488 3748 418494 3800
rect 440878 3748 440884 3800
rect 440936 3788 440942 3800
rect 454494 3788 454500 3800
rect 440936 3760 454500 3788
rect 440936 3748 440942 3760
rect 454494 3748 454500 3760
rect 454552 3748 454558 3800
rect 467282 3748 467288 3800
rect 467340 3788 467346 3800
rect 568022 3788 568028 3800
rect 467340 3760 568028 3788
rect 467340 3748 467346 3760
rect 568022 3748 568028 3760
rect 568080 3748 568086 3800
rect 369946 3720 369952 3732
rect 160244 3692 354674 3720
rect 365548 3692 369952 3720
rect 160244 3680 160250 3692
rect 20622 3612 20628 3664
rect 20680 3652 20686 3664
rect 141602 3652 141608 3664
rect 20680 3624 141608 3652
rect 20680 3612 20686 3624
rect 141602 3612 141608 3624
rect 141660 3612 141666 3664
rect 156598 3612 156604 3664
rect 156656 3652 156662 3664
rect 365548 3652 365576 3692
rect 369946 3680 369952 3692
rect 370004 3680 370010 3732
rect 387150 3680 387156 3732
rect 387208 3720 387214 3732
rect 424134 3720 424140 3732
rect 387208 3692 424140 3720
rect 387208 3680 387214 3692
rect 424134 3680 424140 3692
rect 424192 3680 424198 3732
rect 441062 3680 441068 3732
rect 441120 3720 441126 3732
rect 458082 3720 458088 3732
rect 441120 3692 458088 3720
rect 441120 3680 441126 3692
rect 458082 3680 458088 3692
rect 458140 3680 458146 3732
rect 467098 3680 467104 3732
rect 467156 3720 467162 3732
rect 571518 3720 571524 3732
rect 467156 3692 571524 3720
rect 467156 3680 467162 3692
rect 571518 3680 571524 3692
rect 571576 3680 571582 3732
rect 156656 3624 365576 3652
rect 156656 3612 156662 3624
rect 365622 3612 365628 3664
rect 365680 3652 365686 3664
rect 368566 3652 368572 3664
rect 365680 3624 368572 3652
rect 365680 3612 365686 3624
rect 368566 3612 368572 3624
rect 368624 3612 368630 3664
rect 383562 3612 383568 3664
rect 383620 3652 383626 3664
rect 423950 3652 423956 3664
rect 383620 3624 423956 3652
rect 383620 3612 383626 3624
rect 423950 3612 423956 3624
rect 424008 3612 424014 3664
rect 442258 3612 442264 3664
rect 442316 3652 442322 3664
rect 461578 3652 461584 3664
rect 442316 3624 461584 3652
rect 442316 3612 442322 3624
rect 461578 3612 461584 3624
rect 461636 3612 461642 3664
rect 468478 3612 468484 3664
rect 468536 3652 468542 3664
rect 575106 3652 575112 3664
rect 468536 3624 575112 3652
rect 468536 3612 468542 3624
rect 575106 3612 575112 3624
rect 575164 3612 575170 3664
rect 11146 3544 11152 3596
rect 11204 3584 11210 3596
rect 11204 3556 14596 3584
rect 11204 3544 11210 3556
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 4798 3516 4804 3528
rect 2924 3488 4804 3516
rect 2924 3476 2930 3488
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 13538 3476 13544 3528
rect 13596 3516 13602 3528
rect 14458 3516 14464 3528
rect 13596 3488 14464 3516
rect 13596 3476 13602 3488
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 14568 3516 14596 3556
rect 15930 3544 15936 3596
rect 15988 3584 15994 3596
rect 141418 3584 141424 3596
rect 15988 3556 141424 3584
rect 15988 3544 15994 3556
rect 141418 3544 141424 3556
rect 141476 3544 141482 3596
rect 160094 3544 160100 3596
rect 160152 3584 160158 3596
rect 161290 3584 161296 3596
rect 160152 3556 161296 3584
rect 160152 3544 160158 3556
rect 161290 3544 161296 3556
rect 161348 3544 161354 3596
rect 161382 3544 161388 3596
rect 161440 3584 161446 3596
rect 368474 3584 368480 3596
rect 161440 3556 368480 3584
rect 161440 3544 161446 3556
rect 368474 3544 368480 3556
rect 368532 3544 368538 3596
rect 379974 3544 379980 3596
rect 380032 3584 380038 3596
rect 422294 3584 422300 3596
rect 380032 3556 422300 3584
rect 380032 3544 380038 3556
rect 422294 3544 422300 3556
rect 422352 3544 422358 3596
rect 442442 3544 442448 3596
rect 442500 3584 442506 3596
rect 442500 3556 442580 3584
rect 442500 3544 442506 3556
rect 140222 3516 140228 3528
rect 14568 3488 140228 3516
rect 140222 3476 140228 3488
rect 140280 3476 140286 3528
rect 143534 3476 143540 3528
rect 143592 3516 143598 3528
rect 144730 3516 144736 3528
rect 143592 3488 144736 3516
rect 143592 3476 143598 3488
rect 144730 3476 144736 3488
rect 144788 3476 144794 3528
rect 149514 3476 149520 3528
rect 149572 3516 149578 3528
rect 365622 3516 365628 3528
rect 149572 3488 365628 3516
rect 149572 3476 149578 3488
rect 365622 3476 365628 3488
rect 365680 3476 365686 3528
rect 365714 3476 365720 3528
rect 365772 3516 365778 3528
rect 367002 3516 367008 3528
rect 365772 3488 367008 3516
rect 365772 3476 365778 3488
rect 367002 3476 367008 3488
rect 367060 3476 367066 3528
rect 373994 3476 374000 3528
rect 374052 3516 374058 3528
rect 375282 3516 375288 3528
rect 374052 3488 375288 3516
rect 374052 3476 374058 3488
rect 375282 3476 375288 3488
rect 375340 3476 375346 3528
rect 376478 3476 376484 3528
rect 376536 3516 376542 3528
rect 421098 3516 421104 3528
rect 376536 3488 421104 3516
rect 376536 3476 376542 3488
rect 421098 3476 421104 3488
rect 421156 3476 421162 3528
rect 423766 3476 423772 3528
rect 423824 3516 423830 3528
rect 424962 3516 424968 3528
rect 423824 3488 424968 3516
rect 423824 3476 423830 3488
rect 424962 3476 424968 3488
rect 425020 3476 425026 3528
rect 432138 3516 432144 3528
rect 425072 3488 432144 3516
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 144362 3448 144368 3460
rect 6512 3420 144368 3448
rect 6512 3408 6518 3420
rect 144362 3408 144368 3420
rect 144420 3408 144426 3460
rect 145926 3408 145932 3460
rect 145984 3448 145990 3460
rect 367278 3448 367284 3460
rect 145984 3420 367284 3448
rect 145984 3408 145990 3420
rect 367278 3408 367284 3420
rect 367336 3408 367342 3460
rect 372890 3408 372896 3460
rect 372948 3448 372954 3460
rect 421282 3448 421288 3460
rect 372948 3420 421288 3448
rect 372948 3408 372954 3420
rect 421282 3408 421288 3420
rect 421340 3408 421346 3460
rect 422570 3408 422576 3460
rect 422628 3448 422634 3460
rect 425072 3448 425100 3488
rect 432138 3476 432144 3488
rect 432196 3476 432202 3528
rect 440326 3476 440332 3528
rect 440384 3516 440390 3528
rect 441522 3516 441528 3528
rect 440384 3488 441528 3516
rect 440384 3476 440390 3488
rect 441522 3476 441528 3488
rect 441580 3476 441586 3528
rect 422628 3420 425100 3448
rect 422628 3408 422634 3420
rect 426158 3408 426164 3460
rect 426216 3448 426222 3460
rect 433702 3448 433708 3460
rect 426216 3420 433708 3448
rect 426216 3408 426222 3420
rect 433702 3408 433708 3420
rect 433760 3408 433766 3460
rect 31294 3340 31300 3392
rect 31352 3380 31358 3392
rect 32398 3380 32404 3392
rect 31352 3352 32404 3380
rect 31352 3340 31358 3352
rect 32398 3340 32404 3352
rect 32456 3340 32462 3392
rect 46658 3340 46664 3392
rect 46716 3380 46722 3392
rect 120718 3380 120724 3392
rect 46716 3352 120724 3380
rect 46716 3340 46722 3352
rect 120718 3340 120724 3352
rect 120776 3340 120782 3392
rect 153010 3340 153016 3392
rect 153068 3380 153074 3392
rect 161382 3380 161388 3392
rect 153068 3352 161388 3380
rect 153068 3340 153074 3352
rect 161382 3340 161388 3352
rect 161440 3340 161446 3392
rect 213362 3340 213368 3392
rect 213420 3380 213426 3392
rect 214558 3380 214564 3392
rect 213420 3352 214564 3380
rect 213420 3340 213426 3352
rect 214558 3340 214564 3352
rect 214616 3340 214622 3392
rect 301958 3340 301964 3392
rect 302016 3380 302022 3392
rect 305638 3380 305644 3392
rect 302016 3352 305644 3380
rect 302016 3340 302022 3352
rect 305638 3340 305644 3352
rect 305696 3340 305702 3392
rect 309042 3340 309048 3392
rect 309100 3380 309106 3392
rect 309870 3380 309876 3392
rect 309100 3352 309876 3380
rect 309100 3340 309106 3352
rect 309870 3340 309876 3352
rect 309928 3340 309934 3392
rect 316034 3340 316040 3392
rect 316092 3380 316098 3392
rect 317322 3380 317328 3392
rect 316092 3352 317328 3380
rect 316092 3340 316098 3352
rect 317322 3340 317328 3352
rect 317380 3340 317386 3392
rect 357434 3340 357440 3392
rect 357492 3380 357498 3392
rect 358722 3380 358728 3392
rect 357492 3352 358728 3380
rect 357492 3340 357498 3352
rect 358722 3340 358728 3352
rect 358780 3340 358786 3392
rect 390554 3340 390560 3392
rect 390612 3380 390618 3392
rect 391842 3380 391848 3392
rect 390612 3352 391848 3380
rect 390612 3340 390618 3352
rect 391842 3340 391848 3352
rect 391900 3340 391906 3392
rect 398834 3340 398840 3392
rect 398892 3380 398898 3392
rect 400122 3380 400128 3392
rect 398892 3352 400128 3380
rect 398892 3340 398898 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 408402 3340 408408 3392
rect 408460 3380 408466 3392
rect 429194 3380 429200 3392
rect 408460 3352 429200 3380
rect 408460 3340 408466 3352
rect 429194 3340 429200 3352
rect 429252 3340 429258 3392
rect 436830 3340 436836 3392
rect 436888 3380 436894 3392
rect 440326 3380 440332 3392
rect 436888 3352 440332 3380
rect 436888 3340 436894 3352
rect 440326 3340 440332 3352
rect 440384 3340 440390 3392
rect 442552 3380 442580 3556
rect 445202 3544 445208 3596
rect 445260 3584 445266 3596
rect 472250 3584 472256 3596
rect 445260 3556 472256 3584
rect 445260 3544 445266 3556
rect 472250 3544 472256 3556
rect 472308 3544 472314 3596
rect 472618 3544 472624 3596
rect 472676 3584 472682 3596
rect 582190 3584 582196 3596
rect 472676 3556 582196 3584
rect 472676 3544 472682 3556
rect 582190 3544 582196 3556
rect 582248 3544 582254 3596
rect 444346 3488 448560 3516
rect 443638 3408 443644 3460
rect 443696 3448 443702 3460
rect 444346 3448 444374 3488
rect 443696 3420 444374 3448
rect 448532 3448 448560 3488
rect 449158 3476 449164 3528
rect 449216 3516 449222 3528
rect 465166 3516 465172 3528
rect 449216 3488 465172 3516
rect 449216 3476 449222 3488
rect 465166 3476 465172 3488
rect 465224 3476 465230 3528
rect 470134 3476 470140 3528
rect 470192 3516 470198 3528
rect 578602 3516 578608 3528
rect 470192 3488 578608 3516
rect 470192 3476 470198 3488
rect 578602 3476 578608 3488
rect 578660 3476 578666 3528
rect 468662 3448 468668 3460
rect 448532 3420 468668 3448
rect 443696 3408 443702 3420
rect 468662 3408 468668 3420
rect 468720 3408 468726 3460
rect 471238 3408 471244 3460
rect 471296 3448 471302 3460
rect 580994 3448 581000 3460
rect 471296 3420 581000 3448
rect 471296 3408 471302 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 449158 3380 449164 3392
rect 442552 3352 449164 3380
rect 449158 3340 449164 3352
rect 449216 3340 449222 3392
rect 461670 3340 461676 3392
rect 461728 3380 461734 3392
rect 546678 3380 546684 3392
rect 461728 3352 546684 3380
rect 461728 3340 461734 3352
rect 546678 3340 546684 3352
rect 546736 3340 546742 3392
rect 110506 3272 110512 3324
rect 110564 3312 110570 3324
rect 135898 3312 135904 3324
rect 110564 3284 135904 3312
rect 110564 3272 110570 3284
rect 135898 3272 135904 3284
rect 135956 3272 135962 3324
rect 326798 3272 326804 3324
rect 326856 3312 326862 3324
rect 330570 3312 330576 3324
rect 326856 3284 330576 3312
rect 326856 3272 326862 3284
rect 330570 3272 330576 3284
rect 330628 3272 330634 3324
rect 351638 3272 351644 3324
rect 351696 3312 351702 3324
rect 353938 3312 353944 3324
rect 351696 3284 353944 3312
rect 351696 3272 351702 3284
rect 353938 3272 353944 3284
rect 353996 3272 354002 3324
rect 411898 3272 411904 3324
rect 411956 3312 411962 3324
rect 429286 3312 429292 3324
rect 411956 3284 429292 3312
rect 411956 3272 411962 3284
rect 429286 3272 429292 3284
rect 429344 3272 429350 3324
rect 433242 3272 433248 3324
rect 433300 3312 433306 3324
rect 434806 3312 434812 3324
rect 433300 3284 434812 3312
rect 433300 3272 433306 3284
rect 434806 3272 434812 3284
rect 434864 3272 434870 3324
rect 438302 3272 438308 3324
rect 438360 3312 438366 3324
rect 443822 3312 443828 3324
rect 438360 3284 443828 3312
rect 438360 3272 438366 3284
rect 443822 3272 443828 3284
rect 443880 3272 443886 3324
rect 446398 3272 446404 3324
rect 446456 3312 446462 3324
rect 479334 3312 479340 3324
rect 446456 3284 479340 3312
rect 446456 3272 446462 3284
rect 479334 3272 479340 3284
rect 479392 3272 479398 3324
rect 498194 3272 498200 3324
rect 498252 3312 498258 3324
rect 499022 3312 499028 3324
rect 498252 3284 499028 3312
rect 498252 3272 498258 3284
rect 499022 3272 499028 3284
rect 499080 3272 499086 3324
rect 514754 3272 514760 3324
rect 514812 3312 514818 3324
rect 515582 3312 515588 3324
rect 514812 3284 515588 3312
rect 514812 3272 514818 3284
rect 515582 3272 515588 3284
rect 515640 3272 515646 3324
rect 110414 3204 110420 3256
rect 110472 3244 110478 3256
rect 111610 3244 111616 3256
rect 110472 3216 111616 3244
rect 110472 3204 110478 3216
rect 111610 3204 111616 3216
rect 111668 3204 111674 3256
rect 114002 3204 114008 3256
rect 114060 3244 114066 3256
rect 137462 3244 137468 3256
rect 114060 3216 137468 3244
rect 114060 3204 114066 3216
rect 137462 3204 137468 3216
rect 137520 3204 137526 3256
rect 319714 3204 319720 3256
rect 319772 3244 319778 3256
rect 320818 3244 320824 3256
rect 319772 3216 320824 3244
rect 319772 3204 319778 3216
rect 320818 3204 320824 3216
rect 320876 3204 320882 3256
rect 415486 3204 415492 3256
rect 415544 3244 415550 3256
rect 430666 3244 430672 3256
rect 415544 3216 430672 3244
rect 415544 3204 415550 3216
rect 430666 3204 430672 3216
rect 430724 3204 430730 3256
rect 445110 3204 445116 3256
rect 445168 3244 445174 3256
rect 475746 3244 475752 3256
rect 445168 3216 475752 3244
rect 445168 3204 445174 3216
rect 475746 3204 475752 3216
rect 475804 3204 475810 3256
rect 566 3136 572 3188
rect 624 3176 630 3188
rect 3418 3176 3424 3188
rect 624 3148 3424 3176
rect 624 3136 630 3148
rect 3418 3136 3424 3148
rect 3476 3136 3482 3188
rect 337470 3136 337476 3188
rect 337528 3176 337534 3188
rect 338758 3176 338764 3188
rect 337528 3148 338764 3176
rect 337528 3136 337534 3148
rect 338758 3136 338764 3148
rect 338816 3136 338822 3188
rect 348050 3136 348056 3188
rect 348108 3176 348114 3188
rect 352558 3176 352564 3188
rect 348108 3148 352564 3176
rect 348108 3136 348114 3148
rect 352558 3136 352564 3148
rect 352616 3136 352622 3188
rect 418982 3136 418988 3188
rect 419040 3176 419046 3188
rect 432322 3176 432328 3188
rect 419040 3148 432328 3176
rect 419040 3136 419046 3148
rect 432322 3136 432328 3148
rect 432380 3136 432386 3188
rect 147122 3068 147128 3120
rect 147180 3108 147186 3120
rect 149698 3108 149704 3120
rect 147180 3080 149704 3108
rect 147180 3068 147186 3080
rect 149698 3068 149704 3080
rect 149756 3068 149762 3120
rect 355226 3000 355232 3052
rect 355284 3040 355290 3052
rect 358170 3040 358176 3052
rect 355284 3012 358176 3040
rect 355284 3000 355290 3012
rect 358170 3000 358176 3012
rect 358228 3000 358234 3052
rect 143534 2932 143540 2984
rect 143592 2972 143598 2984
rect 149882 2972 149888 2984
rect 143592 2944 149888 2972
rect 143592 2932 143598 2944
rect 149882 2932 149888 2944
rect 149940 2932 149946 2984
rect 184934 2932 184940 2984
rect 184992 2972 184998 2984
rect 186958 2972 186964 2984
rect 184992 2944 186964 2972
rect 184992 2932 184998 2944
rect 186958 2932 186964 2944
rect 187016 2932 187022 2984
rect 340874 1368 340880 1420
rect 340932 1408 340938 1420
rect 342162 1408 342168 1420
rect 340932 1380 342168 1408
rect 340932 1368 340938 1380
rect 342162 1368 342168 1380
rect 342220 1368 342226 1420
rect 349154 1368 349160 1420
rect 349212 1408 349218 1420
rect 350442 1408 350448 1420
rect 349212 1380 350448 1408
rect 349212 1368 349218 1380
rect 350442 1368 350448 1380
rect 350500 1368 350506 1420
<< via1 >>
rect 1400 448536 1452 448588
rect 57612 448536 57664 448588
rect 314292 59780 314344 59832
rect 315396 59780 315448 59832
rect 357532 59780 357584 59832
rect 359464 59780 359516 59832
rect 422392 59780 422444 59832
rect 424140 59780 424192 59832
rect 63408 59712 63460 59764
rect 64236 59712 64288 59764
rect 67548 59712 67600 59764
rect 68468 59712 68520 59764
rect 68928 59712 68980 59764
rect 70124 59712 70176 59764
rect 72700 59712 72752 59764
rect 74632 59712 74684 59764
rect 81072 59712 81124 59764
rect 83464 59712 83516 59764
rect 86224 59712 86276 59764
rect 88432 59712 88484 59764
rect 88984 59712 89036 59764
rect 91744 59712 91796 59764
rect 96068 59712 96120 59764
rect 98368 59712 98420 59764
rect 98644 59712 98696 59764
rect 100852 59712 100904 59764
rect 113088 59712 113140 59764
rect 115020 59712 115072 59764
rect 122748 59712 122800 59764
rect 123300 59712 123352 59764
rect 125140 59712 125192 59764
rect 127532 59712 127584 59764
rect 134524 59712 134576 59764
rect 136640 59712 136692 59764
rect 140228 59712 140280 59764
rect 142436 59712 142488 59764
rect 148508 59712 148560 59764
rect 149428 59712 149480 59764
rect 151728 59712 151780 59764
rect 152464 59712 152516 59764
rect 154304 59712 154356 59764
rect 156604 59712 156656 59764
rect 158536 59712 158588 59764
rect 160744 59712 160796 59764
rect 165252 59712 165304 59764
rect 167460 59712 167512 59764
rect 173624 59712 173676 59764
rect 175740 59712 175792 59764
rect 180616 59712 180668 59764
rect 182364 59712 182416 59764
rect 184572 59712 184624 59764
rect 185676 59712 185728 59764
rect 188712 59712 188764 59764
rect 189908 59712 189960 59764
rect 202696 59712 202748 59764
rect 204812 59712 204864 59764
rect 209412 59712 209464 59764
rect 209872 59712 209924 59764
rect 210792 59712 210844 59764
rect 213184 59712 213236 59764
rect 216588 59712 216640 59764
rect 218152 59712 218204 59764
rect 219256 59712 219308 59764
rect 221464 59712 221516 59764
rect 238576 59712 238628 59764
rect 240600 59712 240652 59764
rect 242716 59712 242768 59764
rect 244740 59712 244792 59764
rect 248328 59712 248380 59764
rect 249708 59712 249760 59764
rect 251824 59712 251876 59764
rect 253204 59712 253256 59764
rect 267740 59712 267792 59764
rect 269212 59712 269264 59764
rect 272708 59712 272760 59764
rect 274732 59712 274784 59764
rect 276848 59712 276900 59764
rect 278780 59712 278832 59764
rect 286784 59712 286836 59764
rect 288440 59712 288492 59764
rect 291844 59712 291896 59764
rect 294144 59712 294196 59764
rect 300124 59712 300176 59764
rect 303068 59712 303120 59764
rect 303436 59712 303488 59764
rect 305736 59712 305788 59764
rect 310704 59712 310756 59764
rect 312544 59712 312596 59764
rect 318432 59712 318484 59764
rect 320916 59712 320968 59764
rect 326712 59712 326764 59764
rect 329104 59712 329156 59764
rect 330852 59712 330904 59764
rect 331680 59712 331732 59764
rect 337568 59712 337620 59764
rect 340328 59712 340380 59764
rect 345020 59712 345072 59764
rect 347044 59712 347096 59764
rect 356704 59712 356756 59764
rect 359648 59712 359700 59764
rect 360844 59712 360896 59764
rect 363604 59712 363656 59764
rect 373816 59712 373868 59764
rect 375472 59712 375524 59764
rect 379980 59712 380032 59764
rect 380992 59712 381044 59764
rect 406568 59712 406620 59764
rect 408500 59712 408552 59764
rect 409052 59712 409104 59764
rect 410156 59712 410208 59764
rect 417608 59712 417660 59764
rect 419632 59712 419684 59764
rect 422116 59712 422168 59764
rect 423956 59712 424008 59764
rect 425704 59712 425756 59764
rect 428004 59712 428056 59764
rect 429844 59712 429896 59764
rect 432328 59712 432380 59764
rect 435824 59712 435876 59764
rect 438308 59712 438360 59764
rect 442356 59712 442408 59764
rect 445208 59712 445260 59764
rect 445668 59712 445720 59764
rect 447784 59712 447836 59764
rect 456524 59712 456576 59764
rect 458824 59712 458876 59764
rect 461492 59712 461544 59764
rect 462964 59712 463016 59764
rect 158352 59644 158404 59696
rect 159916 59644 159968 59696
rect 257344 59644 257396 59696
rect 258080 59644 258132 59696
rect 301780 59644 301832 59696
rect 304448 59644 304500 59696
rect 319260 59644 319312 59696
rect 320180 59644 320232 59696
rect 320824 59644 320876 59696
rect 322940 59644 322992 59696
rect 325056 59644 325108 59696
rect 327724 59644 327776 59696
rect 330944 59644 330996 59696
rect 333336 59644 333388 59696
rect 438216 59644 438268 59696
rect 440884 59644 440936 59696
rect 454776 59644 454828 59696
rect 457444 59644 457496 59696
rect 57244 59576 57296 59628
rect 62672 59576 62724 59628
rect 75736 59576 75788 59628
rect 77576 59576 77628 59628
rect 94504 59576 94556 59628
rect 96712 59576 96764 59628
rect 102784 59576 102836 59628
rect 105084 59576 105136 59628
rect 108304 59576 108356 59628
rect 110880 59576 110932 59628
rect 117964 59576 118016 59628
rect 119988 59576 120040 59628
rect 129004 59576 129056 59628
rect 131672 59576 131724 59628
rect 131764 59576 131816 59628
rect 134156 59576 134208 59628
rect 146208 59576 146260 59628
rect 147496 59576 147548 59628
rect 179328 59576 179380 59628
rect 180708 59576 180760 59628
rect 198556 59576 198608 59628
rect 200672 59576 200724 59628
rect 227628 59576 227680 59628
rect 228916 59576 228968 59628
rect 255964 59576 256016 59628
rect 257252 59576 257304 59628
rect 258724 59576 258776 59628
rect 260564 59576 260616 59628
rect 293500 59576 293552 59628
rect 295524 59576 295576 59628
rect 296812 59576 296864 59628
rect 298744 59576 298796 59628
rect 305920 59576 305972 59628
rect 307024 59576 307076 59628
rect 316592 59576 316644 59628
rect 318064 59576 318116 59628
rect 342352 59576 342404 59628
rect 344468 59576 344520 59628
rect 353392 59576 353444 59628
rect 354680 59576 354732 59628
rect 360108 59576 360160 59628
rect 361028 59576 361080 59628
rect 369032 59576 369084 59628
rect 369952 59576 370004 59628
rect 384120 59576 384172 59628
rect 385408 59576 385460 59628
rect 393320 59576 393372 59628
rect 394792 59576 394844 59628
rect 431776 59576 431828 59628
rect 433708 59576 433760 59628
rect 450636 59576 450688 59628
rect 451924 59576 451976 59628
rect 458180 59576 458232 59628
rect 460204 59576 460256 59628
rect 146944 59508 146996 59560
rect 149152 59508 149204 59560
rect 446404 59508 446456 59560
rect 448520 59508 448572 59560
rect 115388 59440 115440 59492
rect 117504 59440 117556 59492
rect 157064 59440 157116 59492
rect 157340 59440 157392 59492
rect 176292 59440 176344 59492
rect 178224 59440 178276 59492
rect 205272 59440 205324 59492
rect 207296 59440 207348 59492
rect 215116 59440 215168 59492
rect 215944 59440 215996 59492
rect 259000 59440 259052 59492
rect 260564 59440 260616 59492
rect 282644 59440 282696 59492
rect 284576 59440 284628 59492
rect 306748 59440 306800 59492
rect 307760 59440 307812 59492
rect 321744 59440 321796 59492
rect 323584 59440 323636 59492
rect 331772 59440 331824 59492
rect 333244 59440 333296 59492
rect 333428 59440 333480 59492
rect 336096 59440 336148 59492
rect 347504 59440 347556 59492
rect 349988 59440 350040 59492
rect 362500 59440 362552 59492
rect 364432 59440 364484 59492
rect 364800 59440 364852 59492
rect 365720 59440 365772 59492
rect 366640 59440 366692 59492
rect 368572 59440 368624 59492
rect 385776 59440 385828 59492
rect 388168 59440 388220 59492
rect 419080 59440 419132 59492
rect 421288 59440 421340 59492
rect 448152 59440 448204 59492
rect 450728 59440 450780 59492
rect 452292 59440 452344 59492
rect 454868 59440 454920 59492
rect 463148 59440 463200 59492
rect 465908 59440 465960 59492
rect 3424 59372 3476 59424
rect 57980 59372 58032 59424
rect 169484 59372 169536 59424
rect 171600 59372 171652 59424
rect 194416 59372 194468 59424
rect 196532 59372 196584 59424
rect 246672 59372 246724 59424
rect 248880 59372 248932 59424
rect 135996 59304 136048 59356
rect 137560 59304 137612 59356
rect 156972 59304 157024 59356
rect 160100 59304 160152 59356
rect 451280 59304 451332 59356
rect 453488 59304 453540 59356
rect 461492 59304 461544 59356
rect 463148 59304 463200 59356
rect 350632 58964 350684 59016
rect 352288 58964 352340 59016
rect 174544 58828 174596 58880
rect 234620 58828 234672 58880
rect 236000 58828 236052 58880
rect 280068 58828 280120 58880
rect 305644 58828 305696 58880
rect 401508 58828 401560 58880
rect 186320 58760 186372 58812
rect 268200 58760 268252 58812
rect 305828 58760 305880 58812
rect 342260 58760 342312 58812
rect 351736 58760 351788 58812
rect 538220 58760 538272 58812
rect 40040 58692 40092 58744
rect 67548 58692 67600 58744
rect 81348 58692 81400 58744
rect 89720 58692 89772 58744
rect 125600 58692 125652 58744
rect 146208 58692 146260 58744
rect 194600 58692 194652 58744
rect 376668 58692 376720 58744
rect 6920 58624 6972 58676
rect 60648 58624 60700 58676
rect 88340 58624 88392 58676
rect 131856 58624 131908 58676
rect 232780 58624 232832 58676
rect 483020 58624 483072 58676
rect 142804 58488 142856 58540
rect 144276 58488 144328 58540
rect 417608 58488 417660 58540
rect 418436 58488 418488 58540
rect 222200 57468 222252 57520
rect 277400 57468 277452 57520
rect 273260 57400 273312 57452
rect 394700 57400 394752 57452
rect 165620 57332 165672 57384
rect 262128 57332 262180 57384
rect 307760 57332 307812 57384
rect 346400 57332 346452 57384
rect 354680 57332 354732 57384
rect 545120 57332 545172 57384
rect 46940 57264 46992 57316
rect 68928 57264 68980 57316
rect 88064 57264 88116 57316
rect 118700 57264 118752 57316
rect 162860 57264 162912 57316
rect 369492 57264 369544 57316
rect 32404 57196 32456 57248
rect 91928 57196 91980 57248
rect 235264 57196 235316 57248
rect 494060 57196 494112 57248
rect 218060 56040 218112 56092
rect 278780 56040 278832 56092
rect 314660 56040 314712 56092
rect 371240 56040 371292 56092
rect 168380 55972 168432 56024
rect 262036 55972 262088 56024
rect 267740 55972 267792 56024
rect 287060 55972 287112 56024
rect 320180 55972 320232 56024
rect 398840 55972 398892 56024
rect 251180 55904 251232 55956
rect 389456 55904 389508 55956
rect 448520 55904 448572 55956
rect 489920 55904 489972 55956
rect 20720 55836 20772 55888
rect 63408 55836 63460 55888
rect 87512 55836 87564 55888
rect 121460 55836 121512 55888
rect 236920 55836 236972 55888
rect 500960 55836 501012 55888
rect 190460 54680 190512 54732
rect 271972 54680 272024 54732
rect 353944 54680 353996 54732
rect 412824 54680 412876 54732
rect 198740 54612 198792 54664
rect 379704 54612 379756 54664
rect 29000 54544 29052 54596
rect 64328 54544 64380 54596
rect 226156 54544 226208 54596
rect 465172 54544 465224 54596
rect 52460 54476 52512 54528
rect 96068 54476 96120 54528
rect 106280 54476 106332 54528
rect 136548 54476 136600 54528
rect 237288 54476 237340 54528
rect 512000 54476 512052 54528
rect 129740 53252 129792 53304
rect 253388 53252 253440 53304
rect 320824 53252 320876 53304
rect 408500 53252 408552 53304
rect 170404 53184 170456 53236
rect 372712 53184 372764 53236
rect 222016 53116 222068 53168
rect 451280 53116 451332 53168
rect 451924 53116 451976 53168
rect 503720 53116 503772 53168
rect 33140 53048 33192 53100
rect 64144 53048 64196 53100
rect 69020 53048 69072 53100
rect 100208 53048 100260 53100
rect 239956 53048 240008 53100
rect 514760 53048 514812 53100
rect 240140 51892 240192 51944
rect 282920 51892 282972 51944
rect 315304 51892 315356 51944
rect 374000 51892 374052 51944
rect 136640 51824 136692 51876
rect 254768 51824 254820 51876
rect 291200 51824 291252 51876
rect 401600 51824 401652 51876
rect 190276 51756 190328 51808
rect 316040 51756 316092 51808
rect 322940 51756 322992 51808
rect 407120 51756 407172 51808
rect 44180 51688 44232 51740
rect 66904 51688 66956 51740
rect 244188 51688 244240 51740
rect 543740 51688 543792 51740
rect 183560 50532 183612 50584
rect 270684 50532 270736 50584
rect 330576 50532 330628 50584
rect 409972 50532 410024 50584
rect 169760 50464 169812 50516
rect 372620 50464 372672 50516
rect 222108 50396 222160 50448
rect 448520 50396 448572 50448
rect 48320 50328 48372 50380
rect 95884 50328 95936 50380
rect 245476 50328 245528 50380
rect 547880 50328 547932 50380
rect 172520 49172 172572 49224
rect 268016 49172 268068 49224
rect 338764 49172 338816 49224
rect 412732 49172 412784 49224
rect 186964 49104 187016 49156
rect 376760 49104 376812 49156
rect 219256 49036 219308 49088
rect 440332 49036 440384 49088
rect 14464 48968 14516 49020
rect 87788 48968 87840 49020
rect 246856 48968 246908 49020
rect 554780 48968 554832 49020
rect 176660 47744 176712 47796
rect 267832 47744 267884 47796
rect 337476 47744 337528 47796
rect 470600 47744 470652 47796
rect 214564 47676 214616 47728
rect 383752 47676 383804 47728
rect 215116 47608 215168 47660
rect 423680 47608 423732 47660
rect 17960 47540 18012 47592
rect 89168 47540 89220 47592
rect 248328 47540 248380 47592
rect 561680 47540 561732 47592
rect 193220 46384 193272 46436
rect 271880 46384 271932 46436
rect 336096 46384 336148 46436
rect 459560 46384 459612 46436
rect 206836 46316 206888 46368
rect 387800 46316 387852 46368
rect 138020 46248 138072 46300
rect 365720 46248 365772 46300
rect 27620 46180 27672 46232
rect 90364 46180 90416 46232
rect 249616 46180 249668 46232
rect 564532 46180 564584 46232
rect 316868 45024 316920 45076
rect 378140 45024 378192 45076
rect 201500 44956 201552 45008
rect 274732 44956 274784 45008
rect 333428 44956 333480 45008
rect 448612 44956 448664 45008
rect 194324 44888 194376 44940
rect 333980 44888 334032 44940
rect 352564 44888 352616 44940
rect 414112 44888 414164 44940
rect 34520 44820 34572 44872
rect 91744 44820 91796 44872
rect 158536 44820 158588 44872
rect 182180 44820 182232 44872
rect 250996 44820 251048 44872
rect 572720 44820 572772 44872
rect 177856 43596 177908 43648
rect 263600 43596 263652 43648
rect 322940 43596 322992 43648
rect 408776 43596 408828 43648
rect 194508 43528 194560 43580
rect 331220 43528 331272 43580
rect 348608 43528 348660 43580
rect 516140 43528 516192 43580
rect 205640 43460 205692 43512
rect 380992 43460 381044 43512
rect 9680 43392 9732 43444
rect 113824 43392 113876 43444
rect 217876 43392 217928 43444
rect 430580 43392 430632 43444
rect 259460 42236 259512 42288
rect 393412 42236 393464 42288
rect 201316 42168 201368 42220
rect 362960 42168 363012 42220
rect 186136 42100 186188 42152
rect 295340 42100 295392 42152
rect 352840 42100 352892 42152
rect 534080 42100 534132 42152
rect 49700 42032 49752 42084
rect 122104 42032 122156 42084
rect 224776 42032 224828 42084
rect 462320 42032 462372 42084
rect 158720 40876 158772 40928
rect 258908 40876 258960 40928
rect 319628 40876 319680 40928
rect 389180 40876 389232 40928
rect 244280 40808 244332 40860
rect 390560 40808 390612 40860
rect 190092 40740 190144 40792
rect 313280 40740 313332 40792
rect 344468 40740 344520 40792
rect 495440 40740 495492 40792
rect 205456 40672 205508 40724
rect 376760 40672 376812 40724
rect 456064 40672 456116 40724
rect 521660 40672 521712 40724
rect 326344 39516 326396 39568
rect 420920 39516 420972 39568
rect 188896 39448 188948 39500
rect 309140 39448 309192 39500
rect 309784 39448 309836 39500
rect 405832 39448 405884 39500
rect 204168 39380 204220 39432
rect 374092 39380 374144 39432
rect 449164 39380 449216 39432
rect 492680 39380 492732 39432
rect 227628 39312 227680 39364
rect 473360 39312 473412 39364
rect 278044 38088 278096 38140
rect 397552 38088 397604 38140
rect 202696 38020 202748 38072
rect 369860 38020 369912 38072
rect 188712 37952 188764 38004
rect 306380 37952 306432 38004
rect 354036 37952 354088 38004
rect 540980 37952 541032 38004
rect 225972 37884 226024 37936
rect 469220 37884 469272 37936
rect 266360 36728 266412 36780
rect 396172 36728 396224 36780
rect 202512 36660 202564 36712
rect 365720 36660 365772 36712
rect 187608 36592 187660 36644
rect 302240 36592 302292 36644
rect 352656 36592 352708 36644
rect 531320 36592 531372 36644
rect 223488 36524 223540 36576
rect 455420 36524 455472 36576
rect 262220 35368 262272 35420
rect 394700 35368 394752 35420
rect 201132 35300 201184 35352
rect 358820 35300 358872 35352
rect 185952 35232 186004 35284
rect 299480 35232 299532 35284
rect 351184 35232 351236 35284
rect 527180 35232 527232 35284
rect 220728 35164 220780 35216
rect 444380 35164 444432 35216
rect 184756 33940 184808 33992
rect 292580 33940 292632 33992
rect 336096 33940 336148 33992
rect 411260 33940 411312 33992
rect 216680 33872 216732 33924
rect 383936 33872 383988 33924
rect 197176 33804 197228 33856
rect 340880 33804 340932 33856
rect 349988 33804 350040 33856
rect 520280 33804 520332 33856
rect 92480 33736 92532 33788
rect 131764 33736 131816 33788
rect 219072 33736 219124 33788
rect 437480 33736 437532 33788
rect 177672 32580 177724 32632
rect 259552 32580 259604 32632
rect 320916 32580 320968 32632
rect 396080 32580 396132 32632
rect 193036 32512 193088 32564
rect 324320 32512 324372 32564
rect 344284 32512 344336 32564
rect 498200 32512 498252 32564
rect 214932 32444 214984 32496
rect 419540 32444 419592 32496
rect 70400 32376 70452 32428
rect 127808 32376 127860 32428
rect 142160 32376 142212 32428
rect 367100 32376 367152 32428
rect 457628 32376 457680 32428
rect 528560 32376 528612 32428
rect 147680 31220 147732 31272
rect 257528 31220 257580 31272
rect 343640 31220 343692 31272
rect 414296 31220 414348 31272
rect 201592 31152 201644 31204
rect 380900 31152 380952 31204
rect 217692 31084 217744 31136
rect 433340 31084 433392 31136
rect 63500 31016 63552 31068
rect 125048 31016 125100 31068
rect 175188 31016 175240 31068
rect 249800 31016 249852 31068
rect 251088 31016 251140 31068
rect 575480 31016 575532 31068
rect 309876 29860 309928 29912
rect 349160 29860 349212 29912
rect 229100 29792 229152 29844
rect 280160 29792 280212 29844
rect 319444 29792 319496 29844
rect 391940 29792 391992 29844
rect 140780 29724 140832 29776
rect 254584 29724 254636 29776
rect 269120 29724 269172 29776
rect 396356 29724 396408 29776
rect 191748 29656 191800 29708
rect 320180 29656 320232 29708
rect 358176 29656 358228 29708
rect 416872 29656 416924 29708
rect 60740 29588 60792 29640
rect 124864 29588 124916 29640
rect 249432 29588 249484 29640
rect 568580 29588 568632 29640
rect 311900 28432 311952 28484
rect 405740 28432 405792 28484
rect 216588 28364 216640 28416
rect 426440 28364 426492 28416
rect 126980 28296 127032 28348
rect 363052 28296 363104 28348
rect 56600 28228 56652 28280
rect 123668 28228 123720 28280
rect 173624 28228 173676 28280
rect 245660 28228 245712 28280
rect 246672 28228 246724 28280
rect 557540 28228 557592 28280
rect 338856 27072 338908 27124
rect 473452 27072 473504 27124
rect 191840 27004 191892 27056
rect 378232 27004 378284 27056
rect 212448 26936 212500 26988
rect 408500 26936 408552 26988
rect 52552 26868 52604 26920
rect 123484 26868 123536 26920
rect 173808 26868 173860 26920
rect 242900 26868 242952 26920
rect 245292 26868 245344 26920
rect 550640 26868 550692 26920
rect 172428 25712 172480 25764
rect 238760 25712 238812 25764
rect 337384 25712 337436 25764
rect 466460 25712 466512 25764
rect 210976 25644 211028 25696
rect 401600 25644 401652 25696
rect 131120 25576 131172 25628
rect 364432 25576 364484 25628
rect 44272 25508 44324 25560
rect 94504 25508 94556 25560
rect 238576 25508 238628 25560
rect 523040 25508 523092 25560
rect 318064 24284 318116 24336
rect 385040 24284 385092 24336
rect 127072 24216 127124 24268
rect 251824 24216 251876 24268
rect 336004 24216 336056 24268
rect 463700 24216 463752 24268
rect 195888 24148 195940 24200
rect 338120 24148 338172 24200
rect 22100 24080 22152 24132
rect 88984 24080 89036 24132
rect 235908 24080 235960 24132
rect 507860 24080 507912 24132
rect 316684 22924 316736 22976
rect 382280 22924 382332 22976
rect 133880 22856 133932 22908
rect 253204 22856 253256 22908
rect 329840 22856 329892 22908
rect 410156 22856 410208 22908
rect 192852 22788 192904 22840
rect 327080 22788 327132 22840
rect 332048 22788 332100 22840
rect 445760 22788 445812 22840
rect 77300 22720 77352 22772
rect 102968 22720 103020 22772
rect 234252 22720 234304 22772
rect 505100 22720 505152 22772
rect 280160 21564 280212 21616
rect 398932 21564 398984 21616
rect 151820 21496 151872 21548
rect 257344 21496 257396 21548
rect 334624 21496 334676 21548
rect 456892 21496 456944 21548
rect 208308 21428 208360 21480
rect 390560 21428 390612 21480
rect 84200 21360 84252 21412
rect 104348 21360 104400 21412
rect 168104 21360 168156 21412
rect 220820 21360 220872 21412
rect 232964 21360 233016 21412
rect 498292 21360 498344 21412
rect 293960 20136 294012 20188
rect 401784 20136 401836 20188
rect 143540 20068 143592 20120
rect 255964 20068 256016 20120
rect 260840 20068 260892 20120
rect 288440 20068 288492 20120
rect 333244 20068 333296 20120
rect 452660 20068 452712 20120
rect 206652 20000 206704 20052
rect 383660 20000 383712 20052
rect 461768 20000 461820 20052
rect 542360 20000 542412 20052
rect 80060 19932 80112 19984
rect 102784 19932 102836 19984
rect 168288 19932 168340 19984
rect 218152 19932 218204 19984
rect 231768 19932 231820 19984
rect 490012 19932 490064 19984
rect 357440 18844 357492 18896
rect 417056 18844 417108 18896
rect 247040 18776 247092 18828
rect 284392 18776 284444 18828
rect 322204 18776 322256 18828
rect 403072 18776 403124 18828
rect 205272 18708 205324 18760
rect 380900 18708 380952 18760
rect 66260 18640 66312 18692
rect 100024 18640 100076 18692
rect 135260 18640 135312 18692
rect 364340 18640 364392 18692
rect 460204 18640 460256 18692
rect 539600 18640 539652 18692
rect 99380 18572 99432 18624
rect 133328 18572 133380 18624
rect 164056 18572 164108 18624
rect 202880 18572 202932 18624
rect 230204 18572 230256 18624
rect 487160 18572 487212 18624
rect 200028 17416 200080 17468
rect 356060 17416 356112 17468
rect 209780 17348 209832 17400
rect 382372 17348 382424 17400
rect 60832 17280 60884 17332
rect 71228 17280 71280 17332
rect 242992 17280 243044 17332
rect 284576 17280 284628 17332
rect 305736 17280 305788 17332
rect 332600 17280 332652 17332
rect 349804 17280 349856 17332
rect 523132 17280 523184 17332
rect 16580 17212 16632 17264
rect 61384 17212 61436 17264
rect 79876 17212 79928 17264
rect 93860 17212 93912 17264
rect 102140 17212 102192 17264
rect 108488 17212 108540 17264
rect 163872 17212 163924 17264
rect 200120 17212 200172 17264
rect 228824 17212 228876 17264
rect 480260 17212 480312 17264
rect 340972 16124 341024 16176
rect 412916 16124 412968 16176
rect 272432 16056 272484 16108
rect 291384 16056 291436 16108
rect 316224 16056 316276 16108
rect 407212 16056 407264 16108
rect 162768 15988 162820 16040
rect 196808 15988 196860 16040
rect 233424 15988 233476 16040
rect 281540 15988 281592 16040
rect 305552 15988 305604 16040
rect 404544 15988 404596 16040
rect 98184 15920 98236 15972
rect 107108 15920 107160 15972
rect 184572 15920 184624 15972
rect 288532 15920 288584 15972
rect 298100 15920 298152 15972
rect 402980 15920 403032 15972
rect 446588 15920 446640 15972
rect 482376 15920 482428 15972
rect 59360 15852 59412 15904
rect 98828 15852 98880 15904
rect 180248 15852 180300 15904
rect 269212 15852 269264 15904
rect 287152 15852 287204 15904
rect 400312 15852 400364 15904
rect 459008 15852 459060 15904
rect 536104 15852 536156 15904
rect 289820 15172 289872 15224
rect 295524 15172 295576 15224
rect 255872 14968 255924 15020
rect 393596 14968 393648 15020
rect 248420 14900 248472 14952
rect 392124 14900 392176 14952
rect 241704 14832 241756 14884
rect 389548 14832 389600 14884
rect 237656 14764 237708 14816
rect 389364 14764 389416 14816
rect 234712 14696 234764 14748
rect 387984 14696 388036 14748
rect 231032 14628 231084 14680
rect 388168 14628 388220 14680
rect 227536 14560 227588 14612
rect 386420 14560 386472 14612
rect 223580 14492 223632 14544
rect 385408 14492 385460 14544
rect 84016 14424 84068 14476
rect 114744 14424 114796 14476
rect 161296 14424 161348 14476
rect 193312 14424 193364 14476
rect 219992 14424 220044 14476
rect 385224 14424 385276 14476
rect 450728 14424 450780 14476
rect 497096 14424 497148 14476
rect 155408 13336 155460 13388
rect 258724 13336 258776 13388
rect 340328 13336 340380 13388
rect 478144 13336 478196 13388
rect 188528 13268 188580 13320
rect 376944 13268 376996 13320
rect 180984 13200 181036 13252
rect 375656 13200 375708 13252
rect 177856 13132 177908 13184
rect 375472 13132 375524 13184
rect 26240 13064 26292 13116
rect 62764 13064 62816 13116
rect 82728 13064 82780 13116
rect 108120 13064 108172 13116
rect 173900 13064 173952 13116
rect 374184 13064 374236 13116
rect 376024 13064 376076 13116
rect 418252 13064 418304 13116
rect 454868 13064 454920 13116
rect 514852 13064 514904 13116
rect 300308 12384 300360 12436
rect 307944 12384 307996 12436
rect 323584 12248 323636 12300
rect 410800 12248 410852 12300
rect 153016 12180 153068 12232
rect 157800 12180 157852 12232
rect 325148 12180 325200 12232
rect 414296 12180 414348 12232
rect 324964 12112 325016 12164
rect 417424 12112 417476 12164
rect 226340 12044 226392 12096
rect 280344 12044 280396 12096
rect 327724 12044 327776 12096
rect 423772 12044 423824 12096
rect 215300 11976 215352 12028
rect 277400 11976 277452 12028
rect 327908 11976 327960 12028
rect 427912 11976 427964 12028
rect 211712 11908 211764 11960
rect 276296 11908 276348 11960
rect 329104 11908 329156 11960
rect 432052 11908 432104 11960
rect 208584 11840 208636 11892
rect 276112 11840 276164 11892
rect 329288 11840 329340 11892
rect 434720 11840 434772 11892
rect 81256 11772 81308 11824
rect 100760 11772 100812 11824
rect 11888 11704 11940 11756
rect 57244 11704 57296 11756
rect 78128 11704 78180 11756
rect 129188 11772 129240 11824
rect 205088 11772 205140 11824
rect 274916 11772 274968 11824
rect 283104 11772 283156 11824
rect 294144 11772 294196 11824
rect 330484 11772 330536 11824
rect 439136 11772 439188 11824
rect 126980 11704 127032 11756
rect 128176 11704 128228 11756
rect 158352 11704 158404 11756
rect 178592 11704 178644 11756
rect 197912 11704 197964 11756
rect 273352 11704 273404 11756
rect 279056 11704 279108 11756
rect 292672 11704 292724 11756
rect 331864 11704 331916 11756
rect 442172 11704 442224 11756
rect 447784 11704 447836 11756
rect 486424 11704 486476 11756
rect 218060 11636 218112 11688
rect 219256 11636 219308 11688
rect 234620 11636 234672 11688
rect 235816 11636 235868 11688
rect 251272 10480 251324 10532
rect 285680 10480 285732 10532
rect 313924 10480 313976 10532
rect 367192 10480 367244 10532
rect 162032 10412 162084 10464
rect 260104 10412 260156 10464
rect 284300 10412 284352 10464
rect 400496 10412 400548 10464
rect 58440 10344 58492 10396
rect 71044 10344 71096 10396
rect 77116 10344 77168 10396
rect 86132 10344 86184 10396
rect 224592 10344 224644 10396
rect 459192 10412 459244 10464
rect 458824 10344 458876 10396
rect 532056 10344 532108 10396
rect 4804 10276 4856 10328
rect 58624 10276 58676 10328
rect 84108 10276 84160 10328
rect 110420 10276 110472 10328
rect 229008 10276 229060 10328
rect 476488 10276 476540 10328
rect 76932 9596 76984 9648
rect 83280 9596 83332 9648
rect 72608 9256 72660 9308
rect 73804 9256 73856 9308
rect 209596 9188 209648 9240
rect 395344 9188 395396 9240
rect 209412 9120 209464 9172
rect 398932 9120 398984 9172
rect 453304 9120 453356 9172
rect 507676 9120 507728 9172
rect 210792 9052 210844 9104
rect 406016 9052 406068 9104
rect 453488 9052 453540 9104
rect 511264 9052 511316 9104
rect 81072 8984 81124 9036
rect 104532 8984 104584 9036
rect 157064 8984 157116 9036
rect 175464 8984 175516 9036
rect 213552 8984 213604 9036
rect 413100 8984 413152 9036
rect 454684 8984 454736 9036
rect 518348 8984 518400 9036
rect 51356 8916 51408 8968
rect 68284 8916 68336 8968
rect 96252 8916 96304 8968
rect 133144 8916 133196 8968
rect 161112 8916 161164 8968
rect 189724 8916 189776 8968
rect 213736 8916 213788 8968
rect 416688 8916 416740 8968
rect 457444 8916 457496 8968
rect 525432 8916 525484 8968
rect 75736 8236 75788 8288
rect 79324 8236 79376 8288
rect 356704 8236 356756 8288
rect 361488 8236 361540 8288
rect 312728 8168 312780 8220
rect 364616 8168 364668 8220
rect 450544 8168 450596 8220
rect 500592 8168 500644 8220
rect 356888 8100 356940 8152
rect 549076 8100 549128 8152
rect 358084 8032 358136 8084
rect 359464 7964 359516 8016
rect 361488 8032 361540 8084
rect 552664 8032 552716 8084
rect 311164 7896 311216 7948
rect 354036 7896 354088 7948
rect 359648 7896 359700 7948
rect 361212 7896 361264 7948
rect 311348 7828 311400 7880
rect 357532 7828 357584 7880
rect 361028 7828 361080 7880
rect 556160 7964 556212 8016
rect 361396 7896 361448 7948
rect 559748 7896 559800 7948
rect 312544 7760 312596 7812
rect 361120 7760 361172 7812
rect 563244 7828 563296 7880
rect 566832 7760 566884 7812
rect 91560 7692 91612 7744
rect 105544 7692 105596 7744
rect 79692 7624 79744 7676
rect 97448 7624 97500 7676
rect 157248 7624 157300 7676
rect 171968 7692 172020 7744
rect 196992 7692 197044 7744
rect 345756 7692 345808 7744
rect 360844 7692 360896 7744
rect 570328 7692 570380 7744
rect 168380 7624 168432 7676
rect 169576 7624 169628 7676
rect 198372 7624 198424 7676
rect 349252 7624 349304 7676
rect 362224 7624 362276 7676
rect 573916 7624 573968 7676
rect 54944 7556 54996 7608
rect 69664 7556 69716 7608
rect 73804 7556 73856 7608
rect 101404 7556 101456 7608
rect 103336 7556 103388 7608
rect 134524 7556 134576 7608
rect 160008 7556 160060 7608
rect 186136 7556 186188 7608
rect 198556 7556 198608 7608
rect 352840 7556 352892 7608
rect 363604 7556 363656 7608
rect 577412 7556 577464 7608
rect 105728 7488 105780 7540
rect 108304 7488 108356 7540
rect 448612 7488 448664 7540
rect 449808 7488 449860 7540
rect 265348 6672 265400 6724
rect 288624 6672 288676 6724
rect 176476 6604 176528 6656
rect 253480 6604 253532 6656
rect 254676 6604 254728 6656
rect 287244 6604 287296 6656
rect 300124 6604 300176 6656
rect 311440 6604 311492 6656
rect 340144 6604 340196 6656
rect 481732 6604 481784 6656
rect 82084 6536 82136 6588
rect 129004 6536 129056 6588
rect 176292 6536 176344 6588
rect 257068 6536 257120 6588
rect 258264 6536 258316 6588
rect 287428 6536 287480 6588
rect 301504 6536 301556 6588
rect 315028 6536 315080 6588
rect 341708 6536 341760 6588
rect 485228 6536 485280 6588
rect 41880 6468 41932 6520
rect 93124 6468 93176 6520
rect 179328 6468 179380 6520
rect 267740 6468 267792 6520
rect 303068 6468 303120 6520
rect 318524 6468 318576 6520
rect 341524 6468 341576 6520
rect 488816 6468 488868 6520
rect 75000 6400 75052 6452
rect 127624 6400 127676 6452
rect 180708 6400 180760 6452
rect 271236 6400 271288 6452
rect 302884 6400 302936 6452
rect 322112 6400 322164 6452
rect 342996 6400 343048 6452
rect 492312 6400 492364 6452
rect 38384 6332 38436 6384
rect 93308 6332 93360 6384
rect 180616 6332 180668 6384
rect 274824 6332 274876 6384
rect 276020 6332 276072 6384
rect 291568 6332 291620 6384
rect 304448 6332 304500 6384
rect 325608 6332 325660 6384
rect 345664 6332 345716 6384
rect 502984 6332 503036 6384
rect 67916 6264 67968 6316
rect 126244 6264 126296 6316
rect 181812 6264 181864 6316
rect 278320 6264 278372 6316
rect 304264 6264 304316 6316
rect 329196 6264 329248 6316
rect 345848 6264 345900 6316
rect 506480 6264 506532 6316
rect 19432 6196 19484 6248
rect 115388 6196 115440 6248
rect 181996 6196 182048 6248
rect 281908 6196 281960 6248
rect 307024 6196 307076 6248
rect 336280 6196 336332 6248
rect 347044 6196 347096 6248
rect 510068 6196 510120 6248
rect 14740 6128 14792 6180
rect 115204 6128 115256 6180
rect 129372 6128 129424 6180
rect 145564 6128 145616 6180
rect 155868 6128 155920 6180
rect 168380 6128 168432 6180
rect 183468 6128 183520 6180
rect 285404 6128 285456 6180
rect 286600 6128 286652 6180
rect 294052 6128 294104 6180
rect 307208 6128 307260 6180
rect 339868 6128 339920 6180
rect 348424 6128 348476 6180
rect 513564 6128 513616 6180
rect 298744 5584 298796 5636
rect 304356 5584 304408 5636
rect 293684 5516 293736 5568
rect 295708 5516 295760 5568
rect 298928 5516 298980 5568
rect 300768 5516 300820 5568
rect 165436 5244 165488 5296
rect 207388 5108 207440 5160
rect 238392 5108 238444 5160
rect 519544 5108 519596 5160
rect 63224 5040 63276 5092
rect 98644 5040 98696 5092
rect 165252 5040 165304 5092
rect 210976 5040 211028 5092
rect 240048 5040 240100 5092
rect 526628 5040 526680 5092
rect 56048 4972 56100 5024
rect 97264 4972 97316 5024
rect 111616 4972 111668 5024
rect 116400 4972 116452 5024
rect 166908 4972 166960 5024
rect 214472 4972 214524 5024
rect 241336 4972 241388 5024
rect 530124 4972 530176 5024
rect 37188 4904 37240 4956
rect 65524 4904 65576 4956
rect 85672 4904 85724 4956
rect 130384 4904 130436 4956
rect 136456 4904 136508 4956
rect 148508 4904 148560 4956
rect 169668 4904 169720 4956
rect 225144 4904 225196 4956
rect 241152 4904 241204 4956
rect 533712 4904 533764 4956
rect 8760 4836 8812 4888
rect 87604 4836 87656 4888
rect 95148 4836 95200 4888
rect 106924 4836 106976 4888
rect 112996 4836 113048 4888
rect 119896 4836 119948 4888
rect 169392 4836 169444 4888
rect 228732 4836 228784 4888
rect 242532 4836 242584 4888
rect 537208 4836 537260 4888
rect 4068 4768 4120 4820
rect 86224 4768 86276 4820
rect 87972 4768 88024 4820
rect 104164 4768 104216 4820
rect 113088 4768 113140 4820
rect 123484 4768 123536 4820
rect 132960 4768 133012 4820
rect 146944 4768 146996 4820
rect 154304 4768 154356 4820
rect 164884 4768 164936 4820
rect 171048 4768 171100 4820
rect 232228 4768 232280 4820
rect 242716 4768 242768 4820
rect 540796 4768 540848 4820
rect 65524 4224 65576 4276
rect 72424 4224 72476 4276
rect 69112 4156 69164 4208
rect 72516 4156 72568 4208
rect 111432 4156 111484 4208
rect 112812 4156 112864 4208
rect 153108 4156 153160 4208
rect 154212 4156 154264 4208
rect 43076 4088 43128 4140
rect 120908 4088 120960 4140
rect 167184 4088 167236 4140
rect 170404 4088 170456 4140
rect 277124 4088 277176 4140
rect 278044 4088 278096 4140
rect 333888 4088 333940 4140
rect 336096 4088 336148 4140
rect 404820 4088 404872 4140
rect 428188 4088 428240 4140
rect 463148 4088 463200 4140
rect 550272 4088 550324 4140
rect 39580 4020 39632 4072
rect 119528 4020 119580 4072
rect 401324 4020 401376 4072
rect 428004 4020 428056 4072
rect 462964 4020 463016 4072
rect 553768 4020 553820 4072
rect 35992 3952 36044 4004
rect 119344 3952 119396 4004
rect 362316 3952 362368 4004
rect 376024 3952 376076 4004
rect 397736 3952 397788 4004
rect 426532 3952 426584 4004
rect 429660 3952 429712 4004
rect 433524 3952 433576 4004
rect 464344 3952 464396 4004
rect 557356 3952 557408 4004
rect 32496 3884 32548 3936
rect 117964 3884 118016 3936
rect 124680 3884 124732 3936
rect 140044 3884 140096 3936
rect 394240 3884 394292 3936
rect 425060 3884 425112 3936
rect 438124 3884 438176 3936
rect 447416 3884 447468 3936
rect 465908 3884 465960 3936
rect 560852 3884 560904 3936
rect 28908 3816 28960 3868
rect 116768 3816 116820 3868
rect 121092 3816 121144 3868
rect 138664 3816 138716 3868
rect 24216 3748 24268 3800
rect 116584 3748 116636 3800
rect 117596 3748 117648 3800
rect 137284 3748 137336 3800
rect 140044 3748 140096 3800
rect 148324 3748 148376 3800
rect 193220 3748 193272 3800
rect 194416 3748 194468 3800
rect 251180 3748 251232 3800
rect 252376 3748 252428 3800
rect 371424 3816 371476 3868
rect 390652 3816 390704 3868
rect 425152 3816 425204 3868
rect 439504 3816 439556 3868
rect 450912 3816 450964 3868
rect 465724 3816 465776 3868
rect 564440 3816 564492 3868
rect 25320 3680 25372 3732
rect 142804 3680 142856 3732
rect 160192 3680 160244 3732
rect 365812 3748 365864 3800
rect 418436 3748 418488 3800
rect 440884 3748 440936 3800
rect 454500 3748 454552 3800
rect 467288 3748 467340 3800
rect 568028 3748 568080 3800
rect 20628 3612 20680 3664
rect 141608 3612 141660 3664
rect 156604 3612 156656 3664
rect 369952 3680 370004 3732
rect 387156 3680 387208 3732
rect 424140 3680 424192 3732
rect 441068 3680 441120 3732
rect 458088 3680 458140 3732
rect 467104 3680 467156 3732
rect 571524 3680 571576 3732
rect 365628 3612 365680 3664
rect 368572 3612 368624 3664
rect 383568 3612 383620 3664
rect 423956 3612 424008 3664
rect 442264 3612 442316 3664
rect 461584 3612 461636 3664
rect 468484 3612 468536 3664
rect 575112 3612 575164 3664
rect 11152 3544 11204 3596
rect 2872 3476 2924 3528
rect 4804 3476 4856 3528
rect 13544 3476 13596 3528
rect 14464 3476 14516 3528
rect 15936 3544 15988 3596
rect 141424 3544 141476 3596
rect 160100 3544 160152 3596
rect 161296 3544 161348 3596
rect 161388 3544 161440 3596
rect 368480 3544 368532 3596
rect 379980 3544 380032 3596
rect 422300 3544 422352 3596
rect 442448 3544 442500 3596
rect 140228 3476 140280 3528
rect 143540 3476 143592 3528
rect 144736 3476 144788 3528
rect 149520 3476 149572 3528
rect 365628 3476 365680 3528
rect 365720 3476 365772 3528
rect 367008 3476 367060 3528
rect 374000 3476 374052 3528
rect 375288 3476 375340 3528
rect 376484 3476 376536 3528
rect 421104 3476 421156 3528
rect 423772 3476 423824 3528
rect 424968 3476 425020 3528
rect 6460 3408 6512 3460
rect 144368 3408 144420 3460
rect 145932 3408 145984 3460
rect 367284 3408 367336 3460
rect 372896 3408 372948 3460
rect 421288 3408 421340 3460
rect 422576 3408 422628 3460
rect 432144 3476 432196 3528
rect 440332 3476 440384 3528
rect 441528 3476 441580 3528
rect 426164 3408 426216 3460
rect 433708 3408 433760 3460
rect 31300 3340 31352 3392
rect 32404 3340 32456 3392
rect 46664 3340 46716 3392
rect 120724 3340 120776 3392
rect 153016 3340 153068 3392
rect 161388 3340 161440 3392
rect 213368 3340 213420 3392
rect 214564 3340 214616 3392
rect 301964 3340 302016 3392
rect 305644 3340 305696 3392
rect 309048 3340 309100 3392
rect 309876 3340 309928 3392
rect 316040 3340 316092 3392
rect 317328 3340 317380 3392
rect 357440 3340 357492 3392
rect 358728 3340 358780 3392
rect 390560 3340 390612 3392
rect 391848 3340 391900 3392
rect 398840 3340 398892 3392
rect 400128 3340 400180 3392
rect 408408 3340 408460 3392
rect 429200 3340 429252 3392
rect 436836 3340 436888 3392
rect 440332 3340 440384 3392
rect 445208 3544 445260 3596
rect 472256 3544 472308 3596
rect 472624 3544 472676 3596
rect 582196 3544 582248 3596
rect 443644 3408 443696 3460
rect 449164 3476 449216 3528
rect 465172 3476 465224 3528
rect 470140 3476 470192 3528
rect 578608 3476 578660 3528
rect 468668 3408 468720 3460
rect 471244 3408 471296 3460
rect 581000 3408 581052 3460
rect 449164 3340 449216 3392
rect 461676 3340 461728 3392
rect 546684 3340 546736 3392
rect 110512 3272 110564 3324
rect 135904 3272 135956 3324
rect 326804 3272 326856 3324
rect 330576 3272 330628 3324
rect 351644 3272 351696 3324
rect 353944 3272 353996 3324
rect 411904 3272 411956 3324
rect 429292 3272 429344 3324
rect 433248 3272 433300 3324
rect 434812 3272 434864 3324
rect 438308 3272 438360 3324
rect 443828 3272 443880 3324
rect 446404 3272 446456 3324
rect 479340 3272 479392 3324
rect 498200 3272 498252 3324
rect 499028 3272 499080 3324
rect 514760 3272 514812 3324
rect 515588 3272 515640 3324
rect 110420 3204 110472 3256
rect 111616 3204 111668 3256
rect 114008 3204 114060 3256
rect 137468 3204 137520 3256
rect 319720 3204 319772 3256
rect 320824 3204 320876 3256
rect 415492 3204 415544 3256
rect 430672 3204 430724 3256
rect 445116 3204 445168 3256
rect 475752 3204 475804 3256
rect 572 3136 624 3188
rect 3424 3136 3476 3188
rect 337476 3136 337528 3188
rect 338764 3136 338816 3188
rect 348056 3136 348108 3188
rect 352564 3136 352616 3188
rect 418988 3136 419040 3188
rect 432328 3136 432380 3188
rect 147128 3068 147180 3120
rect 149704 3068 149756 3120
rect 355232 3000 355284 3052
rect 358176 3000 358228 3052
rect 143540 2932 143592 2984
rect 149888 2932 149940 2984
rect 184940 2932 184992 2984
rect 186964 2932 187016 2984
rect 340880 1368 340932 1420
rect 342168 1368 342220 1420
rect 349160 1368 349212 1420
rect 350448 1368 350500 1420
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 57610 449304 57666 449313
rect 57610 449239 57666 449248
rect 57624 448594 57652 449239
rect 1400 448588 1452 448594
rect 1400 448530 1452 448536
rect 57612 448588 57664 448594
rect 57612 448530 57664 448536
rect 572 3188 624 3194
rect 572 3130 624 3136
rect 584 480 612 3130
rect 542 -960 654 480
rect 1412 354 1440 448530
rect 314292 59832 314344 59838
rect 64234 59800 64290 59809
rect 63408 59764 63460 59770
rect 64234 59735 64236 59744
rect 63408 59706 63460 59712
rect 64288 59735 64290 59744
rect 65338 59800 65394 59809
rect 68466 59800 68522 59809
rect 65338 59735 65394 59744
rect 67548 59764 67600 59770
rect 64236 59706 64288 59712
rect 62670 59664 62726 59673
rect 57244 59628 57296 59634
rect 62670 59599 62672 59608
rect 57244 59570 57296 59576
rect 62724 59599 62726 59608
rect 62672 59570 62724 59576
rect 3424 59424 3476 59430
rect 3424 59366 3476 59372
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2884 480 2912 3470
rect 3436 3194 3464 59366
rect 40040 58744 40092 58750
rect 40040 58686 40092 58692
rect 6920 58676 6972 58682
rect 6920 58618 6972 58624
rect 6932 16574 6960 58618
rect 32404 57248 32456 57254
rect 32404 57190 32456 57196
rect 20720 55888 20772 55894
rect 20720 55830 20772 55836
rect 14464 49020 14516 49026
rect 14464 48962 14516 48968
rect 9680 43444 9732 43450
rect 9680 43386 9732 43392
rect 6932 16546 7696 16574
rect 4804 10328 4856 10334
rect 4804 10270 4856 10276
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 4080 480 4108 4762
rect 4816 3534 4844 10270
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 5262 3360 5318 3369
rect 5262 3295 5318 3304
rect 5276 480 5304 3295
rect 6472 480 6500 3402
rect 7668 480 7696 16546
rect 8760 4888 8812 4894
rect 8760 4830 8812 4836
rect 8772 480 8800 4830
rect 1646 354 1758 480
rect 1412 326 1758 354
rect 1646 -960 1758 326
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 43386
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 11164 480 11192 3538
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 11900 354 11928 11698
rect 14476 3534 14504 48962
rect 17960 47592 18012 47598
rect 17960 47534 18012 47540
rect 16580 17264 16632 17270
rect 16580 17206 16632 17212
rect 16592 16574 16620 17206
rect 16592 16546 17080 16574
rect 14740 6180 14792 6186
rect 14740 6122 14792 6128
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 13556 480 13584 3470
rect 14752 480 14780 6122
rect 15936 3596 15988 3602
rect 15936 3538 15988 3544
rect 15948 480 15976 3538
rect 17052 480 17080 16546
rect 12318 354 12430 480
rect 11900 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 47534
rect 20732 16574 20760 55830
rect 29000 54596 29052 54602
rect 29000 54538 29052 54544
rect 27620 46232 27672 46238
rect 27620 46174 27672 46180
rect 22100 24132 22152 24138
rect 22100 24074 22152 24080
rect 22112 16574 22140 24074
rect 27632 16574 27660 46174
rect 29012 16574 29040 54538
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 27632 16546 27752 16574
rect 29012 16546 30144 16574
rect 19432 6248 19484 6254
rect 19432 6190 19484 6196
rect 19444 480 19472 6190
rect 20628 3664 20680 3670
rect 20628 3606 20680 3612
rect 20640 480 20668 3606
rect 21836 480 21864 16546
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 26240 13116 26292 13122
rect 26240 13058 26292 13064
rect 24216 3800 24268 3806
rect 24216 3742 24268 3748
rect 24228 480 24256 3742
rect 25320 3732 25372 3738
rect 25320 3674 25372 3680
rect 25332 480 25360 3674
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 13058
rect 27724 480 27752 16546
rect 28908 3868 28960 3874
rect 28908 3810 28960 3816
rect 28920 480 28948 3810
rect 30116 480 30144 16546
rect 32416 3398 32444 57190
rect 33140 53100 33192 53106
rect 33140 53042 33192 53048
rect 33152 16574 33180 53042
rect 34520 44872 34572 44878
rect 34520 44814 34572 44820
rect 33152 16546 33640 16574
rect 32496 3936 32548 3942
rect 32496 3878 32548 3884
rect 31300 3392 31352 3398
rect 31300 3334 31352 3340
rect 32404 3392 32456 3398
rect 32404 3334 32456 3340
rect 31312 480 31340 3334
rect 32508 1986 32536 3878
rect 32416 1958 32536 1986
rect 32416 480 32444 1958
rect 33612 480 33640 16546
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34532 354 34560 44814
rect 40052 16574 40080 58686
rect 46940 57316 46992 57322
rect 46940 57258 46992 57264
rect 44180 51740 44232 51746
rect 44180 51682 44232 51688
rect 40052 16546 40264 16574
rect 38384 6384 38436 6390
rect 38384 6326 38436 6332
rect 37188 4956 37240 4962
rect 37188 4898 37240 4904
rect 35992 4004 36044 4010
rect 35992 3946 36044 3952
rect 36004 480 36032 3946
rect 37200 480 37228 4898
rect 38396 480 38424 6326
rect 39580 4072 39632 4078
rect 39580 4014 39632 4020
rect 39592 480 39620 4014
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40236 354 40264 16546
rect 44192 6914 44220 51682
rect 44272 25560 44324 25566
rect 44272 25502 44324 25508
rect 44284 16574 44312 25502
rect 46952 16574 46980 57258
rect 52460 54528 52512 54534
rect 52460 54470 52512 54476
rect 48320 50380 48372 50386
rect 48320 50322 48372 50328
rect 48332 16574 48360 50322
rect 49700 42084 49752 42090
rect 49700 42026 49752 42032
rect 49712 16574 49740 42026
rect 44284 16546 45048 16574
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 44192 6886 44312 6914
rect 41880 6520 41932 6526
rect 41880 6462 41932 6468
rect 41892 480 41920 6462
rect 43076 4140 43128 4146
rect 43076 4082 43128 4088
rect 43088 480 43116 4082
rect 44284 480 44312 6886
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 46664 3392 46716 3398
rect 46664 3334 46716 3340
rect 46676 480 46704 3334
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 51356 8968 51408 8974
rect 51356 8910 51408 8916
rect 51368 480 51396 8910
rect 52472 6914 52500 54470
rect 56600 28280 56652 28286
rect 56600 28222 56652 28228
rect 52552 26920 52604 26926
rect 52552 26862 52604 26868
rect 52564 16574 52592 26862
rect 56612 16574 56640 28222
rect 52564 16546 53328 16574
rect 56612 16546 56824 16574
rect 52472 6886 52592 6914
rect 52564 480 52592 6886
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53300 354 53328 16546
rect 54944 7608 54996 7614
rect 54944 7550 54996 7556
rect 54956 480 54984 7550
rect 56048 5024 56100 5030
rect 56048 4966 56100 4972
rect 56060 480 56088 4966
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 57256 11762 57284 59570
rect 57978 59528 58034 59537
rect 57978 59463 58034 59472
rect 57992 59430 58020 59463
rect 57980 59424 58032 59430
rect 57980 59366 58032 59372
rect 58622 59392 58678 59401
rect 58622 59327 58678 59336
rect 62762 59392 62818 59401
rect 62762 59327 62818 59336
rect 57244 11756 57296 11762
rect 57244 11698 57296 11704
rect 58440 10396 58492 10402
rect 58440 10338 58492 10344
rect 58452 480 58480 10338
rect 58636 10334 58664 59327
rect 60646 59256 60702 59265
rect 60646 59191 60702 59200
rect 60660 58682 60688 59191
rect 61382 59120 61438 59129
rect 61382 59055 61438 59064
rect 60648 58676 60700 58682
rect 60648 58618 60700 58624
rect 60740 29640 60792 29646
rect 60740 29582 60792 29588
rect 59360 15904 59412 15910
rect 59360 15846 59412 15852
rect 58624 10328 58676 10334
rect 58624 10270 58676 10276
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 15846
rect 60752 6914 60780 29582
rect 60832 17332 60884 17338
rect 60832 17274 60884 17280
rect 60844 16574 60872 17274
rect 61396 17270 61424 59055
rect 61384 17264 61436 17270
rect 61384 17206 61436 17212
rect 60844 16546 61608 16574
rect 60752 6886 60872 6914
rect 60844 480 60872 6886
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61580 354 61608 16546
rect 62776 13122 62804 59327
rect 63420 55894 63448 59706
rect 64326 59664 64382 59673
rect 64326 59599 64382 59608
rect 64142 59256 64198 59265
rect 64142 59191 64198 59200
rect 63408 55888 63460 55894
rect 63408 55830 63460 55836
rect 64156 53106 64184 59191
rect 64340 54602 64368 59599
rect 65352 59537 65380 59735
rect 69294 59800 69350 59809
rect 68466 59735 68468 59744
rect 67548 59706 67600 59712
rect 68520 59735 68522 59744
rect 68928 59764 68980 59770
rect 68468 59706 68520 59712
rect 69294 59735 69350 59744
rect 70122 59800 70178 59809
rect 70122 59735 70124 59744
rect 68928 59706 68980 59712
rect 66810 59664 66866 59673
rect 66810 59599 66866 59608
rect 65338 59528 65394 59537
rect 65338 59463 65394 59472
rect 65522 59392 65578 59401
rect 65522 59327 65578 59336
rect 64328 54596 64380 54602
rect 64328 54538 64380 54544
rect 64144 53100 64196 53106
rect 64144 53042 64196 53048
rect 63500 31068 63552 31074
rect 63500 31010 63552 31016
rect 63512 16574 63540 31010
rect 63512 16546 64368 16574
rect 62764 13116 62816 13122
rect 62764 13058 62816 13064
rect 63224 5092 63276 5098
rect 63224 5034 63276 5040
rect 63236 480 63264 5034
rect 64340 480 64368 16546
rect 65536 4962 65564 59327
rect 66824 59265 66852 59599
rect 66902 59528 66958 59537
rect 66902 59463 66958 59472
rect 66810 59256 66866 59265
rect 66810 59191 66866 59200
rect 66916 51746 66944 59463
rect 67560 58750 67588 59706
rect 67638 59664 67694 59673
rect 67638 59599 67694 59608
rect 67652 59401 67680 59599
rect 67638 59392 67694 59401
rect 67638 59327 67694 59336
rect 68282 59392 68338 59401
rect 68282 59327 68338 59336
rect 67548 58744 67600 58750
rect 67548 58686 67600 58692
rect 66904 51740 66956 51746
rect 66904 51682 66956 51688
rect 66260 18692 66312 18698
rect 66260 18634 66312 18640
rect 66272 16574 66300 18634
rect 66272 16546 66760 16574
rect 65524 4956 65576 4962
rect 65524 4898 65576 4904
rect 65524 4276 65576 4282
rect 65524 4218 65576 4224
rect 65536 480 65564 4218
rect 66732 480 66760 16546
rect 68296 8974 68324 59327
rect 68940 57322 68968 59706
rect 69308 59537 69336 59735
rect 70176 59735 70178 59744
rect 71778 59800 71834 59809
rect 81346 59800 81402 59809
rect 71778 59735 71834 59744
rect 72700 59764 72752 59770
rect 70124 59706 70176 59712
rect 69294 59528 69350 59537
rect 69294 59463 69350 59472
rect 71042 59528 71098 59537
rect 71042 59463 71098 59472
rect 69662 59392 69718 59401
rect 69662 59327 69718 59336
rect 68928 57316 68980 57322
rect 68928 57258 68980 57264
rect 69020 53100 69072 53106
rect 69020 53042 69072 53048
rect 68284 8968 68336 8974
rect 68284 8910 68336 8916
rect 69032 6914 69060 53042
rect 69676 7614 69704 59327
rect 70400 32428 70452 32434
rect 70400 32370 70452 32376
rect 69664 7608 69716 7614
rect 69664 7550 69716 7556
rect 70412 6914 70440 32370
rect 71056 10402 71084 59463
rect 71792 59401 71820 59735
rect 72700 59706 72752 59712
rect 74632 59764 74684 59770
rect 74632 59706 74684 59712
rect 81072 59764 81124 59770
rect 81346 59735 81402 59744
rect 83462 59800 83518 59809
rect 87510 59800 87566 59809
rect 83462 59735 83464 59744
rect 81072 59706 81124 59712
rect 71778 59392 71834 59401
rect 71778 59327 71834 59336
rect 71226 59256 71282 59265
rect 71226 59191 71282 59200
rect 71240 17338 71268 59191
rect 72422 59120 72478 59129
rect 72422 59055 72478 59064
rect 71228 17332 71280 17338
rect 71228 17274 71280 17280
rect 71044 10396 71096 10402
rect 71044 10338 71096 10344
rect 69032 6886 69888 6914
rect 70412 6886 71544 6914
rect 67916 6316 67968 6322
rect 67916 6258 67968 6264
rect 67928 480 67956 6258
rect 69112 4208 69164 4214
rect 69112 4150 69164 4156
rect 69124 480 69152 4150
rect 61998 354 62110 480
rect 61580 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 69860 354 69888 6886
rect 71516 480 71544 6886
rect 72436 4282 72464 59055
rect 72712 45554 72740 59706
rect 74644 59673 74672 59706
rect 74630 59664 74686 59673
rect 77574 59664 77630 59673
rect 74630 59599 74686 59608
rect 75736 59628 75788 59634
rect 77574 59599 77576 59608
rect 75736 59570 75788 59576
rect 77628 59599 77630 59608
rect 79874 59664 79930 59673
rect 79874 59599 79930 59608
rect 77576 59570 77628 59576
rect 73802 59528 73858 59537
rect 73802 59463 73858 59472
rect 72620 45526 72740 45554
rect 72620 16574 72648 45526
rect 72528 16546 72648 16574
rect 72424 4276 72476 4282
rect 72424 4218 72476 4224
rect 72528 4214 72556 16546
rect 73816 9314 73844 59463
rect 75550 59392 75606 59401
rect 75550 59327 75606 59336
rect 72608 9308 72660 9314
rect 72608 9250 72660 9256
rect 73804 9308 73856 9314
rect 73804 9250 73856 9256
rect 72516 4208 72568 4214
rect 72516 4150 72568 4156
rect 72620 480 72648 9250
rect 73804 7608 73856 7614
rect 73804 7550 73856 7556
rect 73816 480 73844 7550
rect 75564 6914 75592 59327
rect 75748 8294 75776 59570
rect 76930 59528 76986 59537
rect 76930 59463 76986 59472
rect 76944 9654 76972 59463
rect 77114 59392 77170 59401
rect 77114 59327 77170 59336
rect 79690 59392 79746 59401
rect 79690 59327 79746 59336
rect 77128 10402 77156 59327
rect 77300 22772 77352 22778
rect 77300 22714 77352 22720
rect 77312 16574 77340 22714
rect 77312 16546 77432 16574
rect 77116 10396 77168 10402
rect 77116 10338 77168 10344
rect 76932 9648 76984 9654
rect 76932 9590 76984 9596
rect 75736 8288 75788 8294
rect 75736 8230 75788 8236
rect 75564 6886 75868 6914
rect 75000 6452 75052 6458
rect 75000 6394 75052 6400
rect 75012 480 75040 6394
rect 75840 4162 75868 6886
rect 75840 4134 75960 4162
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 75932 354 75960 4134
rect 77404 480 77432 16546
rect 78128 11756 78180 11762
rect 78128 11698 78180 11704
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 11698
rect 79324 8288 79376 8294
rect 79324 8230 79376 8236
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 79336 354 79364 8230
rect 79704 7682 79732 59327
rect 79888 17270 79916 59599
rect 80060 19984 80112 19990
rect 80060 19926 80112 19932
rect 79876 17264 79928 17270
rect 79876 17206 79928 17212
rect 80072 16574 80100 19926
rect 80072 16546 80928 16574
rect 79692 7676 79744 7682
rect 79692 7618 79744 7624
rect 80900 480 80928 16546
rect 81084 9042 81112 59706
rect 81254 59528 81310 59537
rect 81254 59463 81310 59472
rect 81268 11830 81296 59463
rect 81360 58750 81388 59735
rect 83516 59735 83518 59744
rect 86224 59764 86276 59770
rect 83464 59706 83516 59712
rect 87510 59735 87566 59744
rect 88430 59800 88486 59809
rect 91742 59800 91798 59809
rect 88430 59735 88432 59744
rect 86224 59706 86276 59712
rect 81806 59664 81862 59673
rect 81806 59599 81862 59608
rect 81820 59401 81848 59599
rect 84106 59528 84162 59537
rect 84106 59463 84162 59472
rect 81806 59392 81862 59401
rect 81806 59327 81862 59336
rect 82726 59392 82782 59401
rect 82726 59327 82782 59336
rect 84014 59392 84070 59401
rect 84014 59327 84070 59336
rect 81348 58744 81400 58750
rect 81348 58686 81400 58692
rect 82740 13122 82768 59327
rect 84028 14482 84056 59327
rect 84016 14476 84068 14482
rect 84016 14418 84068 14424
rect 82728 13116 82780 13122
rect 82728 13058 82780 13064
rect 81256 11824 81308 11830
rect 81256 11766 81308 11772
rect 84120 10334 84148 59463
rect 84200 21412 84252 21418
rect 84200 21354 84252 21360
rect 84108 10328 84160 10334
rect 84108 10270 84160 10276
rect 83280 9648 83332 9654
rect 83280 9590 83332 9596
rect 81072 9036 81124 9042
rect 81072 8978 81124 8984
rect 82084 6588 82136 6594
rect 82084 6530 82136 6536
rect 82096 480 82124 6530
rect 83292 480 83320 9590
rect 79662 354 79774 480
rect 79336 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84212 354 84240 21354
rect 86132 10396 86184 10402
rect 86132 10338 86184 10344
rect 85672 4956 85724 4962
rect 85672 4898 85724 4904
rect 85684 480 85712 4898
rect 86144 490 86172 10338
rect 86236 4826 86264 59706
rect 87524 55894 87552 59735
rect 88484 59735 88486 59744
rect 88984 59764 89036 59770
rect 88432 59706 88484 59712
rect 98366 59800 98422 59809
rect 91742 59735 91744 59744
rect 88984 59706 89036 59712
rect 91796 59735 91798 59744
rect 96068 59764 96120 59770
rect 91744 59706 91796 59712
rect 100850 59800 100906 59809
rect 98366 59735 98368 59744
rect 96068 59706 96120 59712
rect 98420 59735 98422 59744
rect 98644 59764 98696 59770
rect 98368 59706 98420 59712
rect 100850 59735 100852 59744
rect 98644 59706 98696 59712
rect 100904 59735 100906 59744
rect 102506 59800 102562 59809
rect 102506 59735 102562 59744
rect 103426 59800 103482 59809
rect 103426 59735 103482 59744
rect 107198 59800 107254 59809
rect 107474 59800 107530 59809
rect 107254 59758 107474 59786
rect 107198 59735 107254 59744
rect 107474 59735 107530 59744
rect 111798 59800 111854 59809
rect 115018 59800 115074 59809
rect 111798 59735 111854 59744
rect 113088 59764 113140 59770
rect 100852 59706 100904 59712
rect 88430 59664 88486 59673
rect 87616 59622 88430 59650
rect 87512 55888 87564 55894
rect 87512 55830 87564 55836
rect 87616 4894 87644 59622
rect 88430 59599 88486 59608
rect 88062 59528 88118 59537
rect 88062 59463 88118 59472
rect 87786 59392 87842 59401
rect 87786 59327 87842 59336
rect 87800 49026 87828 59327
rect 88076 57322 88104 59463
rect 88340 58676 88392 58682
rect 88340 58618 88392 58624
rect 88064 57316 88116 57322
rect 88064 57258 88116 57264
rect 87788 49020 87840 49026
rect 87788 48962 87840 48968
rect 88352 16574 88380 58618
rect 88996 24138 89024 59706
rect 90086 59664 90142 59673
rect 93398 59664 93454 59673
rect 90086 59599 90142 59608
rect 93136 59622 93398 59650
rect 89166 59528 89222 59537
rect 89166 59463 89222 59472
rect 89180 47598 89208 59463
rect 90100 59401 90128 59599
rect 93136 59537 93164 59622
rect 93398 59599 93454 59608
rect 94318 59664 94374 59673
rect 95974 59664 96030 59673
rect 94318 59599 94374 59608
rect 94504 59628 94556 59634
rect 91926 59528 91982 59537
rect 91926 59463 91982 59472
rect 93122 59528 93178 59537
rect 93122 59463 93178 59472
rect 93306 59528 93362 59537
rect 93306 59463 93362 59472
rect 90086 59392 90142 59401
rect 90086 59327 90142 59336
rect 90362 59392 90418 59401
rect 90362 59327 90418 59336
rect 91834 59392 91890 59401
rect 91834 59327 91890 59336
rect 89720 58744 89772 58750
rect 89720 58686 89772 58692
rect 89168 47592 89220 47598
rect 89168 47534 89220 47540
rect 88984 24132 89036 24138
rect 88984 24074 89036 24080
rect 89732 16574 89760 58686
rect 90376 46238 90404 59327
rect 90364 46232 90416 46238
rect 90364 46174 90416 46180
rect 91848 45554 91876 59327
rect 91940 57254 91968 59463
rect 93122 59256 93178 59265
rect 93122 59191 93178 59200
rect 91928 57248 91980 57254
rect 91928 57190 91980 57196
rect 91756 45526 91876 45554
rect 91756 44878 91784 45526
rect 91744 44872 91796 44878
rect 91744 44814 91796 44820
rect 92480 33788 92532 33794
rect 92480 33730 92532 33736
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 87604 4888 87656 4894
rect 87604 4830 87656 4836
rect 86224 4820 86276 4826
rect 86224 4762 86276 4768
rect 87972 4820 88024 4826
rect 87972 4762 88024 4768
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86144 462 86540 490
rect 87984 480 88012 4762
rect 89180 480 89208 16546
rect 86512 354 86540 462
rect 86838 354 86950 480
rect 86512 326 86950 354
rect 86838 -960 86950 326
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91560 7744 91612 7750
rect 91560 7686 91612 7692
rect 91572 480 91600 7686
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 33730
rect 93136 6526 93164 59191
rect 93124 6520 93176 6526
rect 93124 6462 93176 6468
rect 93320 6390 93348 59463
rect 94332 59401 94360 59599
rect 95974 59599 96030 59608
rect 94504 59570 94556 59576
rect 94318 59392 94374 59401
rect 94318 59327 94374 59336
rect 94516 25566 94544 59570
rect 95882 59528 95938 59537
rect 95882 59463 95938 59472
rect 95896 50386 95924 59463
rect 95988 59401 96016 59599
rect 95974 59392 96030 59401
rect 95974 59327 96030 59336
rect 96080 54534 96108 59706
rect 96710 59664 96766 59673
rect 96710 59599 96712 59608
rect 96764 59599 96766 59608
rect 96712 59570 96764 59576
rect 97262 59392 97318 59401
rect 97262 59327 97318 59336
rect 96068 54528 96120 54534
rect 96068 54470 96120 54476
rect 95884 50380 95936 50386
rect 95884 50322 95936 50328
rect 94504 25560 94556 25566
rect 94504 25502 94556 25508
rect 93860 17264 93912 17270
rect 93860 17206 93912 17212
rect 93872 16574 93900 17206
rect 93872 16546 93992 16574
rect 93308 6384 93360 6390
rect 93308 6326 93360 6332
rect 93964 480 93992 16546
rect 96252 8968 96304 8974
rect 96252 8910 96304 8916
rect 95148 4888 95200 4894
rect 95148 4830 95200 4836
rect 95160 480 95188 4830
rect 96264 480 96292 8910
rect 97276 5030 97304 59327
rect 98184 15972 98236 15978
rect 98184 15914 98236 15920
rect 97448 7676 97500 7682
rect 97448 7618 97500 7624
rect 97264 5024 97316 5030
rect 97264 4966 97316 4972
rect 97460 480 97488 7618
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98196 354 98224 15914
rect 98656 5098 98684 59706
rect 98826 59528 98882 59537
rect 98826 59463 98882 59472
rect 101402 59528 101458 59537
rect 101402 59463 101458 59472
rect 98840 15910 98868 59463
rect 100022 59392 100078 59401
rect 100022 59327 100078 59336
rect 100036 18698 100064 59327
rect 100206 59256 100262 59265
rect 100206 59191 100262 59200
rect 100220 53106 100248 59191
rect 100208 53100 100260 53106
rect 100208 53042 100260 53048
rect 100024 18692 100076 18698
rect 100024 18634 100076 18640
rect 99380 18624 99432 18630
rect 99380 18566 99432 18572
rect 99392 16574 99420 18566
rect 99392 16546 99880 16574
rect 98828 15904 98880 15910
rect 98828 15846 98880 15852
rect 98644 5092 98696 5098
rect 98644 5034 98696 5040
rect 99852 480 99880 16546
rect 100760 11824 100812 11830
rect 100760 11766 100812 11772
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 11766
rect 101416 7614 101444 59463
rect 102520 59401 102548 59735
rect 102966 59664 103022 59673
rect 102784 59628 102836 59634
rect 102966 59599 103022 59608
rect 102784 59570 102836 59576
rect 102506 59392 102562 59401
rect 102506 59327 102562 59336
rect 102796 19990 102824 59570
rect 102980 22778 103008 59599
rect 103440 59537 103468 59735
rect 105082 59664 105138 59673
rect 107566 59664 107622 59673
rect 105082 59599 105084 59608
rect 105136 59599 105138 59608
rect 106936 59622 107566 59650
rect 105084 59570 105136 59576
rect 103426 59528 103482 59537
rect 103426 59463 103482 59472
rect 104346 59528 104402 59537
rect 104346 59463 104402 59472
rect 104162 59392 104218 59401
rect 104162 59327 104218 59336
rect 102968 22772 103020 22778
rect 102968 22714 103020 22720
rect 102784 19984 102836 19990
rect 102784 19926 102836 19932
rect 102140 17264 102192 17270
rect 102140 17206 102192 17212
rect 102152 16574 102180 17206
rect 102152 16546 102272 16574
rect 101404 7608 101456 7614
rect 101404 7550 101456 7556
rect 102244 480 102272 16546
rect 103336 7608 103388 7614
rect 103336 7550 103388 7556
rect 103348 480 103376 7550
rect 104176 4826 104204 59327
rect 104360 21418 104388 59463
rect 105542 59392 105598 59401
rect 105542 59327 105598 59336
rect 104348 21412 104400 21418
rect 104348 21354 104400 21360
rect 104532 9036 104584 9042
rect 104532 8978 104584 8984
rect 104164 4820 104216 4826
rect 104164 4762 104216 4768
rect 104544 480 104572 8978
rect 105556 7750 105584 59327
rect 106280 54528 106332 54534
rect 106280 54470 106332 54476
rect 106292 16574 106320 54470
rect 106292 16546 106504 16574
rect 105544 7744 105596 7750
rect 105544 7686 105596 7692
rect 105728 7540 105780 7546
rect 105728 7482 105780 7488
rect 105740 480 105768 7482
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 106936 4894 106964 59622
rect 109222 59664 109278 59673
rect 107566 59599 107622 59608
rect 108304 59628 108356 59634
rect 108304 59570 108356 59576
rect 108868 59622 109222 59650
rect 107106 59392 107162 59401
rect 107106 59327 107162 59336
rect 107120 15978 107148 59327
rect 107108 15972 107160 15978
rect 107108 15914 107160 15920
rect 108120 13116 108172 13122
rect 108120 13058 108172 13064
rect 106924 4888 106976 4894
rect 106924 4830 106976 4836
rect 108132 480 108160 13058
rect 108316 7546 108344 59570
rect 108486 59528 108542 59537
rect 108486 59463 108542 59472
rect 108500 17270 108528 59463
rect 108868 59401 108896 59622
rect 109222 59599 109278 59608
rect 110878 59664 110934 59673
rect 111706 59664 111762 59673
rect 110878 59599 110880 59608
rect 110932 59599 110934 59608
rect 111444 59622 111706 59650
rect 110880 59570 110932 59576
rect 108854 59392 108910 59401
rect 108854 59327 108910 59336
rect 109038 59392 109094 59401
rect 109038 59327 109094 59336
rect 108488 17264 108540 17270
rect 108488 17206 108540 17212
rect 108304 7540 108356 7546
rect 108304 7482 108356 7488
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109052 354 109080 59327
rect 110420 10328 110472 10334
rect 110420 10270 110472 10276
rect 110432 3262 110460 10270
rect 111444 4214 111472 59622
rect 111706 59599 111762 59608
rect 111812 59537 111840 59735
rect 115018 59735 115020 59744
rect 113088 59706 113140 59712
rect 115072 59735 115074 59744
rect 121642 59800 121698 59809
rect 123298 59800 123354 59809
rect 121642 59735 121698 59744
rect 122748 59764 122800 59770
rect 115020 59706 115072 59712
rect 111798 59528 111854 59537
rect 111798 59463 111854 59472
rect 112994 59528 113050 59537
rect 112994 59463 113050 59472
rect 111614 59392 111670 59401
rect 111614 59327 111670 59336
rect 111628 5030 111656 59327
rect 111616 5024 111668 5030
rect 111616 4966 111668 4972
rect 113008 4894 113036 59463
rect 112996 4888 113048 4894
rect 112996 4830 113048 4836
rect 113100 4826 113128 59706
rect 113546 59664 113602 59673
rect 119986 59664 120042 59673
rect 113546 59599 113602 59608
rect 117964 59628 118016 59634
rect 113560 59401 113588 59599
rect 119986 59599 119988 59608
rect 117964 59570 118016 59576
rect 120040 59599 120042 59608
rect 120722 59664 120778 59673
rect 120722 59599 120778 59608
rect 119988 59570 120040 59576
rect 115202 59528 115258 59537
rect 117502 59528 117558 59537
rect 115202 59463 115258 59472
rect 115388 59492 115440 59498
rect 113546 59392 113602 59401
rect 113546 59327 113602 59336
rect 114190 59392 114246 59401
rect 114190 59327 114246 59336
rect 114204 45554 114232 59327
rect 113836 45526 114232 45554
rect 113836 43450 113864 45526
rect 113824 43444 113876 43450
rect 113824 43386 113876 43392
rect 114744 14476 114796 14482
rect 114744 14418 114796 14424
rect 113088 4820 113140 4826
rect 113088 4762 113140 4768
rect 111432 4208 111484 4214
rect 111432 4150 111484 4156
rect 112812 4208 112864 4214
rect 112812 4150 112864 4156
rect 110512 3324 110564 3330
rect 110512 3266 110564 3272
rect 110420 3256 110472 3262
rect 110420 3198 110472 3204
rect 110524 480 110552 3266
rect 111616 3256 111668 3262
rect 111616 3198 111668 3204
rect 111628 480 111656 3198
rect 112824 480 112852 4150
rect 114008 3256 114060 3262
rect 114008 3198 114060 3204
rect 114020 480 114048 3198
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 114756 354 114784 14418
rect 115216 6186 115244 59463
rect 117502 59463 117504 59472
rect 115388 59434 115440 59440
rect 117556 59463 117558 59472
rect 117504 59434 117556 59440
rect 115400 6254 115428 59434
rect 116582 59392 116638 59401
rect 116582 59327 116638 59336
rect 115388 6248 115440 6254
rect 115388 6190 115440 6196
rect 115204 6180 115256 6186
rect 115204 6122 115256 6128
rect 116400 5024 116452 5030
rect 116400 4966 116452 4972
rect 116412 480 116440 4966
rect 116596 3806 116624 59327
rect 116766 59256 116822 59265
rect 116766 59191 116822 59200
rect 116780 3874 116808 59191
rect 117976 3942 118004 59570
rect 119986 59528 120042 59537
rect 119356 59486 119986 59514
rect 118700 57316 118752 57322
rect 118700 57258 118752 57264
rect 118712 16574 118740 57258
rect 118712 16546 118832 16574
rect 117964 3936 118016 3942
rect 117964 3878 118016 3884
rect 116768 3868 116820 3874
rect 116768 3810 116820 3816
rect 116584 3800 116636 3806
rect 116584 3742 116636 3748
rect 117596 3800 117648 3806
rect 117596 3742 117648 3748
rect 117608 480 117636 3742
rect 118804 480 118832 16546
rect 119356 4010 119384 59486
rect 119986 59463 120042 59472
rect 119526 59392 119582 59401
rect 119526 59327 119582 59336
rect 119540 4078 119568 59327
rect 119896 4888 119948 4894
rect 119896 4830 119948 4836
rect 119528 4072 119580 4078
rect 119528 4014 119580 4020
rect 119344 4004 119396 4010
rect 119344 3946 119396 3952
rect 119908 480 119936 4830
rect 120736 3398 120764 59599
rect 120906 59528 120962 59537
rect 120906 59463 120962 59472
rect 120920 4146 120948 59463
rect 121656 59401 121684 59735
rect 123298 59735 123300 59744
rect 122748 59706 122800 59712
rect 123352 59735 123354 59744
rect 124218 59800 124274 59809
rect 127530 59800 127586 59809
rect 124218 59735 124274 59744
rect 125140 59764 125192 59770
rect 123300 59706 123352 59712
rect 122760 59673 122788 59706
rect 122746 59664 122802 59673
rect 122746 59599 122802 59608
rect 123482 59664 123538 59673
rect 123482 59599 123538 59608
rect 121642 59392 121698 59401
rect 121642 59327 121698 59336
rect 122102 59392 122158 59401
rect 122102 59327 122158 59336
rect 121460 55888 121512 55894
rect 121460 55830 121512 55836
rect 121472 16574 121500 55830
rect 122116 42090 122144 59327
rect 122104 42084 122156 42090
rect 122104 42026 122156 42032
rect 123496 26926 123524 59599
rect 124232 59401 124260 59735
rect 136638 59800 136694 59809
rect 127530 59735 127532 59744
rect 125140 59706 125192 59712
rect 127584 59735 127586 59744
rect 134524 59764 134576 59770
rect 127532 59706 127584 59712
rect 136638 59735 136640 59744
rect 134524 59706 134576 59712
rect 136692 59735 136694 59744
rect 139214 59800 139270 59809
rect 139214 59735 139270 59744
rect 139950 59800 140006 59809
rect 141698 59800 141754 59809
rect 139950 59735 140006 59744
rect 140228 59764 140280 59770
rect 136640 59706 136692 59712
rect 125046 59528 125102 59537
rect 124876 59486 125046 59514
rect 124218 59392 124274 59401
rect 124218 59327 124274 59336
rect 123666 59256 123722 59265
rect 123666 59191 123722 59200
rect 123680 28286 123708 59191
rect 124876 29646 124904 59486
rect 125046 59463 125102 59472
rect 125152 45554 125180 59706
rect 125874 59664 125930 59673
rect 131670 59664 131726 59673
rect 125874 59599 125930 59608
rect 129004 59628 129056 59634
rect 125888 59401 125916 59599
rect 134154 59664 134210 59673
rect 131670 59599 131672 59608
rect 129004 59570 129056 59576
rect 131724 59599 131726 59608
rect 131764 59628 131816 59634
rect 131672 59570 131724 59576
rect 134154 59599 134156 59608
rect 131764 59570 131816 59576
rect 134208 59599 134210 59608
rect 134156 59570 134208 59576
rect 128358 59528 128414 59537
rect 127820 59486 128358 59514
rect 125874 59392 125930 59401
rect 125874 59327 125930 59336
rect 126242 59392 126298 59401
rect 126242 59327 126298 59336
rect 127714 59392 127770 59401
rect 127714 59327 127770 59336
rect 125600 58744 125652 58750
rect 125600 58686 125652 58692
rect 125060 45526 125180 45554
rect 125060 31074 125088 45526
rect 125048 31068 125100 31074
rect 125048 31010 125100 31016
rect 124864 29640 124916 29646
rect 124864 29582 124916 29588
rect 123668 28280 123720 28286
rect 123668 28222 123720 28228
rect 123484 26920 123536 26926
rect 123484 26862 123536 26868
rect 121472 16546 122328 16574
rect 120908 4140 120960 4146
rect 120908 4082 120960 4088
rect 121092 3868 121144 3874
rect 121092 3810 121144 3816
rect 120724 3392 120776 3398
rect 120724 3334 120776 3340
rect 121104 480 121132 3810
rect 122300 480 122328 16546
rect 123484 4820 123536 4826
rect 123484 4762 123536 4768
rect 123496 480 123524 4762
rect 124680 3936 124732 3942
rect 124680 3878 124732 3884
rect 124692 480 124720 3878
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125612 354 125640 58686
rect 126256 6322 126284 59327
rect 127728 45554 127756 59327
rect 127636 45526 127756 45554
rect 126980 28348 127032 28354
rect 126980 28290 127032 28296
rect 126992 11762 127020 28290
rect 127072 24268 127124 24274
rect 127072 24210 127124 24216
rect 126980 11756 127032 11762
rect 126980 11698 127032 11704
rect 127084 6914 127112 24210
rect 126992 6886 127112 6914
rect 126244 6316 126296 6322
rect 126244 6258 126296 6264
rect 126992 480 127020 6886
rect 127636 6458 127664 45526
rect 127820 32434 127848 59486
rect 128358 59463 128414 59472
rect 127808 32428 127860 32434
rect 127808 32370 127860 32376
rect 128176 11756 128228 11762
rect 128176 11698 128228 11704
rect 127624 6452 127676 6458
rect 127624 6394 127676 6400
rect 128188 480 128216 11698
rect 129016 6594 129044 59570
rect 129186 59256 129242 59265
rect 129186 59191 129242 59200
rect 129200 11830 129228 59191
rect 130382 59120 130438 59129
rect 130382 59055 130438 59064
rect 129740 53304 129792 53310
rect 129740 53246 129792 53252
rect 129752 16574 129780 53246
rect 129752 16546 130332 16574
rect 129188 11824 129240 11830
rect 129188 11766 129240 11772
rect 129004 6588 129056 6594
rect 129004 6530 129056 6536
rect 129372 6180 129424 6186
rect 129372 6122 129424 6128
rect 129384 480 129412 6122
rect 130304 3482 130332 16546
rect 130396 4962 130424 59055
rect 131776 33794 131804 59570
rect 133142 59528 133198 59537
rect 133142 59463 133198 59472
rect 131854 59392 131910 59401
rect 131854 59327 131910 59336
rect 131868 58682 131896 59327
rect 131856 58676 131908 58682
rect 131856 58618 131908 58624
rect 131764 33788 131816 33794
rect 131764 33730 131816 33736
rect 131120 25628 131172 25634
rect 131120 25570 131172 25576
rect 131132 16574 131160 25570
rect 131132 16546 131344 16574
rect 130384 4956 130436 4962
rect 130384 4898 130436 4904
rect 130304 3454 130608 3482
rect 130580 480 130608 3454
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 133156 8974 133184 59463
rect 133418 59392 133474 59401
rect 133418 59327 133474 59336
rect 133432 45554 133460 59327
rect 133340 45526 133460 45554
rect 133340 18630 133368 45526
rect 133880 22908 133932 22914
rect 133880 22850 133932 22856
rect 133328 18624 133380 18630
rect 133328 18566 133380 18572
rect 133144 8968 133196 8974
rect 133144 8910 133196 8916
rect 132960 4820 133012 4826
rect 132960 4762 133012 4768
rect 132972 480 133000 4762
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 133892 354 133920 22850
rect 134536 7614 134564 59706
rect 136638 59664 136694 59673
rect 136560 59622 136638 59650
rect 135996 59356 136048 59362
rect 135996 59298 136048 59304
rect 136008 45554 136036 59298
rect 136560 54534 136588 59622
rect 136638 59599 136694 59608
rect 138478 59664 138534 59673
rect 138478 59599 138534 59608
rect 139122 59664 139178 59673
rect 139122 59599 139178 59608
rect 137466 59528 137522 59537
rect 137466 59463 137522 59472
rect 137282 59256 137338 59265
rect 137282 59191 137338 59200
rect 136548 54528 136600 54534
rect 136548 54470 136600 54476
rect 136640 51876 136692 51882
rect 136640 51818 136692 51824
rect 135916 45526 136036 45554
rect 135260 18692 135312 18698
rect 135260 18634 135312 18640
rect 134524 7608 134576 7614
rect 134524 7550 134576 7556
rect 135272 480 135300 18634
rect 135916 3330 135944 45526
rect 136652 16574 136680 51818
rect 136652 16546 137232 16574
rect 136456 4956 136508 4962
rect 136456 4898 136508 4904
rect 135904 3324 135956 3330
rect 135904 3266 135956 3272
rect 136468 480 136496 4898
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 137296 3806 137324 59191
rect 137284 3800 137336 3806
rect 137284 3742 137336 3748
rect 137480 3262 137508 59463
rect 138492 59401 138520 59599
rect 137558 59392 137614 59401
rect 137558 59327 137560 59336
rect 137612 59327 137614 59336
rect 138478 59392 138534 59401
rect 138478 59327 138534 59336
rect 137560 59298 137612 59304
rect 138020 46300 138072 46306
rect 138020 46242 138072 46248
rect 138032 16574 138060 46242
rect 139136 45554 139164 59599
rect 139228 59537 139256 59735
rect 139214 59528 139270 59537
rect 139214 59463 139270 59472
rect 139964 59401 139992 59735
rect 141698 59735 141754 59744
rect 142434 59800 142490 59809
rect 142434 59735 142436 59744
rect 140228 59706 140280 59712
rect 140042 59528 140098 59537
rect 140042 59463 140098 59472
rect 139950 59392 140006 59401
rect 139950 59327 140006 59336
rect 138676 45526 139164 45554
rect 138032 16546 138612 16574
rect 138584 3482 138612 16546
rect 138676 3874 138704 45526
rect 140056 3942 140084 59463
rect 140044 3936 140096 3942
rect 140044 3878 140096 3884
rect 138664 3868 138716 3874
rect 138664 3810 138716 3816
rect 140044 3800 140096 3806
rect 140044 3742 140096 3748
rect 138584 3454 138888 3482
rect 137468 3256 137520 3262
rect 137468 3198 137520 3204
rect 138860 480 138888 3454
rect 140056 480 140084 3742
rect 140240 3534 140268 59706
rect 141606 59664 141662 59673
rect 141436 59622 141606 59650
rect 140780 29776 140832 29782
rect 140780 29718 140832 29724
rect 140792 16574 140820 29718
rect 140792 16546 141280 16574
rect 140228 3528 140280 3534
rect 140228 3470 140280 3476
rect 141252 480 141280 16546
rect 141436 3602 141464 59622
rect 141606 59599 141662 59608
rect 141712 59537 141740 59735
rect 142488 59735 142490 59744
rect 144274 59800 144330 59809
rect 149426 59800 149482 59809
rect 144274 59735 144330 59744
rect 148508 59764 148560 59770
rect 142436 59706 142488 59712
rect 144182 59664 144238 59673
rect 144182 59599 144238 59608
rect 141698 59528 141754 59537
rect 141698 59463 141754 59472
rect 141606 58984 141662 58993
rect 141606 58919 141662 58928
rect 141620 3670 141648 58919
rect 142804 58540 142856 58546
rect 142804 58482 142856 58488
rect 142160 32428 142212 32434
rect 142160 32370 142212 32376
rect 141608 3664 141660 3670
rect 141608 3606 141660 3612
rect 141424 3596 141476 3602
rect 141424 3538 141476 3544
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142172 354 142200 32370
rect 142816 3738 142844 58482
rect 143540 20120 143592 20126
rect 143540 20062 143592 20068
rect 142804 3732 142856 3738
rect 142804 3674 142856 3680
rect 143552 3534 143580 20062
rect 143540 3528 143592 3534
rect 143540 3470 143592 3476
rect 144196 3369 144224 59599
rect 144288 58546 144316 59735
rect 150806 59800 150862 59809
rect 149426 59735 149428 59744
rect 148508 59706 148560 59712
rect 149480 59735 149482 59744
rect 150268 59758 150806 59786
rect 149428 59706 149480 59712
rect 146666 59664 146722 59673
rect 146208 59628 146260 59634
rect 146666 59599 146722 59608
rect 147494 59664 147550 59673
rect 147494 59599 147496 59608
rect 146208 59570 146260 59576
rect 145562 59528 145618 59537
rect 145562 59463 145618 59472
rect 144366 59392 144422 59401
rect 144366 59327 144422 59336
rect 144276 58540 144328 58546
rect 144276 58482 144328 58488
rect 144380 3466 144408 59327
rect 145576 6186 145604 59463
rect 146220 58750 146248 59570
rect 146680 59401 146708 59599
rect 147548 59599 147550 59608
rect 147496 59570 147548 59576
rect 146944 59560 146996 59566
rect 146944 59502 146996 59508
rect 146666 59392 146722 59401
rect 146666 59327 146722 59336
rect 146208 58744 146260 58750
rect 146208 58686 146260 58692
rect 145564 6180 145616 6186
rect 145564 6122 145616 6128
rect 146956 4826 146984 59502
rect 148322 59392 148378 59401
rect 148322 59327 148378 59336
rect 147680 31272 147732 31278
rect 147680 31214 147732 31220
rect 147692 16574 147720 31214
rect 147692 16546 147904 16574
rect 146944 4820 146996 4826
rect 146944 4762 146996 4768
rect 144736 3528 144788 3534
rect 144736 3470 144788 3476
rect 144368 3460 144420 3466
rect 144368 3402 144420 3408
rect 144182 3360 144238 3369
rect 144182 3295 144238 3304
rect 143540 2984 143592 2990
rect 143540 2926 143592 2932
rect 143552 480 143580 2926
rect 144748 480 144776 3470
rect 145932 3460 145984 3466
rect 145932 3402 145984 3408
rect 145944 480 145972 3402
rect 147128 3120 147180 3126
rect 147128 3062 147180 3068
rect 147140 480 147168 3062
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 148336 3806 148364 59327
rect 148520 4962 148548 59706
rect 149150 59664 149206 59673
rect 149150 59599 149206 59608
rect 149702 59664 149758 59673
rect 149702 59599 149758 59608
rect 149164 59566 149192 59599
rect 149152 59560 149204 59566
rect 149152 59502 149204 59508
rect 148508 4956 148560 4962
rect 148508 4898 148560 4904
rect 148324 3800 148376 3806
rect 148324 3742 148376 3748
rect 149520 3528 149572 3534
rect 149520 3470 149572 3476
rect 149532 480 149560 3470
rect 149716 3126 149744 59599
rect 149886 59528 149942 59537
rect 149886 59463 149942 59472
rect 149704 3120 149756 3126
rect 149704 3062 149756 3068
rect 149900 2990 149928 59463
rect 150268 59401 150296 59758
rect 152462 59800 152518 59809
rect 150806 59735 150862 59744
rect 151728 59764 151780 59770
rect 156602 59800 156658 59809
rect 152462 59735 152464 59744
rect 151728 59706 151780 59712
rect 152516 59735 152518 59744
rect 154304 59764 154356 59770
rect 152464 59706 152516 59712
rect 159914 59800 159970 59809
rect 156602 59735 156604 59744
rect 154304 59706 154356 59712
rect 156656 59735 156658 59744
rect 158536 59764 158588 59770
rect 156604 59706 156656 59712
rect 159914 59735 159970 59744
rect 160742 59800 160798 59809
rect 167458 59800 167514 59809
rect 160742 59735 160744 59744
rect 158536 59706 158588 59712
rect 151740 59673 151768 59706
rect 151726 59664 151782 59673
rect 151726 59599 151782 59608
rect 153106 59528 153162 59537
rect 153106 59463 153162 59472
rect 150254 59392 150310 59401
rect 150254 59327 150310 59336
rect 150438 59392 150494 59401
rect 150438 59327 150494 59336
rect 153014 59392 153070 59401
rect 153014 59327 153070 59336
rect 150452 16574 150480 59327
rect 151820 21548 151872 21554
rect 151820 21490 151872 21496
rect 150452 16546 150664 16574
rect 149888 2984 149940 2990
rect 149888 2926 149940 2932
rect 150636 480 150664 16546
rect 151832 480 151860 21490
rect 153028 12238 153056 59327
rect 153016 12232 153068 12238
rect 153016 12174 153068 12180
rect 153120 4214 153148 59463
rect 154316 4826 154344 59706
rect 158352 59696 158404 59702
rect 156602 59664 156658 59673
rect 158352 59638 158404 59644
rect 156602 59599 156658 59608
rect 156616 59401 156644 59599
rect 156970 59528 157026 59537
rect 157246 59528 157302 59537
rect 156970 59463 157026 59472
rect 157064 59492 157116 59498
rect 155866 59392 155922 59401
rect 155866 59327 155922 59336
rect 156602 59392 156658 59401
rect 156984 59362 157012 59463
rect 157246 59463 157302 59472
rect 157340 59492 157392 59498
rect 157064 59434 157116 59440
rect 156602 59327 156658 59336
rect 156972 59356 157024 59362
rect 155408 13388 155460 13394
rect 155408 13330 155460 13336
rect 154304 4820 154356 4826
rect 154304 4762 154356 4768
rect 153108 4208 153160 4214
rect 153108 4150 153160 4156
rect 154212 4208 154264 4214
rect 154212 4150 154264 4156
rect 153016 3392 153068 3398
rect 153016 3334 153068 3340
rect 153028 480 153056 3334
rect 154224 480 154252 4150
rect 155420 480 155448 13330
rect 155880 6186 155908 59327
rect 156972 59298 157024 59304
rect 157076 9042 157104 59434
rect 157064 9036 157116 9042
rect 157064 8978 157116 8984
rect 157260 7682 157288 59463
rect 157340 59434 157392 59440
rect 157352 59401 157380 59434
rect 157338 59392 157394 59401
rect 157338 59327 157394 59336
rect 157800 12232 157852 12238
rect 157800 12174 157852 12180
rect 157248 7676 157300 7682
rect 157248 7618 157300 7624
rect 155868 6180 155920 6186
rect 155868 6122 155920 6128
rect 156604 3664 156656 3670
rect 156604 3606 156656 3612
rect 156616 480 156644 3606
rect 157812 480 157840 12174
rect 158364 11762 158392 59638
rect 158548 44878 158576 59706
rect 159928 59702 159956 59735
rect 160796 59735 160798 59744
rect 165252 59764 165304 59770
rect 160744 59706 160796 59712
rect 174542 59800 174598 59809
rect 167458 59735 167460 59744
rect 165252 59706 165304 59712
rect 167512 59735 167514 59744
rect 173624 59764 173676 59770
rect 167460 59706 167512 59712
rect 174542 59735 174598 59744
rect 175738 59800 175794 59809
rect 182362 59800 182418 59809
rect 175738 59735 175740 59744
rect 173624 59706 173676 59712
rect 159916 59696 159968 59702
rect 162858 59664 162914 59673
rect 159916 59638 159968 59644
rect 162780 59622 162858 59650
rect 160006 59528 160062 59537
rect 160006 59463 160062 59472
rect 161110 59528 161166 59537
rect 161110 59463 161166 59472
rect 158536 44872 158588 44878
rect 158536 44814 158588 44820
rect 158720 40928 158772 40934
rect 158720 40870 158772 40876
rect 158732 16574 158760 40870
rect 158732 16546 158944 16574
rect 158352 11756 158404 11762
rect 158352 11698 158404 11704
rect 158916 480 158944 16546
rect 160020 7614 160048 59463
rect 160100 59356 160152 59362
rect 160100 59298 160152 59304
rect 160008 7608 160060 7614
rect 160008 7550 160060 7556
rect 160112 3602 160140 59298
rect 161124 8974 161152 59463
rect 161294 59392 161350 59401
rect 161294 59327 161350 59336
rect 161308 14482 161336 59327
rect 162780 16046 162808 59622
rect 162858 59599 162914 59608
rect 163870 59528 163926 59537
rect 163870 59463 163926 59472
rect 162860 57316 162912 57322
rect 162860 57258 162912 57264
rect 162872 16574 162900 57258
rect 163884 17270 163912 59463
rect 164054 59392 164110 59401
rect 164054 59327 164110 59336
rect 164068 18630 164096 59327
rect 164056 18624 164108 18630
rect 164056 18566 164108 18572
rect 163872 17264 163924 17270
rect 163872 17206 163924 17212
rect 162872 16546 163728 16574
rect 162768 16040 162820 16046
rect 162768 15982 162820 15988
rect 161296 14476 161348 14482
rect 161296 14418 161348 14424
rect 162032 10464 162084 10470
rect 162032 10406 162084 10412
rect 161112 8968 161164 8974
rect 161112 8910 161164 8916
rect 160192 3732 160244 3738
rect 160192 3674 160244 3680
rect 160100 3596 160152 3602
rect 160100 3538 160152 3544
rect 160204 1850 160232 3674
rect 161296 3596 161348 3602
rect 161296 3538 161348 3544
rect 161388 3596 161440 3602
rect 161388 3538 161440 3544
rect 160112 1822 160232 1850
rect 160112 480 160140 1822
rect 161308 480 161336 3538
rect 161400 3398 161428 3538
rect 161388 3392 161440 3398
rect 161388 3334 161440 3340
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 10406
rect 163700 480 163728 16546
rect 165264 5098 165292 59706
rect 168286 59528 168342 59537
rect 169942 59528 169998 59537
rect 168286 59463 168342 59472
rect 169404 59486 169942 59514
rect 166906 59392 166962 59401
rect 166906 59327 166962 59336
rect 168102 59392 168158 59401
rect 168102 59327 168158 59336
rect 165434 59256 165490 59265
rect 165434 59191 165490 59200
rect 165448 5302 165476 59191
rect 165620 57384 165672 57390
rect 165620 57326 165672 57332
rect 165632 16574 165660 57326
rect 165632 16546 166120 16574
rect 165436 5296 165488 5302
rect 165436 5238 165488 5244
rect 165252 5092 165304 5098
rect 165252 5034 165304 5040
rect 164884 4820 164936 4826
rect 164884 4762 164936 4768
rect 164896 480 164924 4762
rect 166092 480 166120 16546
rect 166920 5030 166948 59327
rect 168116 21418 168144 59327
rect 168104 21412 168156 21418
rect 168104 21354 168156 21360
rect 168300 19990 168328 59463
rect 169404 59401 169432 59486
rect 169942 59463 169998 59472
rect 171598 59528 171654 59537
rect 171598 59463 171654 59472
rect 171612 59430 171640 59463
rect 169484 59424 169536 59430
rect 169390 59392 169446 59401
rect 171600 59424 171652 59430
rect 169484 59366 169536 59372
rect 169574 59392 169630 59401
rect 169390 59327 169446 59336
rect 168380 56024 168432 56030
rect 168380 55966 168432 55972
rect 168288 19984 168340 19990
rect 168288 19926 168340 19932
rect 168392 7682 168420 55966
rect 169496 45554 169524 59366
rect 171600 59366 171652 59372
rect 169574 59327 169630 59336
rect 169404 45526 169524 45554
rect 168380 7676 168432 7682
rect 168380 7618 168432 7624
rect 168380 6180 168432 6186
rect 168380 6122 168432 6128
rect 166908 5024 166960 5030
rect 166908 4966 166960 4972
rect 167184 4140 167236 4146
rect 167184 4082 167236 4088
rect 167196 480 167224 4082
rect 168392 480 168420 6122
rect 169404 4894 169432 45526
rect 169588 12434 169616 59327
rect 171046 59256 171102 59265
rect 171046 59191 171102 59200
rect 172426 59256 172482 59265
rect 172426 59191 172482 59200
rect 170404 53236 170456 53242
rect 170404 53178 170456 53184
rect 169760 50516 169812 50522
rect 169760 50458 169812 50464
rect 169772 16574 169800 50458
rect 169772 16546 170352 16574
rect 169588 12406 169708 12434
rect 169576 7676 169628 7682
rect 169576 7618 169628 7624
rect 169392 4888 169444 4894
rect 169392 4830 169444 4836
rect 169588 480 169616 7618
rect 169680 4962 169708 12406
rect 169668 4956 169720 4962
rect 169668 4898 169720 4904
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 16546
rect 170416 4146 170444 53178
rect 171060 4826 171088 59191
rect 172440 25770 172468 59191
rect 172520 49224 172572 49230
rect 172520 49166 172572 49172
rect 172428 25764 172480 25770
rect 172428 25706 172480 25712
rect 172532 16574 172560 49166
rect 173636 28286 173664 59706
rect 173806 59528 173862 59537
rect 173806 59463 173862 59472
rect 173624 28280 173676 28286
rect 173624 28222 173676 28228
rect 173820 26926 173848 59463
rect 174556 58886 174584 59735
rect 175792 59735 175794 59744
rect 180616 59764 180668 59770
rect 175740 59706 175792 59712
rect 182362 59735 182364 59744
rect 180616 59706 180668 59712
rect 182416 59735 182418 59744
rect 183190 59800 183246 59809
rect 185674 59800 185730 59809
rect 183190 59735 183246 59744
rect 184572 59764 184624 59770
rect 182364 59706 182416 59712
rect 179328 59628 179380 59634
rect 179328 59570 179380 59576
rect 176474 59528 176530 59537
rect 176292 59492 176344 59498
rect 176474 59463 176530 59472
rect 178222 59528 178278 59537
rect 178222 59463 178224 59472
rect 176292 59434 176344 59440
rect 175186 59392 175242 59401
rect 175186 59327 175242 59336
rect 174544 58880 174596 58886
rect 174544 58822 174596 58828
rect 175200 31074 175228 59327
rect 175188 31068 175240 31074
rect 175188 31010 175240 31016
rect 173808 26920 173860 26926
rect 173808 26862 173860 26868
rect 172532 16546 172744 16574
rect 171968 7744 172020 7750
rect 171968 7686 172020 7692
rect 171048 4820 171100 4826
rect 171048 4762 171100 4768
rect 170404 4140 170456 4146
rect 170404 4082 170456 4088
rect 171980 480 172008 7686
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 173900 13116 173952 13122
rect 173900 13058 173952 13064
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173912 354 173940 13058
rect 175464 9036 175516 9042
rect 175464 8978 175516 8984
rect 175476 480 175504 8978
rect 176304 6594 176332 59434
rect 176488 6662 176516 59463
rect 178276 59463 178278 59472
rect 178224 59434 178276 59440
rect 177670 59392 177726 59401
rect 177670 59327 177726 59336
rect 176660 47796 176712 47802
rect 176660 47738 176712 47744
rect 176476 6656 176528 6662
rect 176476 6598 176528 6604
rect 176292 6588 176344 6594
rect 176292 6530 176344 6536
rect 176672 480 176700 47738
rect 177684 32638 177712 59327
rect 177854 59256 177910 59265
rect 177854 59191 177910 59200
rect 177868 43654 177896 59191
rect 177856 43648 177908 43654
rect 177856 43590 177908 43596
rect 177672 32632 177724 32638
rect 177672 32574 177724 32580
rect 177856 13184 177908 13190
rect 177856 13126 177908 13132
rect 177868 480 177896 13126
rect 178592 11756 178644 11762
rect 178592 11698 178644 11704
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 173134 -960 173246 326
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 11698
rect 179340 6526 179368 59570
rect 180248 15904 180300 15910
rect 180248 15846 180300 15852
rect 179328 6520 179380 6526
rect 179328 6462 179380 6468
rect 180260 480 180288 15846
rect 180628 6390 180656 59706
rect 180706 59664 180762 59673
rect 182362 59664 182418 59673
rect 180706 59599 180708 59608
rect 180760 59599 180762 59608
rect 182008 59622 182362 59650
rect 180708 59570 180760 59576
rect 180706 59528 180762 59537
rect 180706 59463 180762 59472
rect 180720 6458 180748 59463
rect 181810 59392 181866 59401
rect 181810 59327 181866 59336
rect 180984 13252 181036 13258
rect 180984 13194 181036 13200
rect 180708 6452 180760 6458
rect 180708 6394 180760 6400
rect 180616 6384 180668 6390
rect 180616 6326 180668 6332
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 13194
rect 181824 6322 181852 59327
rect 181812 6316 181864 6322
rect 181812 6258 181864 6264
rect 182008 6254 182036 59622
rect 182362 59599 182418 59608
rect 183204 59401 183232 59735
rect 185674 59735 185676 59744
rect 184572 59706 184624 59712
rect 185728 59735 185730 59744
rect 187422 59800 187478 59809
rect 189906 59800 189962 59809
rect 187422 59735 187478 59744
rect 188712 59764 188764 59770
rect 185676 59706 185728 59712
rect 183190 59392 183246 59401
rect 183190 59327 183246 59336
rect 183466 59256 183522 59265
rect 183466 59191 183522 59200
rect 182180 44872 182232 44878
rect 182180 44814 182232 44820
rect 181996 6248 182048 6254
rect 181996 6190 182048 6196
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 44814
rect 183480 6186 183508 59191
rect 183560 50584 183612 50590
rect 183560 50526 183612 50532
rect 183572 16574 183600 50526
rect 183572 16546 183784 16574
rect 183468 6180 183520 6186
rect 183468 6122 183520 6128
rect 183756 480 183784 16546
rect 184584 15978 184612 59706
rect 187330 59664 187386 59673
rect 187330 59599 187386 59608
rect 186134 59528 186190 59537
rect 186134 59463 186190 59472
rect 185950 59392 186006 59401
rect 185950 59327 186006 59336
rect 184754 59256 184810 59265
rect 184754 59191 184810 59200
rect 184768 33998 184796 59191
rect 185964 35290 185992 59327
rect 186148 42158 186176 59463
rect 187344 59401 187372 59599
rect 187436 59537 187464 59735
rect 189906 59735 189908 59744
rect 188712 59706 188764 59712
rect 189960 59735 189962 59744
rect 196530 59800 196586 59809
rect 196530 59735 196586 59744
rect 201498 59800 201554 59809
rect 204810 59800 204866 59809
rect 201498 59735 201554 59744
rect 202696 59764 202748 59770
rect 189908 59706 189960 59712
rect 187422 59528 187478 59537
rect 187422 59463 187478 59472
rect 187330 59392 187386 59401
rect 187330 59327 187386 59336
rect 187606 59392 187662 59401
rect 187606 59327 187662 59336
rect 186320 58812 186372 58818
rect 186320 58754 186372 58760
rect 186136 42152 186188 42158
rect 186136 42094 186188 42100
rect 185952 35284 186004 35290
rect 185952 35226 186004 35232
rect 184756 33992 184808 33998
rect 184756 33934 184808 33940
rect 186332 16574 186360 58754
rect 186964 49156 187016 49162
rect 186964 49098 187016 49104
rect 186332 16546 186912 16574
rect 184572 15972 184624 15978
rect 184572 15914 184624 15920
rect 186136 7608 186188 7614
rect 186136 7550 186188 7556
rect 184940 2984 184992 2990
rect 184940 2926 184992 2932
rect 184952 480 184980 2926
rect 186148 480 186176 7550
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 186976 2990 187004 49098
rect 187620 36650 187648 59327
rect 188724 38010 188752 59706
rect 191746 59664 191802 59673
rect 191576 59622 191746 59650
rect 190090 59528 190146 59537
rect 190090 59463 190146 59472
rect 188894 59256 188950 59265
rect 188894 59191 188950 59200
rect 188908 39506 188936 59191
rect 190104 40798 190132 59463
rect 191576 59401 191604 59622
rect 191746 59599 191802 59608
rect 193034 59528 193090 59537
rect 194874 59528 194930 59537
rect 193034 59463 193090 59472
rect 194336 59486 194874 59514
rect 190274 59392 190330 59401
rect 190274 59327 190330 59336
rect 191562 59392 191618 59401
rect 191562 59327 191618 59336
rect 191746 59392 191802 59401
rect 191746 59327 191802 59336
rect 192850 59392 192906 59401
rect 192850 59327 192906 59336
rect 190288 51814 190316 59327
rect 190460 54732 190512 54738
rect 190460 54674 190512 54680
rect 190276 51808 190328 51814
rect 190276 51750 190328 51756
rect 190092 40792 190144 40798
rect 190092 40734 190144 40740
rect 188896 39500 188948 39506
rect 188896 39442 188948 39448
rect 188712 38004 188764 38010
rect 188712 37946 188764 37952
rect 187608 36644 187660 36650
rect 187608 36586 187660 36592
rect 188528 13320 188580 13326
rect 188528 13262 188580 13268
rect 186964 2984 187016 2990
rect 186964 2926 187016 2932
rect 188540 480 188568 13262
rect 189724 8968 189776 8974
rect 189724 8910 189776 8916
rect 189736 480 189764 8910
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190472 354 190500 54674
rect 191760 29714 191788 59327
rect 191748 29708 191800 29714
rect 191748 29650 191800 29656
rect 191840 27056 191892 27062
rect 191840 26998 191892 27004
rect 191852 16574 191880 26998
rect 192864 22846 192892 59327
rect 193048 32570 193076 59463
rect 194336 59401 194364 59486
rect 194874 59463 194930 59472
rect 196544 59430 196572 59735
rect 200670 59664 200726 59673
rect 198556 59628 198608 59634
rect 200670 59599 200672 59608
rect 198556 59570 198608 59576
rect 200724 59599 200726 59608
rect 200672 59570 200724 59576
rect 197174 59528 197230 59537
rect 197174 59463 197230 59472
rect 194416 59424 194468 59430
rect 194322 59392 194378 59401
rect 196532 59424 196584 59430
rect 194416 59366 194468 59372
rect 194506 59392 194562 59401
rect 194322 59327 194378 59336
rect 193220 46436 193272 46442
rect 193220 46378 193272 46384
rect 193036 32564 193088 32570
rect 193036 32506 193088 32512
rect 192852 22840 192904 22846
rect 192852 22782 192904 22788
rect 191852 16546 192064 16574
rect 192036 480 192064 16546
rect 193232 3806 193260 46378
rect 194428 45554 194456 59366
rect 196532 59366 196584 59372
rect 196990 59392 197046 59401
rect 194506 59327 194562 59336
rect 196990 59327 197046 59336
rect 194336 45526 194456 45554
rect 194336 44946 194364 45526
rect 194324 44940 194376 44946
rect 194324 44882 194376 44888
rect 194520 43586 194548 59327
rect 195886 59256 195942 59265
rect 195886 59191 195942 59200
rect 194600 58744 194652 58750
rect 194600 58686 194652 58692
rect 194508 43580 194560 43586
rect 194508 43522 194560 43528
rect 194612 16574 194640 58686
rect 195900 24206 195928 59191
rect 195888 24200 195940 24206
rect 195888 24142 195940 24148
rect 194612 16546 195192 16574
rect 193312 14476 193364 14482
rect 193312 14418 193364 14424
rect 193220 3800 193272 3806
rect 193220 3742 193272 3748
rect 193324 3482 193352 14418
rect 194416 3800 194468 3806
rect 194416 3742 194468 3748
rect 193232 3454 193352 3482
rect 193232 480 193260 3454
rect 194428 480 194456 3742
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 196808 16040 196860 16046
rect 196808 15982 196860 15988
rect 196820 480 196848 15982
rect 197004 7750 197032 59327
rect 197188 33862 197216 59463
rect 198370 59256 198426 59265
rect 198370 59191 198426 59200
rect 197176 33856 197228 33862
rect 197176 33798 197228 33804
rect 197912 11756 197964 11762
rect 197912 11698 197964 11704
rect 196992 7744 197044 7750
rect 196992 7686 197044 7692
rect 197924 480 197952 11698
rect 198384 7682 198412 59191
rect 198372 7676 198424 7682
rect 198372 7618 198424 7624
rect 198568 7614 198596 59570
rect 201130 59528 201186 59537
rect 201130 59463 201186 59472
rect 200026 59256 200082 59265
rect 200026 59191 200082 59200
rect 198740 54664 198792 54670
rect 198740 54606 198792 54612
rect 198556 7608 198608 7614
rect 198556 7550 198608 7556
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 54606
rect 200040 17474 200068 59191
rect 201144 35358 201172 59463
rect 201512 59401 201540 59735
rect 213182 59800 213238 59809
rect 204810 59735 204812 59744
rect 202696 59706 202748 59712
rect 204864 59735 204866 59744
rect 209412 59764 209464 59770
rect 204812 59706 204864 59712
rect 209412 59706 209464 59712
rect 209872 59764 209924 59770
rect 209872 59706 209924 59712
rect 210792 59764 210844 59770
rect 213182 59735 213184 59744
rect 210792 59706 210844 59712
rect 213236 59735 213238 59744
rect 214010 59800 214066 59809
rect 218150 59800 218206 59809
rect 214010 59735 214066 59744
rect 216588 59764 216640 59770
rect 213184 59706 213236 59712
rect 202510 59528 202566 59537
rect 202510 59463 202566 59472
rect 201498 59392 201554 59401
rect 201498 59327 201554 59336
rect 201314 59256 201370 59265
rect 201314 59191 201370 59200
rect 201328 42226 201356 59191
rect 201500 45008 201552 45014
rect 201500 44950 201552 44956
rect 201316 42220 201368 42226
rect 201316 42162 201368 42168
rect 201132 35352 201184 35358
rect 201132 35294 201184 35300
rect 200028 17468 200080 17474
rect 200028 17410 200080 17416
rect 200120 17264 200172 17270
rect 200120 17206 200172 17212
rect 200132 16574 200160 17206
rect 200132 16546 200344 16574
rect 200316 480 200344 16546
rect 201512 480 201540 44950
rect 202524 36718 202552 59463
rect 202708 38078 202736 59706
rect 203154 59664 203210 59673
rect 203154 59599 203210 59608
rect 203168 59401 203196 59599
rect 205454 59528 205510 59537
rect 205272 59492 205324 59498
rect 205454 59463 205510 59472
rect 207294 59528 207350 59537
rect 207294 59463 207296 59472
rect 205272 59434 205324 59440
rect 203154 59392 203210 59401
rect 203154 59327 203210 59336
rect 204166 59392 204222 59401
rect 204166 59327 204222 59336
rect 204180 39438 204208 59327
rect 204168 39432 204220 39438
rect 204168 39374 204220 39380
rect 202696 38072 202748 38078
rect 202696 38014 202748 38020
rect 202512 36712 202564 36718
rect 202512 36654 202564 36660
rect 201592 31204 201644 31210
rect 201592 31146 201644 31152
rect 201604 16574 201632 31146
rect 205284 18766 205312 59434
rect 205468 40730 205496 59463
rect 207348 59463 207350 59472
rect 207296 59434 207348 59440
rect 206650 59392 206706 59401
rect 206650 59327 206706 59336
rect 205640 43512 205692 43518
rect 205640 43454 205692 43460
rect 205456 40724 205508 40730
rect 205456 40666 205508 40672
rect 205272 18760 205324 18766
rect 205272 18702 205324 18708
rect 202880 18624 202932 18630
rect 202880 18566 202932 18572
rect 202892 16574 202920 18566
rect 205652 16574 205680 43454
rect 206664 20058 206692 59327
rect 206834 59256 206890 59265
rect 206834 59191 206890 59200
rect 206848 46374 206876 59191
rect 208306 59120 208362 59129
rect 208306 59055 208362 59064
rect 206836 46368 206888 46374
rect 206836 46310 206888 46316
rect 208320 21486 208348 59055
rect 208308 21480 208360 21486
rect 208308 21422 208360 21428
rect 206652 20052 206704 20058
rect 206652 19994 206704 20000
rect 201604 16546 202736 16574
rect 202892 16546 203472 16574
rect 205652 16546 206232 16574
rect 202708 480 202736 16546
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 16546
rect 205088 11824 205140 11830
rect 205088 11766 205140 11772
rect 205100 480 205128 11766
rect 206204 480 206232 16546
rect 208584 11892 208636 11898
rect 208584 11834 208636 11840
rect 207388 5160 207440 5166
rect 207388 5102 207440 5108
rect 207400 480 207428 5102
rect 208596 480 208624 11834
rect 209424 9178 209452 59706
rect 209884 59537 209912 59706
rect 210698 59664 210754 59673
rect 210698 59599 210754 59608
rect 209870 59528 209926 59537
rect 209870 59463 209926 59472
rect 210712 59401 210740 59599
rect 209594 59392 209650 59401
rect 209594 59327 209650 59336
rect 210698 59392 210754 59401
rect 210698 59327 210754 59336
rect 209608 9246 209636 59327
rect 209780 17400 209832 17406
rect 209780 17342 209832 17348
rect 209596 9240 209648 9246
rect 209596 9182 209648 9188
rect 209412 9172 209464 9178
rect 209412 9114 209464 9120
rect 209792 480 209820 17342
rect 210804 9110 210832 59706
rect 213550 59664 213606 59673
rect 213550 59599 213606 59608
rect 210974 59392 211030 59401
rect 210974 59327 211030 59336
rect 210988 25702 211016 59327
rect 212446 59256 212502 59265
rect 212446 59191 212502 59200
rect 212460 26994 212488 59191
rect 212448 26988 212500 26994
rect 212448 26930 212500 26936
rect 210976 25696 211028 25702
rect 210976 25638 211028 25644
rect 211712 11960 211764 11966
rect 211712 11902 211764 11908
rect 210792 9104 210844 9110
rect 210792 9046 210844 9052
rect 210976 5092 211028 5098
rect 210976 5034 211028 5040
rect 210988 480 211016 5034
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 11902
rect 213564 9042 213592 59599
rect 214024 59401 214052 59735
rect 221462 59800 221518 59809
rect 218150 59735 218152 59744
rect 216588 59706 216640 59712
rect 218204 59735 218206 59744
rect 219256 59764 219308 59770
rect 218152 59706 218204 59712
rect 225234 59800 225290 59809
rect 221462 59735 221464 59744
rect 219256 59706 219308 59712
rect 221516 59735 221518 59744
rect 224604 59758 225234 59786
rect 221464 59706 221516 59712
rect 215758 59664 215814 59673
rect 215758 59599 215814 59608
rect 214930 59528 214986 59537
rect 214930 59463 214986 59472
rect 215116 59492 215168 59498
rect 214010 59392 214066 59401
rect 214010 59327 214066 59336
rect 213734 59256 213790 59265
rect 213734 59191 213790 59200
rect 213552 9036 213604 9042
rect 213552 8978 213604 8984
rect 213748 8974 213776 59191
rect 214564 47728 214616 47734
rect 214564 47670 214616 47676
rect 213736 8968 213788 8974
rect 213736 8910 213788 8916
rect 214472 5024 214524 5030
rect 214472 4966 214524 4972
rect 213368 3392 213420 3398
rect 213368 3334 213420 3340
rect 213380 480 213408 3334
rect 214484 480 214512 4966
rect 214576 3398 214604 47670
rect 214944 32502 214972 59463
rect 215116 59434 215168 59440
rect 215128 47666 215156 59434
rect 215772 59401 215800 59599
rect 215944 59492 215996 59498
rect 215944 59434 215996 59440
rect 215956 59401 215984 59434
rect 215758 59392 215814 59401
rect 215758 59327 215814 59336
rect 215942 59392 215998 59401
rect 215942 59327 215998 59336
rect 215116 47660 215168 47666
rect 215116 47602 215168 47608
rect 214932 32496 214984 32502
rect 214932 32438 214984 32444
rect 216600 28422 216628 59706
rect 219070 59528 219126 59537
rect 219070 59463 219126 59472
rect 217874 59256 217930 59265
rect 217874 59191 217930 59200
rect 217690 59120 217746 59129
rect 217690 59055 217746 59064
rect 216680 33924 216732 33930
rect 216680 33866 216732 33872
rect 216588 28416 216640 28422
rect 216588 28358 216640 28364
rect 216692 16574 216720 33866
rect 217704 31142 217732 59055
rect 217888 43450 217916 59191
rect 218060 56092 218112 56098
rect 218060 56034 218112 56040
rect 217876 43444 217928 43450
rect 217876 43386 217928 43392
rect 217692 31136 217744 31142
rect 217692 31078 217744 31084
rect 216692 16546 216904 16574
rect 215300 12028 215352 12034
rect 215300 11970 215352 11976
rect 214564 3392 214616 3398
rect 214564 3334 214616 3340
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 11970
rect 216876 480 216904 16546
rect 218072 11694 218100 56034
rect 219084 33794 219112 59463
rect 219268 49094 219296 59706
rect 219806 59664 219862 59673
rect 219806 59599 219862 59608
rect 219820 59401 219848 59599
rect 222106 59528 222162 59537
rect 222106 59463 222162 59472
rect 219806 59392 219862 59401
rect 219806 59327 219862 59336
rect 220726 59392 220782 59401
rect 220726 59327 220782 59336
rect 222014 59392 222070 59401
rect 222014 59327 222070 59336
rect 219256 49088 219308 49094
rect 219256 49030 219308 49036
rect 220740 35222 220768 59327
rect 222028 53174 222056 59327
rect 222016 53168 222068 53174
rect 222016 53110 222068 53116
rect 222120 50454 222148 59463
rect 223486 59256 223542 59265
rect 223486 59191 223542 59200
rect 222200 57520 222252 57526
rect 222200 57462 222252 57468
rect 222108 50448 222160 50454
rect 222108 50390 222160 50396
rect 220728 35216 220780 35222
rect 220728 35158 220780 35164
rect 219072 33788 219124 33794
rect 219072 33730 219124 33736
rect 220820 21412 220872 21418
rect 220820 21354 220872 21360
rect 218152 19984 218204 19990
rect 218152 19926 218204 19932
rect 218060 11688 218112 11694
rect 218060 11630 218112 11636
rect 218164 6914 218192 19926
rect 220832 16574 220860 21354
rect 222212 16574 222240 57462
rect 223500 36582 223528 59191
rect 223488 36576 223540 36582
rect 223488 36518 223540 36524
rect 220832 16546 221136 16574
rect 222212 16546 222792 16574
rect 219992 14476 220044 14482
rect 219992 14418 220044 14424
rect 219256 11688 219308 11694
rect 219256 11630 219308 11636
rect 218072 6886 218192 6914
rect 218072 480 218100 6886
rect 219268 480 219296 11630
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 14418
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 16546
rect 222764 480 222792 16546
rect 223580 14544 223632 14550
rect 223580 14486 223632 14492
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 14486
rect 224604 10402 224632 59758
rect 225234 59735 225290 59744
rect 232778 59800 232834 59809
rect 232778 59735 232834 59744
rect 235262 59800 235318 59809
rect 235262 59735 235318 59744
rect 235446 59800 235502 59809
rect 235446 59735 235502 59744
rect 236918 59800 236974 59809
rect 239954 59800 240010 59809
rect 236918 59735 236974 59744
rect 238576 59764 238628 59770
rect 224958 59664 225014 59673
rect 228914 59664 228970 59673
rect 224958 59599 225014 59608
rect 227628 59628 227680 59634
rect 224774 59528 224830 59537
rect 224774 59463 224830 59472
rect 224788 42090 224816 59463
rect 224972 59401 225000 59599
rect 228914 59599 228916 59608
rect 227628 59570 227680 59576
rect 228968 59599 228970 59608
rect 228916 59570 228968 59576
rect 226154 59528 226210 59537
rect 226154 59463 226210 59472
rect 224958 59392 225014 59401
rect 224958 59327 225014 59336
rect 225970 59392 226026 59401
rect 225970 59327 226026 59336
rect 224776 42084 224828 42090
rect 224776 42026 224828 42032
rect 225984 37942 226012 59327
rect 226168 54602 226196 59463
rect 226156 54596 226208 54602
rect 226156 54538 226208 54544
rect 227640 39370 227668 59570
rect 229006 59528 229062 59537
rect 229006 59463 229062 59472
rect 231766 59528 231822 59537
rect 231766 59463 231822 59472
rect 228914 59392 228970 59401
rect 228914 59327 228970 59336
rect 228928 45554 228956 59327
rect 228836 45526 228956 45554
rect 227628 39364 227680 39370
rect 227628 39306 227680 39312
rect 225972 37936 226024 37942
rect 225972 37878 226024 37884
rect 228836 17270 228864 45526
rect 228824 17264 228876 17270
rect 228824 17206 228876 17212
rect 227536 14612 227588 14618
rect 227536 14554 227588 14560
rect 226340 12096 226392 12102
rect 226340 12038 226392 12044
rect 224592 10396 224644 10402
rect 224592 10338 224644 10344
rect 225144 4956 225196 4962
rect 225144 4898 225196 4904
rect 225156 480 225184 4898
rect 226352 480 226380 12038
rect 227548 480 227576 14554
rect 229020 10334 229048 59463
rect 230202 59256 230258 59265
rect 230202 59191 230258 59200
rect 229100 29844 229152 29850
rect 229100 29786 229152 29792
rect 229112 16574 229140 29786
rect 230216 18630 230244 59191
rect 231780 19990 231808 59463
rect 232792 58682 232820 59735
rect 234250 59664 234306 59673
rect 234250 59599 234306 59608
rect 232962 59392 233018 59401
rect 232962 59327 233018 59336
rect 232780 58676 232832 58682
rect 232780 58618 232832 58624
rect 232976 21418 233004 59327
rect 234264 22778 234292 59599
rect 234620 58880 234672 58886
rect 234620 58822 234672 58828
rect 234252 22772 234304 22778
rect 234252 22714 234304 22720
rect 232964 21412 233016 21418
rect 232964 21354 233016 21360
rect 231768 19984 231820 19990
rect 231768 19926 231820 19932
rect 230204 18624 230256 18630
rect 230204 18566 230256 18572
rect 229112 16546 229416 16574
rect 229008 10328 229060 10334
rect 229008 10270 229060 10276
rect 228732 4888 228784 4894
rect 228732 4830 228784 4836
rect 228744 480 228772 4830
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229388 354 229416 16546
rect 233424 16040 233476 16046
rect 233424 15982 233476 15988
rect 231032 14680 231084 14686
rect 231032 14622 231084 14628
rect 231044 480 231072 14622
rect 232228 4820 232280 4826
rect 232228 4762 232280 4768
rect 232240 480 232268 4762
rect 233436 480 233464 15982
rect 234632 11694 234660 58822
rect 235276 57254 235304 59735
rect 235460 59401 235488 59735
rect 235906 59528 235962 59537
rect 235906 59463 235962 59472
rect 235446 59392 235502 59401
rect 235446 59327 235502 59336
rect 235264 57248 235316 57254
rect 235264 57190 235316 57196
rect 235920 24138 235948 59463
rect 236000 58880 236052 58886
rect 236000 58822 236052 58828
rect 235908 24132 235960 24138
rect 235908 24074 235960 24080
rect 236012 16574 236040 58822
rect 236932 55894 236960 59735
rect 239954 59735 240010 59744
rect 240598 59800 240654 59809
rect 244738 59800 244794 59809
rect 240598 59735 240600 59744
rect 238576 59706 238628 59712
rect 238390 59664 238446 59673
rect 238390 59599 238446 59608
rect 237286 59392 237342 59401
rect 237286 59327 237342 59336
rect 236920 55888 236972 55894
rect 236920 55830 236972 55836
rect 237300 54534 237328 59327
rect 237288 54528 237340 54534
rect 237288 54470 237340 54476
rect 236012 16546 236592 16574
rect 234712 14748 234764 14754
rect 234712 14690 234764 14696
rect 234620 11688 234672 11694
rect 234620 11630 234672 11636
rect 234724 6914 234752 14690
rect 235816 11688 235868 11694
rect 235816 11630 235868 11636
rect 234632 6886 234752 6914
rect 234632 480 234660 6886
rect 235828 480 235856 11630
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 237656 14816 237708 14822
rect 237656 14758 237708 14764
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 14758
rect 238404 5166 238432 59599
rect 238588 25566 238616 59706
rect 239968 53106 239996 59735
rect 240652 59735 240654 59744
rect 242716 59764 242768 59770
rect 240600 59706 240652 59712
rect 249706 59800 249762 59809
rect 244738 59735 244740 59744
rect 242716 59706 242768 59712
rect 244792 59735 244794 59744
rect 248328 59764 248380 59770
rect 244740 59706 244792 59712
rect 249706 59735 249708 59744
rect 248328 59706 248380 59712
rect 249760 59735 249762 59744
rect 250534 59800 250590 59809
rect 253202 59800 253258 59809
rect 250534 59735 250590 59744
rect 251824 59764 251876 59770
rect 249708 59706 249760 59712
rect 241334 59528 241390 59537
rect 241334 59463 241390 59472
rect 240046 59392 240102 59401
rect 240046 59327 240102 59336
rect 241150 59392 241206 59401
rect 241150 59327 241206 59336
rect 239956 53100 240008 53106
rect 239956 53042 240008 53048
rect 238760 25764 238812 25770
rect 238760 25706 238812 25712
rect 238576 25560 238628 25566
rect 238576 25502 238628 25508
rect 238772 16574 238800 25706
rect 238772 16546 239352 16574
rect 238392 5160 238444 5166
rect 238392 5102 238444 5108
rect 239324 480 239352 16546
rect 240060 5098 240088 59327
rect 240140 51944 240192 51950
rect 240140 51886 240192 51892
rect 240048 5092 240100 5098
rect 240048 5034 240100 5040
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240152 354 240180 51886
rect 241164 4962 241192 59327
rect 241348 5030 241376 59463
rect 242530 59256 242586 59265
rect 242530 59191 242586 59200
rect 241704 14884 241756 14890
rect 241704 14826 241756 14832
rect 241336 5024 241388 5030
rect 241336 4966 241388 4972
rect 241152 4956 241204 4962
rect 241152 4898 241204 4904
rect 241716 480 241744 14826
rect 242544 4894 242572 59191
rect 242532 4888 242584 4894
rect 242532 4830 242584 4836
rect 242728 4826 242756 59706
rect 244186 59664 244242 59673
rect 244186 59599 244242 59608
rect 244200 51746 244228 59599
rect 245474 59528 245530 59537
rect 245474 59463 245530 59472
rect 245290 59392 245346 59401
rect 245290 59327 245346 59336
rect 244188 51740 244240 51746
rect 244188 51682 244240 51688
rect 244280 40860 244332 40866
rect 244280 40802 244332 40808
rect 242900 26920 242952 26926
rect 242900 26862 242952 26868
rect 242716 4820 242768 4826
rect 242716 4762 242768 4768
rect 242912 480 242940 26862
rect 242992 17332 243044 17338
rect 242992 17274 243044 17280
rect 243004 16574 243032 17274
rect 244292 16574 244320 40802
rect 245304 26926 245332 59327
rect 245488 50386 245516 59463
rect 246672 59424 246724 59430
rect 246672 59366 246724 59372
rect 245476 50380 245528 50386
rect 245476 50322 245528 50328
rect 246684 28286 246712 59366
rect 246854 59256 246910 59265
rect 246854 59191 246910 59200
rect 246868 49026 246896 59191
rect 246856 49020 246908 49026
rect 246856 48962 246908 48968
rect 248340 47598 248368 59706
rect 249706 59664 249762 59673
rect 249444 59622 249706 59650
rect 248878 59528 248934 59537
rect 248878 59463 248934 59472
rect 248892 59430 248920 59463
rect 248880 59424 248932 59430
rect 248880 59366 248932 59372
rect 248328 47592 248380 47598
rect 248328 47534 248380 47540
rect 249444 29646 249472 59622
rect 249706 59599 249762 59608
rect 250548 59401 250576 59735
rect 253202 59735 253204 59744
rect 251824 59706 251876 59712
rect 253256 59735 253258 59744
rect 257434 59800 257490 59809
rect 257434 59735 257490 59744
rect 267738 59800 267794 59809
rect 272706 59800 272762 59809
rect 267738 59735 267740 59744
rect 253204 59706 253256 59712
rect 251086 59528 251142 59537
rect 251086 59463 251142 59472
rect 249614 59392 249670 59401
rect 249614 59327 249670 59336
rect 250534 59392 250590 59401
rect 250534 59327 250590 59336
rect 250994 59392 251050 59401
rect 250994 59327 251050 59336
rect 249628 46238 249656 59327
rect 249616 46232 249668 46238
rect 249616 46174 249668 46180
rect 251008 44878 251036 59327
rect 250996 44872 251048 44878
rect 250996 44814 251048 44820
rect 251100 31074 251128 59463
rect 251180 55956 251232 55962
rect 251180 55898 251232 55904
rect 249800 31068 249852 31074
rect 249800 31010 249852 31016
rect 251088 31068 251140 31074
rect 251088 31010 251140 31016
rect 249432 29640 249484 29646
rect 249432 29582 249484 29588
rect 245660 28280 245712 28286
rect 245660 28222 245712 28228
rect 246672 28280 246724 28286
rect 246672 28222 246724 28228
rect 245292 26920 245344 26926
rect 245292 26862 245344 26868
rect 245672 16574 245700 28222
rect 247040 18828 247092 18834
rect 247040 18770 247092 18776
rect 247052 16574 247080 18770
rect 249812 16574 249840 31010
rect 243004 16546 244136 16574
rect 244292 16546 245240 16574
rect 245672 16546 245976 16574
rect 247052 16546 247632 16574
rect 249812 16546 250024 16574
rect 244108 480 244136 16546
rect 245212 480 245240 16546
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 16546
rect 247604 480 247632 16546
rect 248420 14952 248472 14958
rect 248420 14894 248472 14900
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248432 354 248460 14894
rect 249996 480 250024 16546
rect 251192 3806 251220 55898
rect 251836 24274 251864 59706
rect 257344 59696 257396 59702
rect 252282 59664 252338 59673
rect 252282 59599 252338 59608
rect 253386 59664 253442 59673
rect 253386 59599 253442 59608
rect 255594 59664 255650 59673
rect 257250 59664 257306 59673
rect 255594 59599 255650 59608
rect 255964 59628 256016 59634
rect 252296 59401 252324 59599
rect 252282 59392 252338 59401
rect 252282 59327 252338 59336
rect 253202 59392 253258 59401
rect 253202 59327 253258 59336
rect 251824 24268 251876 24274
rect 251824 24210 251876 24216
rect 253216 22914 253244 59327
rect 253400 53310 253428 59599
rect 254766 59528 254822 59537
rect 254766 59463 254822 59472
rect 254582 59256 254638 59265
rect 254582 59191 254638 59200
rect 253388 53304 253440 53310
rect 253388 53246 253440 53252
rect 254596 29782 254624 59191
rect 254780 51882 254808 59463
rect 255608 59401 255636 59599
rect 257344 59638 257396 59644
rect 257250 59599 257252 59608
rect 255964 59570 256016 59576
rect 257304 59599 257306 59608
rect 257252 59570 257304 59576
rect 255594 59392 255650 59401
rect 255594 59327 255650 59336
rect 254768 51876 254820 51882
rect 254768 51818 254820 51824
rect 254584 29776 254636 29782
rect 254584 29718 254636 29724
rect 253204 22908 253256 22914
rect 253204 22850 253256 22856
rect 255976 20126 256004 59570
rect 257356 21554 257384 59638
rect 257448 59401 257476 59735
rect 267792 59735 267794 59744
rect 269212 59764 269264 59770
rect 267740 59706 267792 59712
rect 276846 59800 276902 59809
rect 272706 59735 272708 59744
rect 269212 59706 269264 59712
rect 272760 59735 272762 59744
rect 274732 59764 274784 59770
rect 272708 59706 272760 59712
rect 280066 59800 280122 59809
rect 276846 59735 276848 59744
rect 274732 59706 274784 59712
rect 276900 59735 276902 59744
rect 278780 59764 278832 59770
rect 276848 59706 276900 59712
rect 280066 59735 280122 59744
rect 286782 59800 286838 59809
rect 286782 59735 286784 59744
rect 278780 59706 278832 59712
rect 258080 59696 258132 59702
rect 258080 59638 258132 59644
rect 258906 59664 258962 59673
rect 258092 59537 258120 59638
rect 258724 59628 258776 59634
rect 258906 59599 258962 59608
rect 260562 59664 260618 59673
rect 260562 59599 260564 59608
rect 258724 59570 258776 59576
rect 258078 59528 258134 59537
rect 258078 59463 258134 59472
rect 257434 59392 257490 59401
rect 257434 59327 257490 59336
rect 257526 59256 257582 59265
rect 257526 59191 257582 59200
rect 257540 31278 257568 59191
rect 257528 31272 257580 31278
rect 257528 31214 257580 31220
rect 257344 21548 257396 21554
rect 257344 21490 257396 21496
rect 255964 20120 256016 20126
rect 255964 20062 256016 20068
rect 255872 15020 255924 15026
rect 255872 14962 255924 14968
rect 251272 10532 251324 10538
rect 251272 10474 251324 10480
rect 251180 3800 251232 3806
rect 251180 3742 251232 3748
rect 251284 3482 251312 10474
rect 253480 6656 253532 6662
rect 253480 6598 253532 6604
rect 254676 6656 254728 6662
rect 254676 6598 254728 6604
rect 252376 3800 252428 3806
rect 252376 3742 252428 3748
rect 251192 3454 251312 3482
rect 251192 480 251220 3454
rect 252388 480 252416 3742
rect 253492 480 253520 6598
rect 254688 480 254716 6598
rect 255884 480 255912 14962
rect 258736 13394 258764 59570
rect 258920 59401 258948 59599
rect 260616 59599 260618 59608
rect 260564 59570 260616 59576
rect 260562 59528 260618 59537
rect 259000 59492 259052 59498
rect 260562 59463 260564 59472
rect 259000 59434 259052 59440
rect 260616 59463 260618 59472
rect 267738 59528 267794 59537
rect 268198 59528 268254 59537
rect 267794 59486 267872 59514
rect 267738 59463 267794 59472
rect 260564 59434 260616 59440
rect 258906 59392 258962 59401
rect 258906 59327 258962 59336
rect 259012 45554 259040 59434
rect 260102 59392 260158 59401
rect 260102 59327 260158 59336
rect 258920 45526 259040 45554
rect 258920 40934 258948 45526
rect 259460 42288 259512 42294
rect 259460 42230 259512 42236
rect 258908 40928 258960 40934
rect 258908 40870 258960 40876
rect 258724 13388 258776 13394
rect 258724 13330 258776 13336
rect 257068 6588 257120 6594
rect 257068 6530 257120 6536
rect 258264 6588 258316 6594
rect 258264 6530 258316 6536
rect 257080 480 257108 6530
rect 258276 480 258304 6530
rect 259472 480 259500 42230
rect 259552 32632 259604 32638
rect 259552 32574 259604 32580
rect 259564 6914 259592 32574
rect 260116 10470 260144 59327
rect 262126 59256 262182 59265
rect 262126 59191 262182 59200
rect 262034 59120 262090 59129
rect 262034 59055 262090 59064
rect 262048 56030 262076 59055
rect 262140 57390 262168 59191
rect 262128 57384 262180 57390
rect 262128 57326 262180 57332
rect 262036 56024 262088 56030
rect 262036 55966 262088 55972
rect 267740 56024 267792 56030
rect 267740 55966 267792 55972
rect 263600 43648 263652 43654
rect 263600 43590 263652 43596
rect 262220 35420 262272 35426
rect 262220 35362 262272 35368
rect 260840 20120 260892 20126
rect 260840 20062 260892 20068
rect 260852 16574 260880 20062
rect 262232 16574 262260 35362
rect 263612 16574 263640 43590
rect 266360 36780 266412 36786
rect 266360 36722 266412 36728
rect 266372 16574 266400 36722
rect 267752 16574 267780 55966
rect 267844 47802 267872 59486
rect 268198 59463 268254 59472
rect 268014 59256 268070 59265
rect 268014 59191 268070 59200
rect 268028 49230 268056 59191
rect 268212 58818 268240 59463
rect 268200 58812 268252 58818
rect 268200 58754 268252 58760
rect 268016 49224 268068 49230
rect 268016 49166 268068 49172
rect 267832 47796 267884 47802
rect 267832 47738 267884 47744
rect 269120 29776 269172 29782
rect 269120 29718 269172 29724
rect 260852 16546 261800 16574
rect 262232 16546 262536 16574
rect 263612 16546 264192 16574
rect 266372 16546 266584 16574
rect 267752 16546 268424 16574
rect 260104 10464 260156 10470
rect 260104 10406 260156 10412
rect 259564 6886 260696 6914
rect 260668 480 260696 6886
rect 261772 480 261800 16546
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 264164 480 264192 16546
rect 265348 6724 265400 6730
rect 265348 6666 265400 6672
rect 265360 480 265388 6666
rect 266556 480 266584 16546
rect 267740 6520 267792 6526
rect 267740 6462 267792 6468
rect 267752 480 267780 6462
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 16546
rect 269132 6914 269160 29718
rect 269224 15910 269252 59706
rect 271878 59528 271934 59537
rect 271878 59463 271934 59472
rect 270682 59256 270738 59265
rect 270682 59191 270738 59200
rect 270696 50590 270724 59191
rect 270684 50584 270736 50590
rect 270684 50526 270736 50532
rect 271892 46442 271920 59463
rect 271970 59392 272026 59401
rect 271970 59327 272026 59336
rect 271984 54738 272012 59327
rect 273350 59256 273406 59265
rect 273350 59191 273406 59200
rect 273260 57452 273312 57458
rect 273260 57394 273312 57400
rect 271972 54732 272024 54738
rect 271972 54674 272024 54680
rect 271880 46436 271932 46442
rect 271880 46378 271932 46384
rect 272432 16108 272484 16114
rect 272432 16050 272484 16056
rect 269212 15904 269264 15910
rect 269212 15846 269264 15852
rect 269132 6886 270080 6914
rect 270052 480 270080 6886
rect 271236 6452 271288 6458
rect 271236 6394 271288 6400
rect 271248 480 271276 6394
rect 272444 480 272472 16050
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273272 354 273300 57394
rect 273364 11762 273392 59191
rect 274744 45014 274772 59706
rect 276294 59528 276350 59537
rect 276294 59463 276350 59472
rect 274914 59256 274970 59265
rect 274914 59191 274970 59200
rect 276110 59256 276166 59265
rect 276110 59191 276166 59200
rect 274732 45008 274784 45014
rect 274732 44950 274784 44956
rect 274928 11830 274956 59191
rect 276124 11898 276152 59191
rect 276308 11966 276336 59463
rect 277398 59392 277454 59401
rect 277398 59327 277454 59336
rect 277412 57526 277440 59327
rect 277490 59256 277546 59265
rect 277490 59191 277546 59200
rect 277400 57520 277452 57526
rect 277400 57462 277452 57468
rect 277504 45554 277532 59191
rect 278792 56098 278820 59706
rect 280080 58886 280108 59735
rect 286836 59735 286838 59744
rect 287058 59800 287114 59809
rect 291842 59800 291898 59809
rect 287058 59735 287114 59744
rect 288440 59764 288492 59770
rect 286784 59706 286836 59712
rect 285126 59664 285182 59673
rect 285126 59599 285182 59608
rect 280158 59528 280214 59537
rect 280158 59463 280214 59472
rect 282642 59528 282698 59537
rect 282642 59463 282644 59472
rect 280068 58880 280120 58886
rect 280068 58822 280120 58828
rect 278780 56092 278832 56098
rect 278780 56034 278832 56040
rect 277412 45526 277532 45554
rect 277412 12034 277440 45526
rect 278044 38140 278096 38146
rect 278044 38082 278096 38088
rect 277400 12028 277452 12034
rect 277400 11970 277452 11976
rect 276296 11960 276348 11966
rect 276296 11902 276348 11908
rect 276112 11892 276164 11898
rect 276112 11834 276164 11840
rect 274916 11824 274968 11830
rect 274916 11766 274968 11772
rect 273352 11756 273404 11762
rect 273352 11698 273404 11704
rect 274824 6384 274876 6390
rect 274824 6326 274876 6332
rect 276020 6384 276072 6390
rect 276020 6326 276072 6332
rect 274836 480 274864 6326
rect 276032 480 276060 6326
rect 278056 4146 278084 38082
rect 280172 29850 280200 59463
rect 282696 59463 282698 59472
rect 284576 59492 284628 59498
rect 282644 59434 282696 59440
rect 284576 59434 284628 59440
rect 280342 59392 280398 59401
rect 280342 59327 280398 59336
rect 282918 59392 282974 59401
rect 282918 59327 282974 59336
rect 284390 59392 284446 59401
rect 284390 59327 284446 59336
rect 280160 29844 280212 29850
rect 280160 29786 280212 29792
rect 280160 21616 280212 21622
rect 280160 21558 280212 21564
rect 279056 11756 279108 11762
rect 279056 11698 279108 11704
rect 278320 6316 278372 6322
rect 278320 6258 278372 6264
rect 277124 4140 277176 4146
rect 277124 4082 277176 4088
rect 278044 4140 278096 4146
rect 278044 4082 278096 4088
rect 277136 480 277164 4082
rect 278332 480 278360 6258
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 354 279096 11698
rect 280172 6914 280200 21558
rect 280356 12102 280384 59327
rect 281538 59256 281594 59265
rect 281538 59191 281594 59200
rect 281552 16046 281580 59191
rect 282932 51950 282960 59327
rect 282920 51944 282972 51950
rect 282920 51886 282972 51892
rect 284404 18834 284432 59327
rect 284392 18828 284444 18834
rect 284392 18770 284444 18776
rect 284588 17338 284616 59434
rect 285140 59401 285168 59599
rect 285678 59528 285734 59537
rect 285678 59463 285734 59472
rect 285126 59392 285182 59401
rect 285126 59327 285182 59336
rect 284576 17332 284628 17338
rect 284576 17274 284628 17280
rect 281540 16040 281592 16046
rect 281540 15982 281592 15988
rect 280344 12096 280396 12102
rect 280344 12038 280396 12044
rect 283104 11824 283156 11830
rect 283104 11766 283156 11772
rect 280172 6886 280752 6914
rect 280724 480 280752 6886
rect 281908 6248 281960 6254
rect 281908 6190 281960 6196
rect 281920 480 281948 6190
rect 283116 480 283144 11766
rect 285692 10538 285720 59463
rect 287072 56030 287100 59735
rect 300122 59800 300178 59809
rect 291842 59735 291844 59744
rect 288440 59706 288492 59712
rect 291896 59735 291898 59744
rect 294144 59764 294196 59770
rect 291844 59706 291896 59712
rect 300122 59735 300124 59744
rect 294144 59706 294196 59712
rect 300176 59735 300178 59744
rect 300950 59800 301006 59809
rect 300950 59735 301006 59744
rect 301778 59800 301834 59809
rect 303434 59800 303490 59809
rect 301778 59735 301834 59744
rect 303068 59764 303120 59770
rect 300124 59706 300176 59712
rect 287426 59392 287482 59401
rect 287426 59327 287482 59336
rect 287242 59256 287298 59265
rect 287242 59191 287298 59200
rect 287060 56024 287112 56030
rect 287060 55966 287112 55972
rect 287152 15904 287204 15910
rect 287152 15846 287204 15852
rect 285680 10532 285732 10538
rect 285680 10474 285732 10480
rect 284300 10464 284352 10470
rect 284300 10406 284352 10412
rect 284312 480 284340 10406
rect 285404 6180 285456 6186
rect 285404 6122 285456 6128
rect 286600 6180 286652 6186
rect 286600 6122 286652 6128
rect 285416 480 285444 6122
rect 286612 480 286640 6122
rect 287164 490 287192 15846
rect 287256 6662 287284 59191
rect 287244 6656 287296 6662
rect 287244 6598 287296 6604
rect 287440 6594 287468 59327
rect 288452 20126 288480 59706
rect 293498 59664 293554 59673
rect 293498 59599 293500 59608
rect 293552 59599 293554 59608
rect 293500 59570 293552 59576
rect 288622 59528 288678 59537
rect 288622 59463 288678 59472
rect 291566 59528 291622 59537
rect 291566 59463 291622 59472
rect 294050 59528 294106 59537
rect 294050 59463 294106 59472
rect 288440 20120 288492 20126
rect 288440 20062 288492 20068
rect 288532 15972 288584 15978
rect 288532 15914 288584 15920
rect 287428 6588 287480 6594
rect 287428 6530 287480 6536
rect 288544 3482 288572 15914
rect 288636 6730 288664 59463
rect 291382 59256 291438 59265
rect 291382 59191 291438 59200
rect 291200 51876 291252 51882
rect 291200 51818 291252 51824
rect 289820 15224 289872 15230
rect 289820 15166 289872 15172
rect 288624 6724 288676 6730
rect 288624 6666 288676 6672
rect 288544 3454 289032 3482
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287164 462 287376 490
rect 289004 480 289032 3454
rect 287348 354 287376 462
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 289832 354 289860 15166
rect 291212 6914 291240 51818
rect 291396 16114 291424 59191
rect 291384 16108 291436 16114
rect 291384 16050 291436 16056
rect 291212 6886 291424 6914
rect 291396 480 291424 6886
rect 291580 6390 291608 59463
rect 292670 59392 292726 59401
rect 292670 59327 292726 59336
rect 292580 33992 292632 33998
rect 292580 33934 292632 33940
rect 291568 6384 291620 6390
rect 291568 6326 291620 6332
rect 292592 480 292620 33934
rect 292684 11762 292712 59327
rect 293960 20188 294012 20194
rect 293960 20130 294012 20136
rect 292672 11756 292724 11762
rect 292672 11698 292724 11704
rect 293684 5568 293736 5574
rect 293684 5510 293736 5516
rect 293696 480 293724 5510
rect 293972 3482 294000 20130
rect 294064 6186 294092 59463
rect 294156 11830 294184 59706
rect 295982 59664 296038 59673
rect 295524 59628 295576 59634
rect 295982 59599 296038 59608
rect 296810 59664 296866 59673
rect 296810 59599 296812 59608
rect 295524 59570 295576 59576
rect 295340 42152 295392 42158
rect 295340 42094 295392 42100
rect 294144 11824 294196 11830
rect 294144 11766 294196 11772
rect 295352 6914 295380 42094
rect 295536 15230 295564 59570
rect 295996 59401 296024 59599
rect 296864 59599 296866 59608
rect 298744 59628 298796 59634
rect 296812 59570 296864 59576
rect 298744 59570 298796 59576
rect 296718 59528 296774 59537
rect 296718 59463 296774 59472
rect 295982 59392 296038 59401
rect 295982 59327 296038 59336
rect 295706 59256 295762 59265
rect 295706 59191 295762 59200
rect 295524 15224 295576 15230
rect 295524 15166 295576 15172
rect 295352 6886 295656 6914
rect 294052 6180 294104 6186
rect 294052 6122 294104 6128
rect 293972 3454 294920 3482
rect 294892 480 294920 3454
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 295628 354 295656 6886
rect 295720 5574 295748 59191
rect 296732 16574 296760 59463
rect 296732 16546 297312 16574
rect 295708 5568 295760 5574
rect 295708 5510 295760 5516
rect 297284 480 297312 16546
rect 298100 15972 298152 15978
rect 298100 15914 298152 15920
rect 296046 354 296158 480
rect 295628 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298112 354 298140 15914
rect 298756 5642 298784 59570
rect 300122 59528 300178 59537
rect 300122 59463 300178 59472
rect 298926 59256 298982 59265
rect 298926 59191 298982 59200
rect 298744 5636 298796 5642
rect 298744 5578 298796 5584
rect 298940 5574 298968 59191
rect 299480 35284 299532 35290
rect 299480 35226 299532 35232
rect 299492 16574 299520 35226
rect 299492 16546 299704 16574
rect 298928 5568 298980 5574
rect 298928 5510 298980 5516
rect 299676 480 299704 16546
rect 300136 6662 300164 59463
rect 300964 59401 300992 59735
rect 301792 59702 301820 59735
rect 303434 59735 303436 59744
rect 303068 59706 303120 59712
rect 303488 59735 303490 59744
rect 305366 59800 305422 59809
rect 305826 59800 305882 59809
rect 305366 59735 305422 59744
rect 305736 59764 305788 59770
rect 303436 59706 303488 59712
rect 301780 59696 301832 59702
rect 301502 59664 301558 59673
rect 301780 59638 301832 59644
rect 301502 59599 301558 59608
rect 300950 59392 301006 59401
rect 300950 59327 301006 59336
rect 300306 59256 300362 59265
rect 300306 59191 300362 59200
rect 300320 12442 300348 59191
rect 300308 12436 300360 12442
rect 300308 12378 300360 12384
rect 300124 6656 300176 6662
rect 300124 6598 300176 6604
rect 301516 6594 301544 59599
rect 302882 59392 302938 59401
rect 302882 59327 302938 59336
rect 302240 36644 302292 36650
rect 302240 36586 302292 36592
rect 302252 16574 302280 36586
rect 302252 16546 302832 16574
rect 301504 6588 301556 6594
rect 301504 6530 301556 6536
rect 300768 5568 300820 5574
rect 300768 5510 300820 5516
rect 300780 480 300808 5510
rect 302804 3482 302832 16546
rect 302896 6458 302924 59327
rect 303080 6526 303108 59706
rect 304448 59696 304500 59702
rect 304448 59638 304500 59644
rect 304262 59528 304318 59537
rect 304262 59463 304318 59472
rect 303068 6520 303120 6526
rect 303068 6462 303120 6468
rect 302884 6452 302936 6458
rect 302884 6394 302936 6400
rect 304276 6322 304304 59463
rect 304460 6390 304488 59638
rect 305380 59401 305408 59735
rect 305826 59735 305882 59744
rect 309322 59800 309378 59809
rect 309322 59735 309378 59744
rect 310702 59800 310758 59809
rect 310702 59735 310704 59744
rect 305736 59706 305788 59712
rect 305366 59392 305422 59401
rect 305366 59327 305422 59336
rect 305644 58880 305696 58886
rect 305644 58822 305696 58828
rect 305552 16040 305604 16046
rect 305552 15982 305604 15988
rect 304448 6384 304500 6390
rect 304448 6326 304500 6332
rect 304264 6316 304316 6322
rect 304264 6258 304316 6264
rect 304356 5636 304408 5642
rect 304356 5578 304408 5584
rect 302804 3454 303200 3482
rect 301964 3392 302016 3398
rect 301964 3334 302016 3340
rect 301976 480 302004 3334
rect 303172 480 303200 3454
rect 304368 480 304396 5578
rect 305564 480 305592 15982
rect 305656 3398 305684 58822
rect 305748 17338 305776 59706
rect 305840 58818 305868 59735
rect 305918 59664 305974 59673
rect 305918 59599 305920 59608
rect 305972 59599 305974 59608
rect 307024 59628 307076 59634
rect 305920 59570 305972 59576
rect 307024 59570 307076 59576
rect 306746 59528 306802 59537
rect 306746 59463 306748 59472
rect 306800 59463 306802 59472
rect 306748 59434 306800 59440
rect 305828 58812 305880 58818
rect 305828 58754 305880 58760
rect 306380 38004 306432 38010
rect 306380 37946 306432 37952
rect 305736 17332 305788 17338
rect 305736 17274 305788 17280
rect 305644 3392 305696 3398
rect 305644 3334 305696 3340
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306392 354 306420 37946
rect 307036 6254 307064 59570
rect 307760 59492 307812 59498
rect 307760 59434 307812 59440
rect 307206 59392 307262 59401
rect 307206 59327 307262 59336
rect 307024 6248 307076 6254
rect 307024 6190 307076 6196
rect 307220 6186 307248 59327
rect 307772 57390 307800 59434
rect 309336 59401 309364 59735
rect 310756 59735 310758 59744
rect 311806 59800 311862 59809
rect 313462 59800 313518 59809
rect 311806 59735 311862 59744
rect 312544 59764 312596 59770
rect 310704 59706 310756 59712
rect 309874 59528 309930 59537
rect 309874 59463 309930 59472
rect 310702 59528 310758 59537
rect 310702 59463 310758 59472
rect 309322 59392 309378 59401
rect 309322 59327 309378 59336
rect 307760 57384 307812 57390
rect 307760 57326 307812 57332
rect 309140 39500 309192 39506
rect 309140 39442 309192 39448
rect 309784 39500 309836 39506
rect 309784 39442 309836 39448
rect 307944 12436 307996 12442
rect 307944 12378 307996 12384
rect 307208 6180 307260 6186
rect 307208 6122 307260 6128
rect 307956 480 307984 12378
rect 309152 6914 309180 39442
rect 309796 16574 309824 39442
rect 309888 29918 309916 59463
rect 310716 55214 310744 59463
rect 311820 59401 311848 59735
rect 313462 59735 313518 59744
rect 314290 59800 314292 59809
rect 315396 59832 315448 59838
rect 314344 59800 314346 59809
rect 314290 59735 314346 59744
rect 315394 59800 315396 59809
rect 357532 59832 357584 59838
rect 315448 59800 315450 59809
rect 315394 59735 315450 59744
rect 316590 59800 316646 59809
rect 318430 59800 318486 59809
rect 316646 59758 316816 59786
rect 316590 59735 316646 59744
rect 312544 59706 312596 59712
rect 311346 59392 311402 59401
rect 311346 59327 311402 59336
rect 311806 59392 311862 59401
rect 311806 59327 311862 59336
rect 310716 55186 311204 55214
rect 309876 29912 309928 29918
rect 309876 29854 309928 29860
rect 309796 16546 309916 16574
rect 309152 6886 309824 6914
rect 309048 3392 309100 3398
rect 309048 3334 309100 3340
rect 309060 480 309088 3334
rect 306718 354 306830 480
rect 306392 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 6886
rect 309888 3398 309916 16546
rect 311176 7954 311204 55186
rect 311164 7948 311216 7954
rect 311164 7890 311216 7896
rect 311360 7886 311388 59327
rect 311900 28484 311952 28490
rect 311900 28426 311952 28432
rect 311912 16574 311940 28426
rect 311912 16546 312216 16574
rect 311348 7880 311400 7886
rect 311348 7822 311400 7828
rect 311440 6656 311492 6662
rect 311440 6598 311492 6604
rect 309876 3392 309928 3398
rect 309876 3334 309928 3340
rect 311452 480 311480 6598
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312188 354 312216 16546
rect 312556 7818 312584 59706
rect 312726 59528 312782 59537
rect 312726 59463 312782 59472
rect 312740 8226 312768 59463
rect 313476 59401 313504 59735
rect 314290 59664 314346 59673
rect 316590 59664 316646 59673
rect 314346 59622 314700 59650
rect 314290 59599 314346 59608
rect 313462 59392 313518 59401
rect 313462 59327 313518 59336
rect 313922 59256 313978 59265
rect 313922 59191 313978 59200
rect 313280 40792 313332 40798
rect 313280 40734 313332 40740
rect 313292 16574 313320 40734
rect 313292 16546 313872 16574
rect 312728 8220 312780 8226
rect 312728 8162 312780 8168
rect 312544 7812 312596 7818
rect 312544 7754 312596 7760
rect 313844 480 313872 16546
rect 313936 10538 313964 59191
rect 314672 56098 314700 59622
rect 316590 59599 316592 59608
rect 316644 59599 316646 59608
rect 316592 59570 316644 59576
rect 316590 59528 316646 59537
rect 316646 59486 316724 59514
rect 316590 59463 316646 59472
rect 315302 59392 315358 59401
rect 315302 59327 315358 59336
rect 314660 56092 314712 56098
rect 314660 56034 314712 56040
rect 315316 51950 315344 59327
rect 315304 51944 315356 51950
rect 315304 51886 315356 51892
rect 316040 51808 316092 51814
rect 316040 51750 316092 51756
rect 313924 10532 313976 10538
rect 313924 10474 313976 10480
rect 315028 6588 315080 6594
rect 315028 6530 315080 6536
rect 315040 480 315068 6530
rect 316052 3398 316080 51750
rect 316696 22982 316724 59486
rect 316788 55214 316816 59758
rect 318430 59735 318432 59744
rect 318484 59735 318486 59744
rect 319258 59800 319314 59809
rect 319258 59735 319314 59744
rect 320822 59800 320878 59809
rect 325054 59800 325110 59809
rect 320822 59735 320878 59744
rect 320916 59764 320968 59770
rect 318432 59706 318484 59712
rect 319272 59702 319300 59735
rect 320836 59702 320864 59735
rect 325054 59735 325110 59744
rect 325882 59800 325938 59809
rect 325882 59735 325938 59744
rect 326710 59800 326766 59809
rect 330114 59800 330170 59809
rect 326710 59735 326712 59744
rect 320916 59706 320968 59712
rect 319260 59696 319312 59702
rect 319260 59638 319312 59644
rect 320180 59696 320232 59702
rect 320180 59638 320232 59644
rect 320824 59696 320876 59702
rect 320824 59638 320876 59644
rect 318064 59628 318116 59634
rect 318064 59570 318116 59576
rect 316788 55186 316908 55214
rect 316880 45082 316908 55186
rect 316868 45076 316920 45082
rect 316868 45018 316920 45024
rect 318076 24342 318104 59570
rect 319442 59528 319498 59537
rect 319442 59463 319498 59472
rect 319456 29850 319484 59463
rect 319626 59392 319682 59401
rect 319626 59327 319682 59336
rect 319640 40934 319668 59327
rect 320192 56030 320220 59638
rect 320180 56024 320232 56030
rect 320180 55966 320232 55972
rect 320824 53304 320876 53310
rect 320824 53246 320876 53252
rect 319628 40928 319680 40934
rect 319628 40870 319680 40876
rect 319444 29844 319496 29850
rect 319444 29786 319496 29792
rect 320180 29708 320232 29714
rect 320180 29650 320232 29656
rect 318064 24336 318116 24342
rect 318064 24278 318116 24284
rect 316684 22976 316736 22982
rect 316684 22918 316736 22924
rect 320192 16574 320220 29650
rect 320192 16546 320496 16574
rect 316224 16108 316276 16114
rect 316224 16050 316276 16056
rect 316040 3392 316092 3398
rect 316040 3334 316092 3340
rect 316236 480 316264 16050
rect 318524 6520 318576 6526
rect 318524 6462 318576 6468
rect 317328 3392 317380 3398
rect 317328 3334 317380 3340
rect 317340 480 317368 3334
rect 318536 480 318564 6462
rect 319720 3256 319772 3262
rect 319720 3198 319772 3204
rect 319732 480 319760 3198
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 320836 3262 320864 53246
rect 320928 32638 320956 59706
rect 325068 59702 325096 59735
rect 322940 59696 322992 59702
rect 322940 59638 322992 59644
rect 325056 59696 325108 59702
rect 325056 59638 325108 59644
rect 321742 59528 321798 59537
rect 321742 59463 321744 59472
rect 321796 59463 321798 59472
rect 321744 59434 321796 59440
rect 321742 59392 321798 59401
rect 321742 59327 321798 59336
rect 321756 51074 321784 59327
rect 322952 51814 322980 59638
rect 324962 59528 325018 59537
rect 323584 59492 323636 59498
rect 324962 59463 325018 59472
rect 323584 59434 323636 59440
rect 322940 51808 322992 51814
rect 322940 51750 322992 51756
rect 321756 51046 322244 51074
rect 320916 32632 320968 32638
rect 320916 32574 320968 32580
rect 322216 18834 322244 51046
rect 322940 43648 322992 43654
rect 322940 43590 322992 43596
rect 322204 18828 322256 18834
rect 322204 18770 322256 18776
rect 322112 6452 322164 6458
rect 322112 6394 322164 6400
rect 320824 3256 320876 3262
rect 320824 3198 320876 3204
rect 322124 480 322152 6394
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 322952 354 322980 43590
rect 323596 12306 323624 59434
rect 324320 32564 324372 32570
rect 324320 32506 324372 32512
rect 324332 16574 324360 32506
rect 324332 16546 324452 16574
rect 323584 12300 323636 12306
rect 323584 12242 323636 12248
rect 324424 480 324452 16546
rect 324976 12170 325004 59463
rect 325896 59401 325924 59735
rect 326764 59735 326766 59744
rect 329104 59764 329156 59770
rect 326712 59706 326764 59712
rect 330942 59800 330998 59809
rect 330114 59735 330170 59744
rect 330852 59764 330904 59770
rect 329104 59706 329156 59712
rect 327724 59696 327776 59702
rect 326342 59664 326398 59673
rect 327724 59638 327776 59644
rect 328366 59664 328422 59673
rect 326342 59599 326398 59608
rect 325054 59392 325110 59401
rect 325054 59327 325110 59336
rect 325882 59392 325938 59401
rect 325882 59327 325938 59336
rect 325068 51074 325096 59327
rect 325068 51046 325188 51074
rect 325160 12238 325188 51046
rect 326356 39574 326384 59599
rect 326344 39568 326396 39574
rect 326344 39510 326396 39516
rect 327080 22840 327132 22846
rect 327080 22782 327132 22788
rect 325148 12232 325200 12238
rect 325148 12174 325200 12180
rect 324964 12164 325016 12170
rect 324964 12106 325016 12112
rect 327092 6914 327120 22782
rect 327736 12102 327764 59638
rect 328366 59599 328422 59608
rect 328380 59401 328408 59599
rect 327906 59392 327962 59401
rect 327906 59327 327962 59336
rect 328366 59392 328422 59401
rect 328366 59327 328422 59336
rect 327724 12096 327776 12102
rect 327724 12038 327776 12044
rect 327920 12034 327948 59327
rect 327908 12028 327960 12034
rect 327908 11970 327960 11976
rect 329116 11966 329144 59706
rect 329286 59528 329342 59537
rect 329286 59463 329342 59472
rect 329104 11960 329156 11966
rect 329104 11902 329156 11908
rect 329300 11898 329328 59463
rect 330128 59401 330156 59735
rect 337382 59800 337438 59809
rect 330942 59735 330998 59744
rect 331680 59764 331732 59770
rect 330852 59706 330904 59712
rect 330864 59673 330892 59706
rect 330956 59702 330984 59735
rect 337382 59735 337438 59744
rect 337566 59800 337622 59809
rect 341614 59800 341670 59809
rect 337566 59735 337568 59744
rect 331680 59706 331732 59712
rect 330944 59696 330996 59702
rect 330850 59664 330906 59673
rect 330944 59638 330996 59644
rect 330850 59599 330906 59608
rect 330482 59528 330538 59537
rect 330482 59463 330538 59472
rect 330114 59392 330170 59401
rect 330114 59327 330170 59336
rect 329840 22908 329892 22914
rect 329840 22850 329892 22856
rect 329852 16574 329880 22850
rect 329852 16546 330432 16574
rect 329288 11892 329340 11898
rect 329288 11834 329340 11840
rect 327092 6886 328040 6914
rect 325608 6384 325660 6390
rect 325608 6326 325660 6332
rect 325620 480 325648 6326
rect 326804 3324 326856 3330
rect 326804 3266 326856 3272
rect 326816 480 326844 3266
rect 328012 480 328040 6886
rect 329196 6316 329248 6322
rect 329196 6258 329248 6264
rect 329208 480 329236 6258
rect 330404 480 330432 16546
rect 330496 11830 330524 59463
rect 331692 51074 331720 59706
rect 333336 59696 333388 59702
rect 333336 59638 333388 59644
rect 335082 59664 335138 59673
rect 331770 59528 331826 59537
rect 331770 59463 331772 59472
rect 331824 59463 331826 59472
rect 333244 59492 333296 59498
rect 331772 59434 331824 59440
rect 333244 59434 333296 59440
rect 331770 59392 331826 59401
rect 331826 59350 331996 59378
rect 331770 59327 331826 59336
rect 331968 51074 331996 59350
rect 331692 51046 331904 51074
rect 331968 51046 332088 51074
rect 330576 50584 330628 50590
rect 330576 50526 330628 50532
rect 330484 11824 330536 11830
rect 330484 11766 330536 11772
rect 330588 3330 330616 50526
rect 331220 43580 331272 43586
rect 331220 43522 331272 43528
rect 330576 3324 330628 3330
rect 330576 3266 330628 3272
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331232 354 331260 43522
rect 331876 11762 331904 51046
rect 332060 22846 332088 51046
rect 332048 22840 332100 22846
rect 332048 22782 332100 22788
rect 333256 20126 333284 59434
rect 333348 51074 333376 59638
rect 335082 59599 335138 59608
rect 333426 59528 333482 59537
rect 333426 59463 333428 59472
rect 333480 59463 333482 59472
rect 333428 59434 333480 59440
rect 335096 59401 335124 59599
rect 336002 59528 336058 59537
rect 336002 59463 336058 59472
rect 336096 59492 336148 59498
rect 334622 59392 334678 59401
rect 334622 59327 334678 59336
rect 335082 59392 335138 59401
rect 335082 59327 335138 59336
rect 333348 51046 333468 51074
rect 333440 45014 333468 51046
rect 333428 45008 333480 45014
rect 333428 44950 333480 44956
rect 333980 44940 334032 44946
rect 333980 44882 334032 44888
rect 333244 20120 333296 20126
rect 333244 20062 333296 20068
rect 332600 17332 332652 17338
rect 332600 17274 332652 17280
rect 332612 16574 332640 17274
rect 333992 16574 334020 44882
rect 334636 21554 334664 59327
rect 336016 24274 336044 59463
rect 336096 59434 336148 59440
rect 336108 46442 336136 59434
rect 337396 59401 337424 59735
rect 337620 59735 337622 59744
rect 340328 59764 340380 59770
rect 337568 59706 337620 59712
rect 341614 59735 341670 59744
rect 345018 59800 345074 59809
rect 350630 59800 350686 59809
rect 345018 59735 345020 59744
rect 340328 59706 340380 59712
rect 337474 59664 337530 59673
rect 337474 59599 337530 59608
rect 339222 59664 339278 59673
rect 339222 59599 339278 59608
rect 337198 59392 337254 59401
rect 337198 59327 337254 59336
rect 337382 59392 337438 59401
rect 337382 59327 337438 59336
rect 337212 51074 337240 59327
rect 337212 51046 337424 51074
rect 336096 46436 336148 46442
rect 336096 46378 336148 46384
rect 336096 33992 336148 33998
rect 336096 33934 336148 33940
rect 336004 24268 336056 24274
rect 336004 24210 336056 24216
rect 334624 21548 334676 21554
rect 334624 21490 334676 21496
rect 332612 16546 332732 16574
rect 333992 16546 334664 16574
rect 331864 11756 331916 11762
rect 331864 11698 331916 11704
rect 332704 480 332732 16546
rect 333888 4140 333940 4146
rect 333888 4082 333940 4088
rect 333900 480 333928 4082
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 336108 4146 336136 33934
rect 337396 25770 337424 51046
rect 337488 47802 337516 59599
rect 339236 59401 339264 59599
rect 340142 59528 340198 59537
rect 340142 59463 340198 59472
rect 338854 59392 338910 59401
rect 338854 59327 338910 59336
rect 339222 59392 339278 59401
rect 339222 59327 339278 59336
rect 338764 49224 338816 49230
rect 338764 49166 338816 49172
rect 337476 47796 337528 47802
rect 337476 47738 337528 47744
rect 337384 25764 337436 25770
rect 337384 25706 337436 25712
rect 338120 24200 338172 24206
rect 338120 24142 338172 24148
rect 338132 16574 338160 24142
rect 338132 16546 338712 16574
rect 336280 6248 336332 6254
rect 336280 6190 336332 6196
rect 336096 4140 336148 4146
rect 336096 4082 336148 4088
rect 336292 480 336320 6190
rect 337476 3188 337528 3194
rect 337476 3130 337528 3136
rect 337488 480 337516 3130
rect 338684 480 338712 16546
rect 338776 3194 338804 49166
rect 338868 27130 338896 59327
rect 338856 27124 338908 27130
rect 338856 27066 338908 27072
rect 340156 6662 340184 59463
rect 340340 13394 340368 59706
rect 341522 59664 341578 59673
rect 341522 59599 341578 59608
rect 340880 33856 340932 33862
rect 340880 33798 340932 33804
rect 340328 13388 340380 13394
rect 340328 13330 340380 13336
rect 340144 6656 340196 6662
rect 340144 6598 340196 6604
rect 339868 6180 339920 6186
rect 339868 6122 339920 6128
rect 338764 3188 338816 3194
rect 338764 3130 338816 3136
rect 339880 480 339908 6122
rect 340892 1426 340920 33798
rect 340972 16176 341024 16182
rect 340972 16118 341024 16124
rect 340880 1420 340932 1426
rect 340880 1362 340932 1368
rect 340984 480 341012 16118
rect 341536 6526 341564 59599
rect 341628 59537 341656 59735
rect 345072 59735 345074 59744
rect 347044 59764 347096 59770
rect 345020 59706 345072 59712
rect 350630 59735 350686 59744
rect 351734 59800 351790 59809
rect 351734 59735 351790 59744
rect 356702 59800 356758 59809
rect 356702 59735 356704 59744
rect 347044 59706 347096 59712
rect 342350 59664 342406 59673
rect 342350 59599 342352 59608
rect 342404 59599 342406 59608
rect 343362 59664 343418 59673
rect 345018 59664 345074 59673
rect 343362 59599 343418 59608
rect 344468 59628 344520 59634
rect 342352 59570 342404 59576
rect 341614 59528 341670 59537
rect 341614 59463 341670 59472
rect 343376 59401 343404 59599
rect 345074 59622 345152 59650
rect 345018 59599 345074 59608
rect 344468 59570 344520 59576
rect 344282 59528 344338 59537
rect 344282 59463 344338 59472
rect 341614 59392 341670 59401
rect 341614 59327 341670 59336
rect 342902 59392 342958 59401
rect 342902 59327 342958 59336
rect 343362 59392 343418 59401
rect 343362 59327 343418 59336
rect 341628 55214 341656 59327
rect 342260 58812 342312 58818
rect 342260 58754 342312 58760
rect 341628 55186 341748 55214
rect 341720 6594 341748 55186
rect 342272 6914 342300 58754
rect 342916 16574 342944 59327
rect 344296 32570 344324 59463
rect 344480 40798 344508 59570
rect 345018 59392 345074 59401
rect 345018 59327 345074 59336
rect 345032 55214 345060 59327
rect 345124 58562 345152 59622
rect 345124 58534 345796 58562
rect 345768 55214 345796 58534
rect 346400 57384 346452 57390
rect 346400 57326 346452 57332
rect 345032 55186 345704 55214
rect 345768 55186 345888 55214
rect 344468 40792 344520 40798
rect 344468 40734 344520 40740
rect 344284 32564 344336 32570
rect 344284 32506 344336 32512
rect 343640 31272 343692 31278
rect 343640 31214 343692 31220
rect 343652 16574 343680 31214
rect 342916 16546 343036 16574
rect 343652 16546 344600 16574
rect 342272 6886 342944 6914
rect 341708 6588 341760 6594
rect 341708 6530 341760 6536
rect 341524 6520 341576 6526
rect 341524 6462 341576 6468
rect 342168 1420 342220 1426
rect 342168 1362 342220 1368
rect 342180 480 342208 1362
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 6886
rect 343008 6458 343036 16546
rect 342996 6452 343048 6458
rect 342996 6394 343048 6400
rect 344572 480 344600 16546
rect 345676 6390 345704 55186
rect 345756 7744 345808 7750
rect 345756 7686 345808 7692
rect 345664 6384 345716 6390
rect 345664 6326 345716 6332
rect 345768 480 345796 7686
rect 345860 6322 345888 55186
rect 346412 16574 346440 57326
rect 346412 16546 346992 16574
rect 345848 6316 345900 6322
rect 345848 6258 345900 6264
rect 346964 480 346992 16546
rect 347056 6254 347084 59706
rect 347502 59528 347558 59537
rect 347502 59463 347504 59472
rect 347556 59463 347558 59472
rect 349802 59528 349858 59537
rect 349802 59463 349858 59472
rect 349988 59492 350040 59498
rect 347504 59434 347556 59440
rect 348606 59392 348662 59401
rect 348606 59327 348662 59336
rect 348422 59256 348478 59265
rect 348422 59191 348478 59200
rect 347044 6248 347096 6254
rect 347044 6190 347096 6196
rect 348436 6186 348464 59191
rect 348620 43586 348648 59327
rect 348608 43580 348660 43586
rect 348608 43522 348660 43528
rect 349160 29912 349212 29918
rect 349160 29854 349212 29860
rect 348424 6180 348476 6186
rect 348424 6122 348476 6128
rect 348056 3188 348108 3194
rect 348056 3130 348108 3136
rect 348068 480 348096 3130
rect 349172 1426 349200 29854
rect 349816 17338 349844 59463
rect 349988 59434 350040 59440
rect 350000 33862 350028 59434
rect 350644 59022 350672 59735
rect 350906 59664 350962 59673
rect 350906 59599 350962 59608
rect 350632 59016 350684 59022
rect 350632 58958 350684 58964
rect 350920 51074 350948 59599
rect 351748 58818 351776 59735
rect 356756 59735 356758 59744
rect 357530 59800 357532 59809
rect 359464 59832 359516 59838
rect 357584 59800 357586 59809
rect 422392 59832 422444 59838
rect 359464 59774 359516 59780
rect 360842 59800 360898 59809
rect 357530 59735 357586 59744
rect 356704 59706 356756 59712
rect 353390 59664 353446 59673
rect 353390 59599 353392 59608
rect 353444 59599 353446 59608
rect 354218 59664 354274 59673
rect 357530 59664 357586 59673
rect 354218 59599 354274 59608
rect 354680 59628 354732 59634
rect 353392 59570 353444 59576
rect 354034 59528 354090 59537
rect 354034 59463 354090 59472
rect 352288 59016 352340 59022
rect 352288 58958 352340 58964
rect 352746 58984 352802 58993
rect 351736 58812 351788 58818
rect 351736 58754 351788 58760
rect 352300 51074 352328 58958
rect 352746 58919 352802 58928
rect 352760 51074 352788 58919
rect 353944 54732 353996 54738
rect 353944 54674 353996 54680
rect 350920 51046 351224 51074
rect 352300 51046 352696 51074
rect 352760 51046 352880 51074
rect 351196 35290 351224 51046
rect 352564 44940 352616 44946
rect 352564 44882 352616 44888
rect 351184 35284 351236 35290
rect 351184 35226 351236 35232
rect 349988 33856 350040 33862
rect 349988 33798 350040 33804
rect 349804 17332 349856 17338
rect 349804 17274 349856 17280
rect 349252 7676 349304 7682
rect 349252 7618 349304 7624
rect 349160 1420 349212 1426
rect 349160 1362 349212 1368
rect 349264 480 349292 7618
rect 351644 3324 351696 3330
rect 351644 3266 351696 3272
rect 350448 1420 350500 1426
rect 350448 1362 350500 1368
rect 350460 480 350488 1362
rect 351656 480 351684 3266
rect 352576 3194 352604 44882
rect 352668 36650 352696 51046
rect 352852 42158 352880 51046
rect 352840 42152 352892 42158
rect 352840 42094 352892 42100
rect 352656 36644 352708 36650
rect 352656 36586 352708 36592
rect 352840 7608 352892 7614
rect 352840 7550 352892 7556
rect 352564 3188 352616 3194
rect 352564 3130 352616 3136
rect 352852 480 352880 7550
rect 353956 3330 353984 54674
rect 354048 38010 354076 59463
rect 354232 59401 354260 59599
rect 357530 59599 357586 59608
rect 354680 59570 354732 59576
rect 354218 59392 354274 59401
rect 354218 59327 354274 59336
rect 354692 57390 354720 59570
rect 356702 59528 356758 59537
rect 356702 59463 356758 59472
rect 354680 57384 354732 57390
rect 354680 57326 354732 57332
rect 354036 38004 354088 38010
rect 354036 37946 354088 37952
rect 356060 17468 356112 17474
rect 356060 17410 356112 17416
rect 356072 16574 356100 17410
rect 356072 16546 356376 16574
rect 354036 7948 354088 7954
rect 354036 7890 354088 7896
rect 353944 3324 353996 3330
rect 353944 3266 353996 3272
rect 354048 480 354076 7890
rect 355232 3052 355284 3058
rect 355232 2994 355284 3000
rect 355244 480 355272 2994
rect 356348 480 356376 16546
rect 356716 8294 356744 59463
rect 356886 59256 356942 59265
rect 356886 59191 356942 59200
rect 356704 8288 356756 8294
rect 356704 8230 356756 8236
rect 356900 8158 356928 59191
rect 357544 51074 357572 59599
rect 357544 51046 358124 51074
rect 357440 18896 357492 18902
rect 357440 18838 357492 18844
rect 356888 8152 356940 8158
rect 356888 8094 356940 8100
rect 357452 3398 357480 18838
rect 358096 8090 358124 51046
rect 358820 35352 358872 35358
rect 358820 35294 358872 35300
rect 358176 29708 358228 29714
rect 358176 29650 358228 29656
rect 358084 8084 358136 8090
rect 358084 8026 358136 8032
rect 357532 7880 357584 7886
rect 357532 7822 357584 7828
rect 357440 3392 357492 3398
rect 357440 3334 357492 3340
rect 357544 480 357572 7822
rect 358188 3058 358216 29650
rect 358832 6914 358860 35294
rect 359476 8022 359504 59774
rect 359648 59764 359700 59770
rect 360842 59735 360844 59744
rect 359648 59706 359700 59712
rect 360896 59735 360898 59744
rect 361578 59800 361634 59809
rect 369122 59800 369178 59809
rect 361578 59735 361634 59744
rect 363604 59764 363656 59770
rect 360844 59706 360896 59712
rect 359464 8016 359516 8022
rect 359464 7958 359516 7964
rect 359660 7954 359688 59706
rect 360108 59628 360160 59634
rect 360108 59570 360160 59576
rect 361028 59628 361080 59634
rect 361028 59570 361080 59576
rect 360120 59401 360148 59570
rect 360842 59528 360898 59537
rect 360842 59463 360898 59472
rect 360106 59392 360162 59401
rect 360106 59327 360162 59336
rect 359648 7948 359700 7954
rect 359648 7890 359700 7896
rect 360856 7750 360884 59463
rect 361040 7886 361068 59570
rect 361592 59401 361620 59735
rect 369122 59735 369178 59744
rect 369490 59800 369546 59809
rect 376482 59800 376538 59809
rect 369490 59735 369546 59744
rect 373816 59764 373868 59770
rect 363604 59706 363656 59712
rect 361670 59664 361726 59673
rect 361670 59599 361726 59608
rect 361578 59392 361634 59401
rect 361578 59327 361634 59336
rect 361684 55214 361712 59599
rect 362498 59528 362554 59537
rect 362498 59463 362500 59472
rect 362552 59463 362554 59472
rect 362500 59434 362552 59440
rect 363050 59256 363106 59265
rect 363050 59191 363106 59200
rect 361684 55186 362264 55214
rect 361488 8288 361540 8294
rect 361488 8230 361540 8236
rect 361500 8090 361528 8230
rect 361488 8084 361540 8090
rect 361488 8026 361540 8032
rect 361224 7954 361436 7970
rect 361212 7948 361448 7954
rect 361264 7942 361396 7948
rect 361212 7890 361264 7896
rect 361396 7890 361448 7896
rect 361028 7880 361080 7886
rect 361028 7822 361080 7828
rect 361120 7812 361172 7818
rect 361120 7754 361172 7760
rect 360844 7744 360896 7750
rect 360844 7686 360896 7692
rect 358832 6886 359504 6914
rect 358728 3392 358780 3398
rect 358728 3334 358780 3340
rect 358176 3052 358228 3058
rect 358176 2994 358228 3000
rect 358740 480 358768 3334
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 6886
rect 361132 480 361160 7754
rect 362236 7682 362264 55186
rect 362960 42220 363012 42226
rect 362960 42162 363012 42168
rect 362972 16574 363000 42162
rect 363064 28354 363092 59191
rect 363052 28348 363104 28354
rect 363052 28290 363104 28296
rect 362972 16546 363552 16574
rect 362224 7676 362276 7682
rect 362224 7618 362276 7624
rect 362316 4004 362368 4010
rect 362316 3946 362368 3952
rect 362328 480 362356 3946
rect 363524 480 363552 16546
rect 363616 7614 363644 59706
rect 369030 59664 369086 59673
rect 369030 59599 369032 59608
rect 369084 59599 369086 59608
rect 369032 59570 369084 59576
rect 364798 59528 364854 59537
rect 364432 59492 364484 59498
rect 366638 59528 366694 59537
rect 364798 59463 364800 59472
rect 364432 59434 364484 59440
rect 364852 59463 364854 59472
rect 365720 59492 365772 59498
rect 364800 59434 364852 59440
rect 366638 59463 366640 59472
rect 365720 59434 365772 59440
rect 366692 59463 366694 59472
rect 368478 59528 368534 59537
rect 368478 59463 368534 59472
rect 368572 59492 368624 59498
rect 366640 59434 366692 59440
rect 364338 59392 364394 59401
rect 364338 59327 364394 59336
rect 364352 18698 364380 59327
rect 364444 25634 364472 59434
rect 365732 46306 365760 59434
rect 367282 59392 367338 59401
rect 367282 59327 367338 59336
rect 367098 59256 367154 59265
rect 367098 59191 367154 59200
rect 365720 46300 365772 46306
rect 365720 46242 365772 46248
rect 365720 36712 365772 36718
rect 365720 36654 365772 36660
rect 364432 25628 364484 25634
rect 364432 25570 364484 25576
rect 364340 18692 364392 18698
rect 364340 18634 364392 18640
rect 364616 8220 364668 8226
rect 364616 8162 364668 8168
rect 363604 7608 363656 7614
rect 363604 7550 363656 7556
rect 364628 480 364656 8162
rect 365628 3664 365680 3670
rect 365628 3606 365680 3612
rect 365640 3534 365668 3606
rect 365732 3534 365760 36654
rect 367112 32434 367140 59191
rect 367100 32428 367152 32434
rect 367100 32370 367152 32376
rect 367192 10532 367244 10538
rect 367192 10474 367244 10480
rect 365812 3800 365864 3806
rect 365812 3742 365864 3748
rect 365628 3528 365680 3534
rect 365628 3470 365680 3476
rect 365720 3528 365772 3534
rect 365720 3470 365772 3476
rect 365824 480 365852 3742
rect 367008 3528 367060 3534
rect 367008 3470 367060 3476
rect 367020 480 367048 3470
rect 367204 490 367232 10474
rect 367296 3466 367324 59327
rect 368492 3602 368520 59463
rect 368572 59434 368624 59440
rect 368584 3670 368612 59434
rect 369136 59401 369164 59735
rect 369122 59392 369178 59401
rect 369122 59327 369178 59336
rect 369504 57322 369532 59735
rect 373816 59706 373868 59712
rect 375472 59764 375524 59770
rect 376482 59735 376538 59744
rect 376666 59800 376722 59809
rect 376666 59735 376722 59744
rect 379978 59800 380034 59809
rect 381634 59800 381690 59809
rect 379978 59735 379980 59744
rect 375472 59706 375524 59712
rect 373828 59673 373856 59706
rect 372526 59664 372582 59673
rect 369952 59628 370004 59634
rect 372526 59599 372582 59608
rect 373814 59664 373870 59673
rect 373814 59599 373870 59608
rect 369952 59570 370004 59576
rect 369492 57316 369544 57322
rect 369492 57258 369544 57264
rect 369860 38072 369912 38078
rect 369860 38014 369912 38020
rect 368572 3664 368624 3670
rect 368572 3606 368624 3612
rect 368480 3596 368532 3602
rect 368480 3538 368532 3544
rect 367284 3460 367336 3466
rect 367284 3402 367336 3408
rect 369398 3360 369454 3369
rect 369398 3295 369454 3304
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367204 462 367784 490
rect 369412 480 369440 3295
rect 369872 490 369900 38014
rect 369964 3738 369992 59570
rect 372540 59401 372568 59599
rect 372618 59528 372674 59537
rect 372618 59463 372674 59472
rect 372526 59392 372582 59401
rect 372526 59327 372582 59336
rect 371422 59256 371478 59265
rect 371422 59191 371478 59200
rect 371240 56092 371292 56098
rect 371240 56034 371292 56040
rect 369952 3732 370004 3738
rect 369952 3674 370004 3680
rect 367756 354 367784 462
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 369872 462 370176 490
rect 370148 354 370176 462
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 371252 354 371280 56034
rect 371436 3874 371464 59191
rect 372632 50522 372660 59463
rect 374182 59392 374238 59401
rect 374182 59327 374238 59336
rect 372710 59256 372766 59265
rect 372710 59191 372766 59200
rect 372724 53242 372752 59191
rect 372712 53236 372764 53242
rect 372712 53178 372764 53184
rect 374000 51944 374052 51950
rect 374000 51886 374052 51892
rect 372620 50516 372672 50522
rect 372620 50458 372672 50464
rect 371424 3868 371476 3874
rect 371424 3810 371476 3816
rect 374012 3534 374040 51886
rect 374092 39432 374144 39438
rect 374092 39374 374144 39380
rect 374000 3528 374052 3534
rect 374000 3470 374052 3476
rect 372896 3460 372948 3466
rect 372896 3402 372948 3408
rect 372908 480 372936 3402
rect 374104 480 374132 39374
rect 374196 13122 374224 59327
rect 375484 13190 375512 59706
rect 376496 59401 376524 59735
rect 375654 59392 375710 59401
rect 375654 59327 375710 59336
rect 376482 59392 376538 59401
rect 376482 59327 376538 59336
rect 375668 13258 375696 59327
rect 376680 58750 376708 59735
rect 380032 59735 380034 59744
rect 380992 59764 381044 59770
rect 379980 59706 380032 59712
rect 381634 59735 381690 59744
rect 389454 59800 389510 59809
rect 389454 59735 389510 59744
rect 398838 59800 398894 59809
rect 400678 59800 400734 59809
rect 398894 59758 399156 59786
rect 398838 59735 398894 59744
rect 380992 59706 381044 59712
rect 376942 59664 376998 59673
rect 376942 59599 376998 59608
rect 376758 59528 376814 59537
rect 376758 59463 376814 59472
rect 376668 58744 376720 58750
rect 376668 58686 376720 58692
rect 376772 49162 376800 59463
rect 376760 49156 376812 49162
rect 376760 49098 376812 49104
rect 376760 40724 376812 40730
rect 376760 40666 376812 40672
rect 375656 13252 375708 13258
rect 375656 13194 375708 13200
rect 375472 13184 375524 13190
rect 375472 13126 375524 13132
rect 374184 13116 374236 13122
rect 374184 13058 374236 13064
rect 376024 13116 376076 13122
rect 376024 13058 376076 13064
rect 376036 4010 376064 13058
rect 376772 6914 376800 40666
rect 376956 13326 376984 59599
rect 379702 59528 379758 59537
rect 379702 59463 379758 59472
rect 378230 59392 378286 59401
rect 378230 59327 378286 59336
rect 378140 45076 378192 45082
rect 378140 45018 378192 45024
rect 378152 16574 378180 45018
rect 378244 27062 378272 59327
rect 379716 54670 379744 59463
rect 380898 59256 380954 59265
rect 380898 59191 380954 59200
rect 379704 54664 379756 54670
rect 379704 54606 379756 54612
rect 380912 31210 380940 59191
rect 381004 43518 381032 59706
rect 381648 59265 381676 59735
rect 383106 59664 383162 59673
rect 383106 59599 383162 59608
rect 384118 59664 384174 59673
rect 387430 59664 387486 59673
rect 384118 59599 384120 59608
rect 383120 59401 383148 59599
rect 384172 59599 384174 59608
rect 385408 59628 385460 59634
rect 384120 59570 384172 59576
rect 387430 59599 387486 59608
rect 385408 59570 385460 59576
rect 383934 59528 383990 59537
rect 383934 59463 383990 59472
rect 382370 59392 382426 59401
rect 382370 59327 382426 59336
rect 383106 59392 383162 59401
rect 383106 59327 383162 59336
rect 381634 59256 381690 59265
rect 381634 59191 381690 59200
rect 380992 43512 381044 43518
rect 380992 43454 381044 43460
rect 380900 31204 380952 31210
rect 380900 31146 380952 31152
rect 378232 27056 378284 27062
rect 378232 26998 378284 27004
rect 382280 22976 382332 22982
rect 382280 22918 382332 22924
rect 380900 18760 380952 18766
rect 380900 18702 380952 18708
rect 380912 16574 380940 18702
rect 382292 16574 382320 22918
rect 382384 17406 382412 59327
rect 383750 59256 383806 59265
rect 383750 59191 383806 59200
rect 383764 47734 383792 59191
rect 383752 47728 383804 47734
rect 383752 47670 383804 47676
rect 383948 33930 383976 59463
rect 385222 59256 385278 59265
rect 385222 59191 385278 59200
rect 383936 33924 383988 33930
rect 383936 33866 383988 33872
rect 385040 24336 385092 24342
rect 385040 24278 385092 24284
rect 383660 20052 383712 20058
rect 383660 19994 383712 20000
rect 382372 17400 382424 17406
rect 382372 17342 382424 17348
rect 383672 16574 383700 19994
rect 378152 16546 378456 16574
rect 380912 16546 381216 16574
rect 382292 16546 382412 16574
rect 383672 16546 384344 16574
rect 376944 13320 376996 13326
rect 376944 13262 376996 13268
rect 376772 6886 377720 6914
rect 376024 4004 376076 4010
rect 376024 3946 376076 3952
rect 375288 3528 375340 3534
rect 375288 3470 375340 3476
rect 376484 3528 376536 3534
rect 376484 3470 376536 3476
rect 375300 480 375328 3470
rect 376496 480 376524 3470
rect 377692 480 377720 6886
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 379980 3596 380032 3602
rect 379980 3538 380032 3544
rect 379992 480 380020 3538
rect 381188 480 381216 16546
rect 382384 480 382412 16546
rect 383568 3664 383620 3670
rect 383568 3606 383620 3612
rect 383580 480 383608 3606
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 378846 -960 378958 326
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 16546
rect 385052 6914 385080 24278
rect 385236 14482 385264 59191
rect 385420 14550 385448 59570
rect 385774 59528 385830 59537
rect 385774 59463 385776 59472
rect 385828 59463 385830 59472
rect 385776 59434 385828 59440
rect 387444 59401 387472 59599
rect 387982 59528 388038 59537
rect 387982 59463 388038 59472
rect 388168 59492 388220 59498
rect 386418 59392 386474 59401
rect 386418 59327 386474 59336
rect 387430 59392 387486 59401
rect 387430 59327 387486 59336
rect 386432 14618 386460 59327
rect 387800 46368 387852 46374
rect 387800 46310 387852 46316
rect 386420 14612 386472 14618
rect 386420 14554 386472 14560
rect 385408 14544 385460 14550
rect 385408 14486 385460 14492
rect 385224 14476 385276 14482
rect 385224 14418 385276 14424
rect 385052 6886 386000 6914
rect 385972 480 386000 6886
rect 387156 3732 387208 3738
rect 387156 3674 387208 3680
rect 387168 480 387196 3674
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 387812 354 387840 46310
rect 387996 14754 388024 59463
rect 388168 59434 388220 59440
rect 387984 14748 388036 14754
rect 387984 14690 388036 14696
rect 388180 14686 388208 59434
rect 389362 59256 389418 59265
rect 389362 59191 389418 59200
rect 389180 40928 389232 40934
rect 389180 40870 389232 40876
rect 388168 14680 388220 14686
rect 388168 14622 388220 14628
rect 389192 6914 389220 40870
rect 389376 14822 389404 59191
rect 389468 55962 389496 59735
rect 393318 59664 393374 59673
rect 393318 59599 393320 59608
rect 393372 59599 393374 59608
rect 394792 59628 394844 59634
rect 393320 59570 393372 59576
rect 394792 59570 394844 59576
rect 390558 59528 390614 59537
rect 390558 59463 390614 59472
rect 393318 59528 393374 59537
rect 394698 59528 394754 59537
rect 393374 59486 393452 59514
rect 393318 59463 393374 59472
rect 389546 59392 389602 59401
rect 389546 59327 389602 59336
rect 389456 55956 389508 55962
rect 389456 55898 389508 55904
rect 389560 14890 389588 59327
rect 390572 40866 390600 59463
rect 392122 59256 392178 59265
rect 392122 59191 392178 59200
rect 390560 40860 390612 40866
rect 390560 40802 390612 40808
rect 391940 29844 391992 29850
rect 391940 29786 391992 29792
rect 390560 21480 390612 21486
rect 390560 21422 390612 21428
rect 389548 14884 389600 14890
rect 389548 14826 389600 14832
rect 389364 14816 389416 14822
rect 389364 14758 389416 14764
rect 389192 6886 389496 6914
rect 389468 480 389496 6886
rect 390572 3398 390600 21422
rect 391952 6914 391980 29786
rect 392136 14958 392164 59191
rect 393424 42294 393452 59486
rect 394698 59463 394754 59472
rect 393594 59256 393650 59265
rect 393594 59191 393650 59200
rect 393412 42288 393464 42294
rect 393412 42230 393464 42236
rect 393608 15026 393636 59191
rect 394712 57458 394740 59463
rect 394700 57452 394752 57458
rect 394700 57394 394752 57400
rect 394804 45554 394832 59570
rect 397550 59528 397606 59537
rect 397550 59463 397606 59472
rect 396354 59392 396410 59401
rect 396354 59327 396410 59336
rect 396170 59256 396226 59265
rect 396170 59191 396226 59200
rect 394712 45526 394832 45554
rect 394712 35426 394740 45526
rect 396184 36786 396212 59191
rect 396172 36780 396224 36786
rect 396172 36722 396224 36728
rect 394700 35420 394752 35426
rect 394700 35362 394752 35368
rect 396080 32632 396132 32638
rect 396080 32574 396132 32580
rect 393596 15020 393648 15026
rect 393596 14962 393648 14968
rect 392124 14952 392176 14958
rect 392124 14894 392176 14900
rect 395344 9240 395396 9246
rect 395344 9182 395396 9188
rect 391952 6886 392624 6914
rect 390652 3868 390704 3874
rect 390652 3810 390704 3816
rect 390560 3392 390612 3398
rect 390560 3334 390612 3340
rect 390664 480 390692 3810
rect 391848 3392 391900 3398
rect 391848 3334 391900 3340
rect 391860 480 391888 3334
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 6886
rect 394240 3936 394292 3942
rect 394240 3878 394292 3884
rect 394252 480 394280 3878
rect 395356 480 395384 9182
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 32574
rect 396368 29782 396396 59327
rect 397564 38146 397592 59463
rect 399128 59401 399156 59758
rect 400954 59800 401010 59809
rect 400734 59758 400954 59786
rect 400678 59735 400734 59744
rect 400954 59735 401010 59744
rect 401782 59800 401838 59809
rect 401782 59735 401838 59744
rect 406566 59800 406622 59809
rect 409050 59800 409106 59809
rect 406566 59735 406568 59744
rect 400310 59528 400366 59537
rect 400310 59463 400366 59472
rect 401506 59528 401562 59537
rect 401506 59463 401562 59472
rect 398930 59392 398986 59401
rect 398930 59327 398986 59336
rect 399114 59392 399170 59401
rect 399114 59327 399170 59336
rect 398840 56024 398892 56030
rect 398840 55966 398892 55972
rect 397552 38140 397604 38146
rect 397552 38082 397604 38088
rect 396356 29776 396408 29782
rect 396356 29718 396408 29724
rect 397736 4004 397788 4010
rect 397736 3946 397788 3952
rect 397748 480 397776 3946
rect 398852 3398 398880 55966
rect 398944 21622 398972 59327
rect 398932 21616 398984 21622
rect 398932 21558 398984 21564
rect 400324 15910 400352 59463
rect 400494 59392 400550 59401
rect 400494 59327 400550 59336
rect 400312 15904 400364 15910
rect 400312 15846 400364 15852
rect 400508 10470 400536 59327
rect 401520 58886 401548 59463
rect 401598 59256 401654 59265
rect 401598 59191 401654 59200
rect 401508 58880 401560 58886
rect 401508 58822 401560 58828
rect 401612 51882 401640 59191
rect 401600 51876 401652 51882
rect 401600 51818 401652 51824
rect 401600 25696 401652 25702
rect 401600 25638 401652 25644
rect 401612 16574 401640 25638
rect 401796 20194 401824 59735
rect 406620 59735 406622 59744
rect 408500 59764 408552 59770
rect 406568 59706 406620 59712
rect 412822 59800 412878 59809
rect 409050 59735 409052 59744
rect 408500 59706 408552 59712
rect 409104 59735 409106 59744
rect 410156 59764 410208 59770
rect 409052 59706 409104 59712
rect 412822 59735 412878 59744
rect 417606 59800 417662 59809
rect 422390 59800 422392 59809
rect 424140 59832 424192 59838
rect 422444 59800 422446 59809
rect 417606 59735 417608 59744
rect 410156 59706 410208 59712
rect 405738 59528 405794 59537
rect 405738 59463 405794 59472
rect 402978 59256 403034 59265
rect 402978 59191 403034 59200
rect 404542 59256 404598 59265
rect 404542 59191 404598 59200
rect 401784 20188 401836 20194
rect 401784 20130 401836 20136
rect 401612 16546 402560 16574
rect 400496 10464 400548 10470
rect 400496 10406 400548 10412
rect 398932 9172 398984 9178
rect 398932 9114 398984 9120
rect 398840 3392 398892 3398
rect 398840 3334 398892 3340
rect 398944 480 398972 9114
rect 401324 4072 401376 4078
rect 401324 4014 401376 4020
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 400140 480 400168 3334
rect 401336 480 401364 4014
rect 402532 480 402560 16546
rect 402992 15978 403020 59191
rect 403072 18828 403124 18834
rect 403072 18770 403124 18776
rect 403084 16574 403112 18770
rect 403084 16546 403664 16574
rect 402980 15972 403032 15978
rect 402980 15914 403032 15920
rect 403636 480 403664 16546
rect 404556 16046 404584 59191
rect 405752 28490 405780 59463
rect 405830 59392 405886 59401
rect 405830 59327 405886 59336
rect 407210 59392 407266 59401
rect 407210 59327 407266 59336
rect 405844 39506 405872 59327
rect 407120 51808 407172 51814
rect 407120 51750 407172 51756
rect 405832 39500 405884 39506
rect 405832 39442 405884 39448
rect 405740 28484 405792 28490
rect 405740 28426 405792 28432
rect 404544 16040 404596 16046
rect 404544 15982 404596 15988
rect 406016 9104 406068 9110
rect 406016 9046 406068 9052
rect 404820 4140 404872 4146
rect 404820 4082 404872 4088
rect 404832 480 404860 4082
rect 406028 480 406056 9046
rect 407132 6914 407160 51750
rect 407224 16114 407252 59327
rect 408512 53310 408540 59706
rect 408774 59528 408830 59537
rect 408774 59463 408830 59472
rect 408500 53304 408552 53310
rect 408500 53246 408552 53252
rect 408788 43654 408816 59463
rect 409970 59256 410026 59265
rect 409970 59191 410026 59200
rect 409984 50590 410012 59191
rect 409972 50584 410024 50590
rect 409972 50526 410024 50532
rect 408776 43648 408828 43654
rect 408776 43590 408828 43596
rect 408500 26988 408552 26994
rect 408500 26930 408552 26936
rect 408512 16574 408540 26930
rect 410168 22914 410196 59706
rect 411534 59664 411590 59673
rect 411534 59599 411590 59608
rect 412362 59664 412418 59673
rect 412730 59664 412786 59673
rect 412418 59622 412730 59650
rect 412362 59599 412418 59608
rect 412730 59599 412786 59608
rect 411548 59401 411576 59599
rect 412362 59528 412418 59537
rect 412418 59486 412772 59514
rect 412362 59463 412418 59472
rect 411534 59392 411590 59401
rect 411534 59327 411590 59336
rect 411258 59256 411314 59265
rect 411258 59191 411314 59200
rect 411272 33998 411300 59191
rect 412744 49230 412772 59486
rect 412836 54738 412864 59735
rect 417660 59735 417662 59744
rect 419632 59764 419684 59770
rect 417608 59706 417660 59712
rect 419632 59706 419684 59712
rect 422116 59764 422168 59770
rect 424140 59774 424192 59780
rect 425702 59800 425758 59809
rect 422390 59735 422446 59744
rect 423956 59764 424008 59770
rect 422116 59706 422168 59712
rect 423956 59706 424008 59712
rect 414110 59664 414166 59673
rect 417606 59664 417662 59673
rect 414166 59622 414336 59650
rect 414110 59599 414166 59608
rect 414110 59528 414166 59537
rect 414110 59463 414166 59472
rect 412914 59392 412970 59401
rect 412914 59327 412970 59336
rect 412824 54732 412876 54738
rect 412824 54674 412876 54680
rect 412732 49224 412784 49230
rect 412732 49166 412784 49172
rect 411260 33992 411312 33998
rect 411260 33934 411312 33940
rect 410156 22908 410208 22914
rect 410156 22850 410208 22856
rect 408512 16546 409184 16574
rect 407212 16108 407264 16114
rect 407212 16050 407264 16056
rect 407132 6886 407252 6914
rect 407224 480 407252 6886
rect 408408 3392 408460 3398
rect 408408 3334 408460 3340
rect 408420 480 408448 3334
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 412928 16182 412956 59327
rect 414124 44946 414152 59463
rect 414112 44940 414164 44946
rect 414112 44882 414164 44888
rect 414308 31278 414336 59622
rect 417606 59599 417662 59608
rect 417054 59392 417110 59401
rect 417054 59327 417110 59336
rect 416870 59256 416926 59265
rect 416870 59191 416926 59200
rect 414296 31272 414348 31278
rect 414296 31214 414348 31220
rect 416884 29714 416912 59191
rect 416872 29708 416924 29714
rect 416872 29650 416924 29656
rect 417068 18902 417096 59327
rect 417620 58546 417648 59599
rect 418250 59528 418306 59537
rect 418250 59463 418306 59472
rect 419078 59528 419134 59537
rect 419078 59463 419080 59472
rect 417608 58540 417660 58546
rect 417608 58482 417660 58488
rect 417056 18896 417108 18902
rect 417056 18838 417108 18844
rect 412916 16176 412968 16182
rect 412916 16118 412968 16124
rect 418264 13122 418292 59463
rect 419132 59463 419134 59472
rect 419080 59434 419132 59440
rect 418436 58540 418488 58546
rect 418436 58482 418488 58488
rect 418252 13116 418304 13122
rect 418252 13058 418304 13064
rect 410800 12300 410852 12306
rect 410800 12242 410852 12248
rect 410812 480 410840 12242
rect 414296 12232 414348 12238
rect 414296 12174 414348 12180
rect 413100 9036 413152 9042
rect 413100 8978 413152 8984
rect 411904 3324 411956 3330
rect 411904 3266 411956 3272
rect 411916 480 411944 3266
rect 413112 480 413140 8978
rect 414308 480 414336 12174
rect 417424 12164 417476 12170
rect 417424 12106 417476 12112
rect 416688 8968 416740 8974
rect 416688 8910 416740 8916
rect 415492 3256 415544 3262
rect 415492 3198 415544 3204
rect 415504 480 415532 3198
rect 416700 480 416728 8910
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 12106
rect 418448 3806 418476 58482
rect 419540 32496 419592 32502
rect 419540 32438 419592 32444
rect 418436 3800 418488 3806
rect 418436 3742 418488 3748
rect 419552 3482 419580 32438
rect 419644 3641 419672 59706
rect 422128 59673 422156 59706
rect 420734 59664 420790 59673
rect 420734 59599 420790 59608
rect 422114 59664 422170 59673
rect 422114 59599 422170 59608
rect 422298 59664 422354 59673
rect 422298 59599 422354 59608
rect 420748 59401 420776 59599
rect 421102 59528 421158 59537
rect 421102 59463 421158 59472
rect 421288 59492 421340 59498
rect 420734 59392 420790 59401
rect 420734 59327 420790 59336
rect 420920 39568 420972 39574
rect 420920 39510 420972 39516
rect 419630 3632 419686 3641
rect 419630 3567 419686 3576
rect 419552 3454 420224 3482
rect 418988 3188 419040 3194
rect 418988 3130 419040 3136
rect 419000 480 419028 3130
rect 420196 480 420224 3454
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 417854 -960 417966 326
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 420932 354 420960 39510
rect 421116 3534 421144 59463
rect 421288 59434 421340 59440
rect 421104 3528 421156 3534
rect 421104 3470 421156 3476
rect 421300 3466 421328 59434
rect 422312 3602 422340 59599
rect 423680 47660 423732 47666
rect 423680 47602 423732 47608
rect 422300 3596 422352 3602
rect 422300 3538 422352 3544
rect 421288 3460 421340 3466
rect 421288 3402 421340 3408
rect 422576 3460 422628 3466
rect 422576 3402 422628 3408
rect 422588 480 422616 3402
rect 423692 3346 423720 47602
rect 423772 12096 423824 12102
rect 423772 12038 423824 12044
rect 423784 3534 423812 12038
rect 423968 3670 423996 59706
rect 424152 3738 424180 59774
rect 428094 59800 428150 59809
rect 425702 59735 425704 59744
rect 425756 59735 425758 59744
rect 428004 59764 428056 59770
rect 425704 59706 425756 59712
rect 428094 59735 428150 59744
rect 429014 59800 429070 59809
rect 429014 59735 429070 59744
rect 429842 59800 429898 59809
rect 435822 59800 435878 59809
rect 429842 59735 429844 59744
rect 428004 59706 428056 59712
rect 425058 59528 425114 59537
rect 425058 59463 425114 59472
rect 425072 3942 425100 59463
rect 425150 59392 425206 59401
rect 425150 59327 425206 59336
rect 426530 59392 426586 59401
rect 426530 59327 426586 59336
rect 425060 3936 425112 3942
rect 425060 3878 425112 3884
rect 425164 3874 425192 59327
rect 426440 28416 426492 28422
rect 426440 28358 426492 28364
rect 425152 3868 425204 3874
rect 425152 3810 425204 3816
rect 424140 3732 424192 3738
rect 424140 3674 424192 3680
rect 423956 3664 424008 3670
rect 423956 3606 424008 3612
rect 423772 3528 423824 3534
rect 423772 3470 423824 3476
rect 424968 3528 425020 3534
rect 424968 3470 425020 3476
rect 423692 3318 423812 3346
rect 423784 480 423812 3318
rect 424980 480 425008 3470
rect 426164 3460 426216 3466
rect 426164 3402 426216 3408
rect 426176 480 426204 3402
rect 426452 490 426480 28358
rect 426544 4010 426572 59327
rect 427912 12028 427964 12034
rect 427912 11970 427964 11976
rect 426532 4004 426584 4010
rect 426532 3946 426584 3952
rect 427924 3482 427952 11970
rect 428016 4078 428044 59706
rect 428108 59401 428136 59735
rect 429028 59537 429056 59735
rect 429896 59735 429898 59744
rect 432328 59764 432380 59770
rect 429844 59706 429896 59712
rect 435822 59735 435824 59744
rect 432328 59706 432380 59712
rect 435876 59735 435878 59744
rect 438214 59800 438270 59809
rect 438766 59800 438822 59809
rect 438214 59735 438270 59744
rect 438308 59764 438360 59770
rect 435824 59706 435876 59712
rect 429198 59664 429254 59673
rect 429198 59599 429254 59608
rect 430578 59664 430634 59673
rect 430578 59599 430634 59608
rect 431776 59628 431828 59634
rect 428186 59528 428242 59537
rect 428186 59463 428242 59472
rect 429014 59528 429070 59537
rect 429014 59463 429070 59472
rect 428094 59392 428150 59401
rect 428094 59327 428150 59336
rect 428200 4146 428228 59463
rect 428188 4140 428240 4146
rect 428188 4082 428240 4088
rect 428004 4072 428056 4078
rect 428004 4014 428056 4020
rect 427924 3454 428504 3482
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 426452 462 426848 490
rect 428476 480 428504 3454
rect 429212 3398 429240 59599
rect 430592 59401 430620 59599
rect 431776 59570 431828 59576
rect 431788 59537 431816 59570
rect 430670 59528 430726 59537
rect 430670 59463 430726 59472
rect 431774 59528 431830 59537
rect 431774 59463 431830 59472
rect 429290 59392 429346 59401
rect 429290 59327 429346 59336
rect 430578 59392 430634 59401
rect 430578 59327 430634 59336
rect 429200 3392 429252 3398
rect 429200 3334 429252 3340
rect 429304 3330 429332 59327
rect 430580 43444 430632 43450
rect 430580 43386 430632 43392
rect 429660 4004 429712 4010
rect 429660 3946 429712 3952
rect 429292 3324 429344 3330
rect 429292 3266 429344 3272
rect 429672 480 429700 3946
rect 430592 3074 430620 43386
rect 430684 3262 430712 59463
rect 432142 59392 432198 59401
rect 432142 59327 432198 59336
rect 432052 11960 432104 11966
rect 432052 11902 432104 11908
rect 430672 3256 430724 3262
rect 430672 3198 430724 3204
rect 430592 3046 430896 3074
rect 430868 480 430896 3046
rect 432064 480 432092 11902
rect 432156 3534 432184 59327
rect 432144 3528 432196 3534
rect 432144 3470 432196 3476
rect 432340 3194 432368 59706
rect 438228 59702 438256 59735
rect 438766 59735 438822 59744
rect 440698 59800 440754 59809
rect 440698 59735 440754 59744
rect 441250 59800 441306 59809
rect 441250 59735 441306 59744
rect 442354 59800 442410 59809
rect 445666 59800 445722 59809
rect 442354 59735 442356 59744
rect 438308 59706 438360 59712
rect 438216 59696 438268 59702
rect 433982 59664 434038 59673
rect 433708 59628 433760 59634
rect 438216 59638 438268 59644
rect 433982 59599 434038 59608
rect 433708 59570 433760 59576
rect 433522 59392 433578 59401
rect 433522 59327 433578 59336
rect 433340 31136 433392 31142
rect 433340 31078 433392 31084
rect 433352 16574 433380 31078
rect 433352 16546 433472 16574
rect 433248 3324 433300 3330
rect 433248 3266 433300 3272
rect 432328 3188 432380 3194
rect 432328 3130 432380 3136
rect 433260 480 433288 3266
rect 433444 490 433472 16546
rect 433536 4010 433564 59327
rect 433524 4004 433576 4010
rect 433524 3946 433576 3952
rect 433720 3466 433748 59570
rect 433996 59401 434024 59599
rect 434810 59528 434866 59537
rect 434810 59463 434866 59472
rect 438122 59528 438178 59537
rect 438122 59463 438178 59472
rect 433982 59392 434038 59401
rect 433982 59327 434038 59336
rect 434720 11892 434772 11898
rect 434720 11834 434772 11840
rect 433708 3460 433760 3466
rect 433708 3402 433760 3408
rect 434732 490 434760 11834
rect 434824 3330 434852 59463
rect 436742 59392 436798 59401
rect 436742 59327 436798 59336
rect 436098 59256 436154 59265
rect 436098 59191 436154 59200
rect 436112 6914 436140 59191
rect 436756 16574 436784 59327
rect 437480 33788 437532 33794
rect 437480 33730 437532 33736
rect 436756 16546 436876 16574
rect 436112 6886 436784 6914
rect 434812 3324 434864 3330
rect 434812 3266 434864 3272
rect 426820 354 426848 462
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433444 462 434024 490
rect 433996 354 434024 462
rect 434414 354 434526 480
rect 434732 462 435128 490
rect 436756 480 436784 6886
rect 436848 3398 436876 16546
rect 436836 3392 436888 3398
rect 436836 3334 436888 3340
rect 433996 326 434526 354
rect 435100 354 435128 462
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 33730
rect 438136 3942 438164 59463
rect 438124 3936 438176 3942
rect 438124 3878 438176 3884
rect 438320 3330 438348 59706
rect 438780 59401 438808 59735
rect 440712 59537 440740 59735
rect 440884 59696 440936 59702
rect 440884 59638 440936 59644
rect 439502 59528 439558 59537
rect 439502 59463 439558 59472
rect 440698 59528 440754 59537
rect 440698 59463 440754 59472
rect 438766 59392 438822 59401
rect 438766 59327 438822 59336
rect 439136 11824 439188 11830
rect 439136 11766 439188 11772
rect 438308 3324 438360 3330
rect 438308 3266 438360 3272
rect 439148 480 439176 11766
rect 439516 3874 439544 59463
rect 440332 49088 440384 49094
rect 440332 49030 440384 49036
rect 439504 3868 439556 3874
rect 439504 3810 439556 3816
rect 440344 3534 440372 49030
rect 440896 3806 440924 59638
rect 441264 59401 441292 59735
rect 442408 59735 442410 59744
rect 445208 59764 445260 59770
rect 442356 59706 442408 59712
rect 450542 59800 450598 59809
rect 445666 59735 445668 59744
rect 445208 59706 445260 59712
rect 445720 59735 445722 59744
rect 447784 59764 447836 59770
rect 445668 59706 445720 59712
rect 450542 59735 450598 59744
rect 454774 59800 454830 59809
rect 454774 59735 454830 59744
rect 455602 59800 455658 59809
rect 455602 59735 455658 59744
rect 456522 59800 456578 59809
rect 461490 59800 461546 59809
rect 456522 59735 456524 59744
rect 447784 59706 447836 59712
rect 442262 59664 442318 59673
rect 442262 59599 442318 59608
rect 444010 59664 444066 59673
rect 444010 59599 444066 59608
rect 441066 59392 441122 59401
rect 441066 59327 441122 59336
rect 441250 59392 441306 59401
rect 441250 59327 441306 59336
rect 440884 3800 440936 3806
rect 440884 3742 440936 3748
rect 441080 3738 441108 59327
rect 442172 11756 442224 11762
rect 442172 11698 442224 11704
rect 441068 3732 441120 3738
rect 441068 3674 441120 3680
rect 440332 3528 440384 3534
rect 440332 3470 440384 3476
rect 441528 3528 441580 3534
rect 441528 3470 441580 3476
rect 442184 3482 442212 11698
rect 442276 3670 442304 59599
rect 442354 59528 442410 59537
rect 442410 59486 442488 59514
rect 442354 59463 442410 59472
rect 442264 3664 442316 3670
rect 442264 3606 442316 3612
rect 442460 3602 442488 59486
rect 444024 59401 444052 59599
rect 445022 59528 445078 59537
rect 445022 59463 445078 59472
rect 443642 59392 443698 59401
rect 443642 59327 443698 59336
rect 444010 59392 444066 59401
rect 444010 59327 444066 59336
rect 442448 3596 442500 3602
rect 442448 3538 442500 3544
rect 440332 3392 440384 3398
rect 440332 3334 440384 3340
rect 440344 480 440372 3334
rect 441540 480 441568 3470
rect 442184 3454 442672 3482
rect 443656 3466 443684 59327
rect 444380 35216 444432 35222
rect 444380 35158 444432 35164
rect 444392 6914 444420 35158
rect 445036 16574 445064 59463
rect 445036 16546 445156 16574
rect 444392 6886 445064 6914
rect 442644 480 442672 3454
rect 443644 3460 443696 3466
rect 443644 3402 443696 3408
rect 443828 3324 443880 3330
rect 443828 3266 443880 3272
rect 443840 480 443868 3266
rect 445036 480 445064 6886
rect 445128 3262 445156 16546
rect 445220 3602 445248 59706
rect 445666 59664 445722 59673
rect 445722 59622 446628 59650
rect 445666 59599 445722 59608
rect 446404 59560 446456 59566
rect 446402 59528 446404 59537
rect 446456 59528 446458 59537
rect 446402 59463 446458 59472
rect 446402 59392 446458 59401
rect 446402 59327 446458 59336
rect 445760 22840 445812 22846
rect 445760 22782 445812 22788
rect 445208 3596 445260 3602
rect 445208 3538 445260 3544
rect 445116 3256 445168 3262
rect 445116 3198 445168 3204
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 354 445800 22782
rect 446416 3330 446444 59327
rect 446600 15978 446628 59622
rect 446588 15972 446640 15978
rect 446588 15914 446640 15920
rect 447796 11762 447824 59706
rect 448520 59560 448572 59566
rect 448150 59528 448206 59537
rect 448520 59502 448572 59508
rect 450450 59528 450506 59537
rect 448150 59463 448152 59472
rect 448204 59463 448206 59472
rect 448152 59434 448204 59440
rect 448532 55962 448560 59502
rect 450450 59463 450506 59472
rect 449162 59392 449218 59401
rect 449162 59327 449218 59336
rect 448520 55956 448572 55962
rect 448520 55898 448572 55904
rect 448520 50448 448572 50454
rect 448520 50390 448572 50396
rect 447784 11756 447836 11762
rect 447784 11698 447836 11704
rect 447416 3936 447468 3942
rect 447416 3878 447468 3884
rect 446404 3324 446456 3330
rect 446404 3266 446456 3272
rect 447428 480 447456 3878
rect 448532 2774 448560 50390
rect 448612 45008 448664 45014
rect 448612 44950 448664 44956
rect 448624 7546 448652 44950
rect 449176 39438 449204 59327
rect 450464 55214 450492 59463
rect 450556 59401 450584 59735
rect 454788 59702 454816 59735
rect 454776 59696 454828 59702
rect 450634 59664 450690 59673
rect 454776 59638 454828 59644
rect 450634 59599 450636 59608
rect 450688 59599 450690 59608
rect 451924 59628 451976 59634
rect 450636 59570 450688 59576
rect 451924 59570 451976 59576
rect 450728 59492 450780 59498
rect 450728 59434 450780 59440
rect 450542 59392 450598 59401
rect 450542 59327 450598 59336
rect 450464 55186 450584 55214
rect 449164 39432 449216 39438
rect 449164 39374 449216 39380
rect 450556 8226 450584 55186
rect 450740 14482 450768 59434
rect 451278 59392 451334 59401
rect 451278 59327 451280 59336
rect 451332 59327 451334 59336
rect 451280 59298 451332 59304
rect 451936 53174 451964 59570
rect 452290 59528 452346 59537
rect 452290 59463 452292 59472
rect 452344 59463 452346 59472
rect 454682 59528 454738 59537
rect 454682 59463 454738 59472
rect 454868 59492 454920 59498
rect 452292 59434 452344 59440
rect 453302 59392 453358 59401
rect 453302 59327 453358 59336
rect 453488 59356 453540 59362
rect 451280 53168 451332 53174
rect 451280 53110 451332 53116
rect 451924 53168 451976 53174
rect 451924 53110 451976 53116
rect 451292 16574 451320 53110
rect 452660 20120 452712 20126
rect 452660 20062 452712 20068
rect 451292 16546 451688 16574
rect 450728 14476 450780 14482
rect 450728 14418 450780 14424
rect 450544 8220 450596 8226
rect 450544 8162 450596 8168
rect 448612 7540 448664 7546
rect 448612 7482 448664 7488
rect 449808 7540 449860 7546
rect 449808 7482 449860 7488
rect 449164 3528 449216 3534
rect 449164 3470 449216 3476
rect 449176 3398 449204 3470
rect 449164 3392 449216 3398
rect 449164 3334 449216 3340
rect 448532 2746 448652 2774
rect 448624 480 448652 2746
rect 449820 480 449848 7482
rect 450912 3868 450964 3874
rect 450912 3810 450964 3816
rect 450924 480 450952 3810
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 452672 2774 452700 20062
rect 453316 9178 453344 59327
rect 453488 59298 453540 59304
rect 453304 9172 453356 9178
rect 453304 9114 453356 9120
rect 453500 9110 453528 59298
rect 453488 9104 453540 9110
rect 453488 9046 453540 9052
rect 454696 9042 454724 59463
rect 454868 59434 454920 59440
rect 454880 13122 454908 59434
rect 455616 59401 455644 59735
rect 456576 59735 456578 59744
rect 458824 59764 458876 59770
rect 456524 59706 456576 59712
rect 467930 59800 467986 59809
rect 461490 59735 461492 59744
rect 458824 59706 458876 59712
rect 461544 59735 461546 59744
rect 462964 59764 463016 59770
rect 461492 59706 461544 59712
rect 467930 59735 467986 59744
rect 462964 59706 463016 59712
rect 457444 59696 457496 59702
rect 456062 59664 456118 59673
rect 457444 59638 457496 59644
rect 458178 59664 458234 59673
rect 456062 59599 456118 59608
rect 455602 59392 455658 59401
rect 455602 59327 455658 59336
rect 456076 40730 456104 59599
rect 456064 40724 456116 40730
rect 456064 40666 456116 40672
rect 455420 36576 455472 36582
rect 455420 36518 455472 36524
rect 455432 16574 455460 36518
rect 456892 21548 456944 21554
rect 456892 21490 456944 21496
rect 455432 16546 455736 16574
rect 454868 13116 454920 13122
rect 454868 13058 454920 13064
rect 454684 9036 454736 9042
rect 454684 8978 454736 8984
rect 454500 3800 454552 3806
rect 454500 3742 454552 3748
rect 452672 2746 453344 2774
rect 453316 480 453344 2746
rect 454512 480 454540 3742
rect 455708 480 455736 16546
rect 456904 480 456932 21490
rect 457456 8974 457484 59638
rect 458178 59599 458180 59608
rect 458232 59599 458234 59608
rect 458180 59570 458232 59576
rect 457626 59392 457682 59401
rect 457626 59327 457682 59336
rect 457640 32434 457668 59327
rect 457628 32428 457680 32434
rect 457628 32370 457680 32376
rect 458836 10402 458864 59706
rect 458914 59664 458970 59673
rect 460478 59664 460534 59673
rect 458914 59599 458970 59608
rect 460204 59628 460256 59634
rect 458928 59401 458956 59599
rect 460478 59599 460534 59608
rect 460204 59570 460256 59576
rect 459006 59528 459062 59537
rect 459006 59463 459062 59472
rect 458914 59392 458970 59401
rect 458914 59327 458970 59336
rect 459020 15910 459048 59463
rect 459560 46436 459612 46442
rect 459560 46378 459612 46384
rect 459572 16574 459600 46378
rect 460216 18698 460244 59570
rect 460492 59401 460520 59599
rect 461490 59528 461546 59537
rect 461546 59486 461624 59514
rect 461490 59463 461546 59472
rect 460478 59392 460534 59401
rect 460478 59327 460534 59336
rect 461490 59392 461546 59401
rect 461490 59327 461492 59336
rect 461544 59327 461546 59336
rect 461492 59298 461544 59304
rect 460204 18692 460256 18698
rect 460204 18634 460256 18640
rect 461596 16574 461624 59486
rect 461766 59256 461822 59265
rect 461766 59191 461822 59200
rect 461780 20058 461808 59191
rect 462320 42084 462372 42090
rect 462320 42026 462372 42032
rect 461768 20052 461820 20058
rect 461768 19994 461820 20000
rect 459572 16546 459968 16574
rect 461596 16546 461716 16574
rect 459008 15904 459060 15910
rect 459008 15846 459060 15852
rect 459192 10464 459244 10470
rect 459192 10406 459244 10412
rect 458824 10396 458876 10402
rect 458824 10338 458876 10344
rect 457444 8968 457496 8974
rect 457444 8910 457496 8916
rect 458088 3732 458140 3738
rect 458088 3674 458140 3680
rect 458100 480 458128 3674
rect 459204 480 459232 10406
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 461584 3664 461636 3670
rect 461584 3606 461636 3612
rect 461596 480 461624 3606
rect 461688 3398 461716 16546
rect 461676 3392 461728 3398
rect 461676 3334 461728 3340
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 42026
rect 462976 4078 463004 59706
rect 464802 59664 464858 59673
rect 464802 59599 464858 59608
rect 467102 59664 467158 59673
rect 467102 59599 467158 59608
rect 463146 59528 463202 59537
rect 463146 59463 463148 59472
rect 463200 59463 463202 59472
rect 463148 59434 463200 59440
rect 464816 59401 464844 59599
rect 465722 59528 465778 59537
rect 465722 59463 465778 59472
rect 465908 59492 465960 59498
rect 464342 59392 464398 59401
rect 463148 59356 463200 59362
rect 464342 59327 464398 59336
rect 464802 59392 464858 59401
rect 464802 59327 464858 59336
rect 463148 59298 463200 59304
rect 463160 4146 463188 59298
rect 463700 24268 463752 24274
rect 463700 24210 463752 24216
rect 463712 16574 463740 24210
rect 463712 16546 464016 16574
rect 463148 4140 463200 4146
rect 463148 4082 463200 4088
rect 462964 4072 463016 4078
rect 462964 4014 463016 4020
rect 463988 480 464016 16546
rect 464356 4010 464384 59327
rect 465172 54596 465224 54602
rect 465172 54538 465224 54544
rect 465184 16574 465212 54538
rect 465184 16546 465672 16574
rect 464344 4004 464396 4010
rect 464344 3946 464396 3952
rect 465172 3528 465224 3534
rect 465172 3470 465224 3476
rect 465184 480 465212 3470
rect 465644 490 465672 16546
rect 465736 3874 465764 59463
rect 465908 59434 465960 59440
rect 465920 3942 465948 59434
rect 466460 25764 466512 25770
rect 466460 25706 466512 25712
rect 466472 16574 466500 25706
rect 466472 16546 467052 16574
rect 465908 3936 465960 3942
rect 465908 3878 465960 3884
rect 465724 3868 465776 3874
rect 465724 3810 465776 3816
rect 467024 3482 467052 16546
rect 467116 3738 467144 59599
rect 467286 59392 467342 59401
rect 467286 59327 467342 59336
rect 467300 3806 467328 59327
rect 467944 55214 467972 59735
rect 472622 59664 472678 59673
rect 472622 59599 472678 59608
rect 471426 59528 471482 59537
rect 471426 59463 471482 59472
rect 471242 59392 471298 59401
rect 471242 59327 471298 59336
rect 470138 59256 470194 59265
rect 470138 59191 470194 59200
rect 467944 55186 468524 55214
rect 467288 3800 467340 3806
rect 467288 3742 467340 3748
rect 467104 3732 467156 3738
rect 467104 3674 467156 3680
rect 468496 3670 468524 55186
rect 469220 37936 469272 37942
rect 469220 37878 469272 37884
rect 469232 16574 469260 37878
rect 469232 16546 469904 16574
rect 468484 3664 468536 3670
rect 468484 3606 468536 3612
rect 467024 3454 467512 3482
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465644 462 465856 490
rect 467484 480 467512 3454
rect 468668 3460 468720 3466
rect 468668 3402 468720 3408
rect 468680 480 468708 3402
rect 469876 480 469904 16546
rect 470152 3534 470180 59191
rect 470600 47796 470652 47802
rect 470600 47738 470652 47744
rect 470140 3528 470192 3534
rect 470140 3470 470192 3476
rect 465828 354 465856 462
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 354 470640 47738
rect 471256 3466 471284 59327
rect 471244 3460 471296 3466
rect 471244 3402 471296 3408
rect 471440 3369 471468 59463
rect 472636 3602 472664 59599
rect 538220 58812 538272 58818
rect 538220 58754 538272 58760
rect 483020 58676 483072 58682
rect 483020 58618 483072 58624
rect 473360 39364 473412 39370
rect 473360 39306 473412 39312
rect 473372 6914 473400 39306
rect 473452 27124 473504 27130
rect 473452 27066 473504 27072
rect 473464 16574 473492 27066
rect 480260 17264 480312 17270
rect 480260 17206 480312 17212
rect 480272 16574 480300 17206
rect 483032 16574 483060 58618
rect 494060 57248 494112 57254
rect 494060 57190 494112 57196
rect 489920 55956 489972 55962
rect 489920 55898 489972 55904
rect 487160 18624 487212 18630
rect 487160 18566 487212 18572
rect 473464 16546 474136 16574
rect 480272 16546 480576 16574
rect 483032 16546 484072 16574
rect 473372 6886 473492 6914
rect 472256 3596 472308 3602
rect 472256 3538 472308 3544
rect 472624 3596 472676 3602
rect 472624 3538 472676 3544
rect 471426 3360 471482 3369
rect 471426 3295 471482 3304
rect 472268 480 472296 3538
rect 473464 480 473492 6886
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 16546
rect 478144 13388 478196 13394
rect 478144 13330 478196 13336
rect 476488 10328 476540 10334
rect 476488 10270 476540 10276
rect 475752 3256 475804 3262
rect 475752 3198 475804 3204
rect 475764 480 475792 3198
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 10270
rect 478156 480 478184 13330
rect 479340 3324 479392 3330
rect 479340 3266 479392 3272
rect 479352 480 479380 3266
rect 480548 480 480576 16546
rect 482376 15972 482428 15978
rect 482376 15914 482428 15920
rect 481732 6656 481784 6662
rect 481732 6598 481784 6604
rect 481744 480 481772 6598
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 354 482416 15914
rect 484044 480 484072 16546
rect 486424 11756 486476 11762
rect 486424 11698 486476 11704
rect 485228 6588 485280 6594
rect 485228 6530 485280 6536
rect 485240 480 485268 6530
rect 486436 480 486464 11698
rect 482806 354 482918 480
rect 482388 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487172 354 487200 18566
rect 488816 6520 488868 6526
rect 488816 6462 488868 6468
rect 488828 480 488856 6462
rect 489932 480 489960 55898
rect 492680 39432 492732 39438
rect 492680 39374 492732 39380
rect 490012 19984 490064 19990
rect 490012 19926 490064 19932
rect 490024 16574 490052 19926
rect 492692 16574 492720 39374
rect 494072 16574 494100 57190
rect 500960 55888 501012 55894
rect 500960 55830 501012 55836
rect 495440 40792 495492 40798
rect 495440 40734 495492 40740
rect 490024 16546 490696 16574
rect 492692 16546 493088 16574
rect 494072 16546 494744 16574
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490668 354 490696 16546
rect 492312 6452 492364 6458
rect 492312 6394 492364 6400
rect 492324 480 492352 6394
rect 491086 354 491198 480
rect 490668 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494716 480 494744 16546
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 40734
rect 498200 32564 498252 32570
rect 498200 32506 498252 32512
rect 497096 14476 497148 14482
rect 497096 14418 497148 14424
rect 497108 480 497136 14418
rect 498212 3330 498240 32506
rect 498292 21412 498344 21418
rect 498292 21354 498344 21360
rect 498200 3324 498252 3330
rect 498200 3266 498252 3272
rect 498304 3210 498332 21354
rect 500972 16574 501000 55830
rect 512000 54528 512052 54534
rect 512000 54470 512052 54476
rect 503720 53168 503772 53174
rect 503720 53110 503772 53116
rect 500972 16546 501368 16574
rect 500592 8220 500644 8226
rect 500592 8162 500644 8168
rect 499028 3324 499080 3330
rect 499028 3266 499080 3272
rect 498212 3182 498332 3210
rect 498212 480 498240 3182
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499040 354 499068 3266
rect 500604 480 500632 8162
rect 499366 354 499478 480
rect 499040 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501340 354 501368 16546
rect 502984 6384 503036 6390
rect 502984 6326 503036 6332
rect 502996 480 503024 6326
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503732 354 503760 53110
rect 507860 24132 507912 24138
rect 507860 24074 507912 24080
rect 505100 22772 505152 22778
rect 505100 22714 505152 22720
rect 505112 16574 505140 22714
rect 507872 16574 507900 24074
rect 505112 16546 505416 16574
rect 507872 16546 508912 16574
rect 505388 480 505416 16546
rect 507676 9172 507728 9178
rect 507676 9114 507728 9120
rect 506480 6316 506532 6322
rect 506480 6258 506532 6264
rect 506492 480 506520 6258
rect 507688 480 507716 9114
rect 508884 480 508912 16546
rect 511264 9104 511316 9110
rect 511264 9046 511316 9052
rect 510068 6248 510120 6254
rect 510068 6190 510120 6196
rect 510080 480 510108 6190
rect 511276 480 511304 9046
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512012 354 512040 54470
rect 514760 53100 514812 53106
rect 514760 53042 514812 53048
rect 513564 6180 513616 6186
rect 513564 6122 513616 6128
rect 513576 480 513604 6122
rect 514772 3330 514800 53042
rect 516140 43580 516192 43586
rect 516140 43522 516192 43528
rect 516152 16574 516180 43522
rect 534080 42152 534132 42158
rect 534080 42094 534132 42100
rect 521660 40724 521712 40730
rect 521660 40666 521712 40672
rect 520280 33856 520332 33862
rect 520280 33798 520332 33804
rect 516152 16546 517192 16574
rect 514852 13116 514904 13122
rect 514852 13058 514904 13064
rect 514760 3324 514812 3330
rect 514760 3266 514812 3272
rect 514864 3210 514892 13058
rect 515588 3324 515640 3330
rect 515588 3266 515640 3272
rect 514772 3182 514892 3210
rect 514772 480 514800 3182
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 512430 -960 512542 326
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515600 354 515628 3266
rect 517164 480 517192 16546
rect 518348 9036 518400 9042
rect 518348 8978 518400 8984
rect 518360 480 518388 8978
rect 519544 5160 519596 5166
rect 519544 5102 519596 5108
rect 519556 480 519584 5102
rect 515926 354 516038 480
rect 515600 326 516038 354
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520292 354 520320 33798
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 40666
rect 531320 36644 531372 36650
rect 531320 36586 531372 36592
rect 527180 35284 527232 35290
rect 527180 35226 527232 35232
rect 523040 25560 523092 25566
rect 523040 25502 523092 25508
rect 523052 480 523080 25502
rect 523132 17332 523184 17338
rect 523132 17274 523184 17280
rect 523144 16574 523172 17274
rect 527192 16574 527220 35226
rect 528560 32428 528612 32434
rect 528560 32370 528612 32376
rect 523144 16546 523816 16574
rect 527192 16546 527864 16574
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523788 354 523816 16546
rect 525432 8968 525484 8974
rect 525432 8910 525484 8916
rect 525444 480 525472 8910
rect 526628 5092 526680 5098
rect 526628 5034 526680 5040
rect 526640 480 526668 5034
rect 527836 480 527864 16546
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528572 354 528600 32370
rect 530124 5024 530176 5030
rect 530124 4966 530176 4972
rect 530136 480 530164 4966
rect 531332 480 531360 36586
rect 534092 16574 534120 42094
rect 534092 16546 534488 16574
rect 532056 10396 532108 10402
rect 532056 10338 532108 10344
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 528990 -960 529102 326
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532068 354 532096 10338
rect 533712 4956 533764 4962
rect 533712 4898 533764 4904
rect 533724 480 533752 4898
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536104 15904 536156 15910
rect 536104 15846 536156 15852
rect 536116 480 536144 15846
rect 537208 4888 537260 4894
rect 537208 4830 537260 4836
rect 537220 480 537248 4830
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 58754
rect 545120 57384 545172 57390
rect 545120 57326 545172 57332
rect 543740 51740 543792 51746
rect 543740 51682 543792 51688
rect 540980 38004 541032 38010
rect 540980 37946 541032 37952
rect 539600 18692 539652 18698
rect 539600 18634 539652 18640
rect 539612 480 539640 18634
rect 540992 16574 541020 37946
rect 542360 20052 542412 20058
rect 542360 19994 542412 20000
rect 542372 16574 542400 19994
rect 543752 16574 543780 51682
rect 545132 16574 545160 57326
rect 547880 50380 547932 50386
rect 547880 50322 547932 50328
rect 540992 16546 542032 16574
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 545132 16546 545528 16574
rect 540796 4820 540848 4826
rect 540796 4762 540848 4768
rect 540808 480 540836 4762
rect 542004 480 542032 16546
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545500 480 545528 16546
rect 546684 3392 546736 3398
rect 546684 3334 546736 3340
rect 546696 480 546724 3334
rect 547892 480 547920 50322
rect 554780 49020 554832 49026
rect 554780 48962 554832 48968
rect 550640 26920 550692 26926
rect 550640 26862 550692 26868
rect 550652 16574 550680 26862
rect 550652 16546 551048 16574
rect 549076 8152 549128 8158
rect 549076 8094 549128 8100
rect 549088 480 549116 8094
rect 550272 4140 550324 4146
rect 550272 4082 550324 4088
rect 550284 480 550312 4082
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 552664 8084 552716 8090
rect 552664 8026 552716 8032
rect 552676 480 552704 8026
rect 553768 4072 553820 4078
rect 553768 4014 553820 4020
rect 553780 480 553808 4014
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 48962
rect 561680 47592 561732 47598
rect 561680 47534 561732 47540
rect 557540 28280 557592 28286
rect 557540 28222 557592 28228
rect 557552 16574 557580 28222
rect 561692 16574 561720 47534
rect 564532 46232 564584 46238
rect 564532 46174 564584 46180
rect 564544 16574 564572 46174
rect 572720 44872 572772 44878
rect 572720 44814 572772 44820
rect 568580 29640 568632 29646
rect 568580 29582 568632 29588
rect 568592 16574 568620 29582
rect 557552 16546 558592 16574
rect 561692 16546 562088 16574
rect 564544 16546 565216 16574
rect 568592 16546 568712 16574
rect 556160 8016 556212 8022
rect 556160 7958 556212 7964
rect 556172 480 556200 7958
rect 557356 4004 557408 4010
rect 557356 3946 557408 3952
rect 557368 480 557396 3946
rect 558564 480 558592 16546
rect 559748 7948 559800 7954
rect 559748 7890 559800 7896
rect 559760 480 559788 7890
rect 560852 3936 560904 3942
rect 560852 3878 560904 3884
rect 560864 480 560892 3878
rect 562060 480 562088 16546
rect 563244 7880 563296 7886
rect 563244 7822 563296 7828
rect 563256 480 563284 7822
rect 564440 3868 564492 3874
rect 564440 3810 564492 3816
rect 564452 480 564480 3810
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565188 354 565216 16546
rect 566832 7812 566884 7818
rect 566832 7754 566884 7760
rect 566844 480 566872 7754
rect 568028 3800 568080 3806
rect 568028 3742 568080 3748
rect 568040 480 568068 3742
rect 565606 354 565718 480
rect 565188 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 568684 354 568712 16546
rect 570328 7744 570380 7750
rect 570328 7686 570380 7692
rect 570340 480 570368 7686
rect 571524 3732 571576 3738
rect 571524 3674 571576 3680
rect 571536 480 571564 3674
rect 572732 480 572760 44814
rect 575480 31068 575532 31074
rect 575480 31010 575532 31016
rect 575492 16574 575520 31010
rect 575492 16546 575888 16574
rect 573916 7676 573968 7682
rect 573916 7618 573968 7624
rect 573928 480 573956 7618
rect 575112 3664 575164 3670
rect 575112 3606 575164 3612
rect 575124 480 575152 3606
rect 569102 354 569214 480
rect 568684 326 569214 354
rect 569102 -960 569214 326
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 575860 354 575888 16546
rect 577412 7608 577464 7614
rect 577412 7550 577464 7556
rect 577424 480 577452 7550
rect 582196 3596 582248 3602
rect 582196 3538 582248 3544
rect 578608 3528 578660 3534
rect 578608 3470 578660 3476
rect 578620 480 578648 3470
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 581012 480 581040 3402
rect 582208 480 582236 3538
rect 583390 3360 583446 3369
rect 583390 3295 583446 3304
rect 583404 480 583432 3295
rect 576278 354 576390 480
rect 575860 326 576390 354
rect 576278 -960 576390 326
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 57610 449248 57666 449304
rect 64234 59764 64290 59800
rect 64234 59744 64236 59764
rect 64236 59744 64288 59764
rect 64288 59744 64290 59764
rect 65338 59744 65394 59800
rect 62670 59628 62726 59664
rect 62670 59608 62672 59628
rect 62672 59608 62724 59628
rect 62724 59608 62726 59628
rect 5262 3304 5318 3360
rect 57978 59472 58034 59528
rect 58622 59336 58678 59392
rect 62762 59336 62818 59392
rect 60646 59200 60702 59256
rect 61382 59064 61438 59120
rect 64326 59608 64382 59664
rect 64142 59200 64198 59256
rect 68466 59764 68522 59800
rect 68466 59744 68468 59764
rect 68468 59744 68520 59764
rect 68520 59744 68522 59764
rect 69294 59744 69350 59800
rect 70122 59764 70178 59800
rect 70122 59744 70124 59764
rect 70124 59744 70176 59764
rect 70176 59744 70178 59764
rect 66810 59608 66866 59664
rect 65338 59472 65394 59528
rect 65522 59336 65578 59392
rect 66902 59472 66958 59528
rect 66810 59200 66866 59256
rect 67638 59608 67694 59664
rect 67638 59336 67694 59392
rect 68282 59336 68338 59392
rect 71778 59744 71834 59800
rect 69294 59472 69350 59528
rect 71042 59472 71098 59528
rect 69662 59336 69718 59392
rect 81346 59744 81402 59800
rect 83462 59764 83518 59800
rect 83462 59744 83464 59764
rect 83464 59744 83516 59764
rect 83516 59744 83518 59764
rect 71778 59336 71834 59392
rect 71226 59200 71282 59256
rect 72422 59064 72478 59120
rect 74630 59608 74686 59664
rect 77574 59628 77630 59664
rect 77574 59608 77576 59628
rect 77576 59608 77628 59628
rect 77628 59608 77630 59628
rect 79874 59608 79930 59664
rect 73802 59472 73858 59528
rect 75550 59336 75606 59392
rect 76930 59472 76986 59528
rect 77114 59336 77170 59392
rect 79690 59336 79746 59392
rect 81254 59472 81310 59528
rect 87510 59744 87566 59800
rect 88430 59764 88486 59800
rect 88430 59744 88432 59764
rect 88432 59744 88484 59764
rect 88484 59744 88486 59764
rect 81806 59608 81862 59664
rect 84106 59472 84162 59528
rect 81806 59336 81862 59392
rect 82726 59336 82782 59392
rect 84014 59336 84070 59392
rect 91742 59764 91798 59800
rect 91742 59744 91744 59764
rect 91744 59744 91796 59764
rect 91796 59744 91798 59764
rect 98366 59764 98422 59800
rect 98366 59744 98368 59764
rect 98368 59744 98420 59764
rect 98420 59744 98422 59764
rect 100850 59764 100906 59800
rect 100850 59744 100852 59764
rect 100852 59744 100904 59764
rect 100904 59744 100906 59764
rect 102506 59744 102562 59800
rect 103426 59744 103482 59800
rect 107198 59744 107254 59800
rect 107474 59744 107530 59800
rect 111798 59744 111854 59800
rect 88430 59608 88486 59664
rect 88062 59472 88118 59528
rect 87786 59336 87842 59392
rect 90086 59608 90142 59664
rect 89166 59472 89222 59528
rect 93398 59608 93454 59664
rect 94318 59608 94374 59664
rect 91926 59472 91982 59528
rect 93122 59472 93178 59528
rect 93306 59472 93362 59528
rect 90086 59336 90142 59392
rect 90362 59336 90418 59392
rect 91834 59336 91890 59392
rect 93122 59200 93178 59256
rect 95974 59608 96030 59664
rect 94318 59336 94374 59392
rect 95882 59472 95938 59528
rect 95974 59336 96030 59392
rect 96710 59628 96766 59664
rect 96710 59608 96712 59628
rect 96712 59608 96764 59628
rect 96764 59608 96766 59628
rect 97262 59336 97318 59392
rect 98826 59472 98882 59528
rect 101402 59472 101458 59528
rect 100022 59336 100078 59392
rect 100206 59200 100262 59256
rect 102966 59608 103022 59664
rect 102506 59336 102562 59392
rect 105082 59628 105138 59664
rect 105082 59608 105084 59628
rect 105084 59608 105136 59628
rect 105136 59608 105138 59628
rect 103426 59472 103482 59528
rect 104346 59472 104402 59528
rect 104162 59336 104218 59392
rect 105542 59336 105598 59392
rect 107566 59608 107622 59664
rect 107106 59336 107162 59392
rect 108486 59472 108542 59528
rect 109222 59608 109278 59664
rect 110878 59628 110934 59664
rect 110878 59608 110880 59628
rect 110880 59608 110932 59628
rect 110932 59608 110934 59628
rect 108854 59336 108910 59392
rect 109038 59336 109094 59392
rect 111706 59608 111762 59664
rect 115018 59764 115074 59800
rect 115018 59744 115020 59764
rect 115020 59744 115072 59764
rect 115072 59744 115074 59764
rect 121642 59744 121698 59800
rect 111798 59472 111854 59528
rect 112994 59472 113050 59528
rect 111614 59336 111670 59392
rect 113546 59608 113602 59664
rect 119986 59628 120042 59664
rect 119986 59608 119988 59628
rect 119988 59608 120040 59628
rect 120040 59608 120042 59628
rect 120722 59608 120778 59664
rect 115202 59472 115258 59528
rect 113546 59336 113602 59392
rect 114190 59336 114246 59392
rect 117502 59492 117558 59528
rect 117502 59472 117504 59492
rect 117504 59472 117556 59492
rect 117556 59472 117558 59492
rect 116582 59336 116638 59392
rect 116766 59200 116822 59256
rect 119986 59472 120042 59528
rect 119526 59336 119582 59392
rect 120906 59472 120962 59528
rect 123298 59764 123354 59800
rect 123298 59744 123300 59764
rect 123300 59744 123352 59764
rect 123352 59744 123354 59764
rect 124218 59744 124274 59800
rect 122746 59608 122802 59664
rect 123482 59608 123538 59664
rect 121642 59336 121698 59392
rect 122102 59336 122158 59392
rect 127530 59764 127586 59800
rect 127530 59744 127532 59764
rect 127532 59744 127584 59764
rect 127584 59744 127586 59764
rect 136638 59764 136694 59800
rect 136638 59744 136640 59764
rect 136640 59744 136692 59764
rect 136692 59744 136694 59764
rect 139214 59744 139270 59800
rect 139950 59744 140006 59800
rect 124218 59336 124274 59392
rect 123666 59200 123722 59256
rect 125046 59472 125102 59528
rect 125874 59608 125930 59664
rect 131670 59628 131726 59664
rect 131670 59608 131672 59628
rect 131672 59608 131724 59628
rect 131724 59608 131726 59628
rect 134154 59628 134210 59664
rect 134154 59608 134156 59628
rect 134156 59608 134208 59628
rect 134208 59608 134210 59628
rect 125874 59336 125930 59392
rect 126242 59336 126298 59392
rect 127714 59336 127770 59392
rect 128358 59472 128414 59528
rect 129186 59200 129242 59256
rect 130382 59064 130438 59120
rect 133142 59472 133198 59528
rect 131854 59336 131910 59392
rect 133418 59336 133474 59392
rect 136638 59608 136694 59664
rect 138478 59608 138534 59664
rect 139122 59608 139178 59664
rect 137466 59472 137522 59528
rect 137282 59200 137338 59256
rect 137558 59356 137614 59392
rect 137558 59336 137560 59356
rect 137560 59336 137612 59356
rect 137612 59336 137614 59356
rect 138478 59336 138534 59392
rect 139214 59472 139270 59528
rect 141698 59744 141754 59800
rect 142434 59764 142490 59800
rect 142434 59744 142436 59764
rect 142436 59744 142488 59764
rect 142488 59744 142490 59764
rect 140042 59472 140098 59528
rect 139950 59336 140006 59392
rect 141606 59608 141662 59664
rect 144274 59744 144330 59800
rect 144182 59608 144238 59664
rect 141698 59472 141754 59528
rect 141606 58928 141662 58984
rect 149426 59764 149482 59800
rect 149426 59744 149428 59764
rect 149428 59744 149480 59764
rect 149480 59744 149482 59764
rect 146666 59608 146722 59664
rect 147494 59628 147550 59664
rect 147494 59608 147496 59628
rect 147496 59608 147548 59628
rect 147548 59608 147550 59628
rect 145562 59472 145618 59528
rect 144366 59336 144422 59392
rect 146666 59336 146722 59392
rect 148322 59336 148378 59392
rect 144182 3304 144238 3360
rect 149150 59608 149206 59664
rect 149702 59608 149758 59664
rect 149886 59472 149942 59528
rect 150806 59744 150862 59800
rect 152462 59764 152518 59800
rect 152462 59744 152464 59764
rect 152464 59744 152516 59764
rect 152516 59744 152518 59764
rect 156602 59764 156658 59800
rect 156602 59744 156604 59764
rect 156604 59744 156656 59764
rect 156656 59744 156658 59764
rect 159914 59744 159970 59800
rect 160742 59764 160798 59800
rect 160742 59744 160744 59764
rect 160744 59744 160796 59764
rect 160796 59744 160798 59764
rect 151726 59608 151782 59664
rect 153106 59472 153162 59528
rect 150254 59336 150310 59392
rect 150438 59336 150494 59392
rect 153014 59336 153070 59392
rect 156602 59608 156658 59664
rect 156970 59472 157026 59528
rect 155866 59336 155922 59392
rect 156602 59336 156658 59392
rect 157246 59472 157302 59528
rect 157338 59336 157394 59392
rect 167458 59764 167514 59800
rect 167458 59744 167460 59764
rect 167460 59744 167512 59764
rect 167512 59744 167514 59764
rect 174542 59744 174598 59800
rect 175738 59764 175794 59800
rect 175738 59744 175740 59764
rect 175740 59744 175792 59764
rect 175792 59744 175794 59764
rect 160006 59472 160062 59528
rect 161110 59472 161166 59528
rect 161294 59336 161350 59392
rect 162858 59608 162914 59664
rect 163870 59472 163926 59528
rect 164054 59336 164110 59392
rect 168286 59472 168342 59528
rect 166906 59336 166962 59392
rect 168102 59336 168158 59392
rect 165434 59200 165490 59256
rect 169942 59472 169998 59528
rect 171598 59472 171654 59528
rect 169390 59336 169446 59392
rect 169574 59336 169630 59392
rect 171046 59200 171102 59256
rect 172426 59200 172482 59256
rect 173806 59472 173862 59528
rect 182362 59764 182418 59800
rect 182362 59744 182364 59764
rect 182364 59744 182416 59764
rect 182416 59744 182418 59764
rect 183190 59744 183246 59800
rect 176474 59472 176530 59528
rect 178222 59492 178278 59528
rect 178222 59472 178224 59492
rect 178224 59472 178276 59492
rect 178276 59472 178278 59492
rect 175186 59336 175242 59392
rect 177670 59336 177726 59392
rect 177854 59200 177910 59256
rect 180706 59628 180762 59664
rect 180706 59608 180708 59628
rect 180708 59608 180760 59628
rect 180760 59608 180762 59628
rect 180706 59472 180762 59528
rect 181810 59336 181866 59392
rect 182362 59608 182418 59664
rect 185674 59764 185730 59800
rect 185674 59744 185676 59764
rect 185676 59744 185728 59764
rect 185728 59744 185730 59764
rect 187422 59744 187478 59800
rect 183190 59336 183246 59392
rect 183466 59200 183522 59256
rect 187330 59608 187386 59664
rect 186134 59472 186190 59528
rect 185950 59336 186006 59392
rect 184754 59200 184810 59256
rect 189906 59764 189962 59800
rect 189906 59744 189908 59764
rect 189908 59744 189960 59764
rect 189960 59744 189962 59764
rect 196530 59744 196586 59800
rect 201498 59744 201554 59800
rect 187422 59472 187478 59528
rect 187330 59336 187386 59392
rect 187606 59336 187662 59392
rect 190090 59472 190146 59528
rect 188894 59200 188950 59256
rect 191746 59608 191802 59664
rect 193034 59472 193090 59528
rect 190274 59336 190330 59392
rect 191562 59336 191618 59392
rect 191746 59336 191802 59392
rect 192850 59336 192906 59392
rect 194874 59472 194930 59528
rect 200670 59628 200726 59664
rect 200670 59608 200672 59628
rect 200672 59608 200724 59628
rect 200724 59608 200726 59628
rect 197174 59472 197230 59528
rect 194322 59336 194378 59392
rect 194506 59336 194562 59392
rect 196990 59336 197046 59392
rect 195886 59200 195942 59256
rect 198370 59200 198426 59256
rect 201130 59472 201186 59528
rect 200026 59200 200082 59256
rect 204810 59764 204866 59800
rect 204810 59744 204812 59764
rect 204812 59744 204864 59764
rect 204864 59744 204866 59764
rect 213182 59764 213238 59800
rect 213182 59744 213184 59764
rect 213184 59744 213236 59764
rect 213236 59744 213238 59764
rect 214010 59744 214066 59800
rect 202510 59472 202566 59528
rect 201498 59336 201554 59392
rect 201314 59200 201370 59256
rect 203154 59608 203210 59664
rect 205454 59472 205510 59528
rect 207294 59492 207350 59528
rect 207294 59472 207296 59492
rect 207296 59472 207348 59492
rect 207348 59472 207350 59492
rect 203154 59336 203210 59392
rect 204166 59336 204222 59392
rect 206650 59336 206706 59392
rect 206834 59200 206890 59256
rect 208306 59064 208362 59120
rect 210698 59608 210754 59664
rect 209870 59472 209926 59528
rect 209594 59336 209650 59392
rect 210698 59336 210754 59392
rect 213550 59608 213606 59664
rect 210974 59336 211030 59392
rect 212446 59200 212502 59256
rect 218150 59764 218206 59800
rect 218150 59744 218152 59764
rect 218152 59744 218204 59764
rect 218204 59744 218206 59764
rect 221462 59764 221518 59800
rect 221462 59744 221464 59764
rect 221464 59744 221516 59764
rect 221516 59744 221518 59764
rect 215758 59608 215814 59664
rect 214930 59472 214986 59528
rect 214010 59336 214066 59392
rect 213734 59200 213790 59256
rect 215758 59336 215814 59392
rect 215942 59336 215998 59392
rect 219070 59472 219126 59528
rect 217874 59200 217930 59256
rect 217690 59064 217746 59120
rect 219806 59608 219862 59664
rect 222106 59472 222162 59528
rect 219806 59336 219862 59392
rect 220726 59336 220782 59392
rect 222014 59336 222070 59392
rect 223486 59200 223542 59256
rect 225234 59744 225290 59800
rect 232778 59744 232834 59800
rect 235262 59744 235318 59800
rect 235446 59744 235502 59800
rect 236918 59744 236974 59800
rect 224958 59608 225014 59664
rect 224774 59472 224830 59528
rect 228914 59628 228970 59664
rect 228914 59608 228916 59628
rect 228916 59608 228968 59628
rect 228968 59608 228970 59628
rect 226154 59472 226210 59528
rect 224958 59336 225014 59392
rect 225970 59336 226026 59392
rect 229006 59472 229062 59528
rect 231766 59472 231822 59528
rect 228914 59336 228970 59392
rect 230202 59200 230258 59256
rect 234250 59608 234306 59664
rect 232962 59336 233018 59392
rect 235906 59472 235962 59528
rect 235446 59336 235502 59392
rect 239954 59744 240010 59800
rect 240598 59764 240654 59800
rect 240598 59744 240600 59764
rect 240600 59744 240652 59764
rect 240652 59744 240654 59764
rect 238390 59608 238446 59664
rect 237286 59336 237342 59392
rect 244738 59764 244794 59800
rect 244738 59744 244740 59764
rect 244740 59744 244792 59764
rect 244792 59744 244794 59764
rect 249706 59764 249762 59800
rect 249706 59744 249708 59764
rect 249708 59744 249760 59764
rect 249760 59744 249762 59764
rect 250534 59744 250590 59800
rect 241334 59472 241390 59528
rect 240046 59336 240102 59392
rect 241150 59336 241206 59392
rect 242530 59200 242586 59256
rect 244186 59608 244242 59664
rect 245474 59472 245530 59528
rect 245290 59336 245346 59392
rect 246854 59200 246910 59256
rect 248878 59472 248934 59528
rect 249706 59608 249762 59664
rect 253202 59764 253258 59800
rect 253202 59744 253204 59764
rect 253204 59744 253256 59764
rect 253256 59744 253258 59764
rect 257434 59744 257490 59800
rect 267738 59764 267794 59800
rect 267738 59744 267740 59764
rect 267740 59744 267792 59764
rect 267792 59744 267794 59764
rect 251086 59472 251142 59528
rect 249614 59336 249670 59392
rect 250534 59336 250590 59392
rect 250994 59336 251050 59392
rect 252282 59608 252338 59664
rect 253386 59608 253442 59664
rect 255594 59608 255650 59664
rect 252282 59336 252338 59392
rect 253202 59336 253258 59392
rect 254766 59472 254822 59528
rect 254582 59200 254638 59256
rect 257250 59628 257306 59664
rect 257250 59608 257252 59628
rect 257252 59608 257304 59628
rect 257304 59608 257306 59628
rect 255594 59336 255650 59392
rect 272706 59764 272762 59800
rect 272706 59744 272708 59764
rect 272708 59744 272760 59764
rect 272760 59744 272762 59764
rect 276846 59764 276902 59800
rect 276846 59744 276848 59764
rect 276848 59744 276900 59764
rect 276900 59744 276902 59764
rect 280066 59744 280122 59800
rect 286782 59764 286838 59800
rect 286782 59744 286784 59764
rect 286784 59744 286836 59764
rect 286836 59744 286838 59764
rect 258906 59608 258962 59664
rect 260562 59628 260618 59664
rect 260562 59608 260564 59628
rect 260564 59608 260616 59628
rect 260616 59608 260618 59628
rect 258078 59472 258134 59528
rect 257434 59336 257490 59392
rect 257526 59200 257582 59256
rect 260562 59492 260618 59528
rect 260562 59472 260564 59492
rect 260564 59472 260616 59492
rect 260616 59472 260618 59492
rect 267738 59472 267794 59528
rect 258906 59336 258962 59392
rect 260102 59336 260158 59392
rect 262126 59200 262182 59256
rect 262034 59064 262090 59120
rect 268198 59472 268254 59528
rect 268014 59200 268070 59256
rect 271878 59472 271934 59528
rect 270682 59200 270738 59256
rect 271970 59336 272026 59392
rect 273350 59200 273406 59256
rect 276294 59472 276350 59528
rect 274914 59200 274970 59256
rect 276110 59200 276166 59256
rect 277398 59336 277454 59392
rect 277490 59200 277546 59256
rect 287058 59744 287114 59800
rect 285126 59608 285182 59664
rect 280158 59472 280214 59528
rect 282642 59492 282698 59528
rect 282642 59472 282644 59492
rect 282644 59472 282696 59492
rect 282696 59472 282698 59492
rect 280342 59336 280398 59392
rect 282918 59336 282974 59392
rect 284390 59336 284446 59392
rect 281538 59200 281594 59256
rect 285678 59472 285734 59528
rect 285126 59336 285182 59392
rect 291842 59764 291898 59800
rect 291842 59744 291844 59764
rect 291844 59744 291896 59764
rect 291896 59744 291898 59764
rect 300122 59764 300178 59800
rect 300122 59744 300124 59764
rect 300124 59744 300176 59764
rect 300176 59744 300178 59764
rect 300950 59744 301006 59800
rect 301778 59744 301834 59800
rect 287426 59336 287482 59392
rect 287242 59200 287298 59256
rect 293498 59628 293554 59664
rect 293498 59608 293500 59628
rect 293500 59608 293552 59628
rect 293552 59608 293554 59628
rect 288622 59472 288678 59528
rect 291566 59472 291622 59528
rect 294050 59472 294106 59528
rect 291382 59200 291438 59256
rect 292670 59336 292726 59392
rect 295982 59608 296038 59664
rect 296810 59628 296866 59664
rect 296810 59608 296812 59628
rect 296812 59608 296864 59628
rect 296864 59608 296866 59628
rect 296718 59472 296774 59528
rect 295982 59336 296038 59392
rect 295706 59200 295762 59256
rect 300122 59472 300178 59528
rect 298926 59200 298982 59256
rect 303434 59764 303490 59800
rect 303434 59744 303436 59764
rect 303436 59744 303488 59764
rect 303488 59744 303490 59764
rect 305366 59744 305422 59800
rect 301502 59608 301558 59664
rect 300950 59336 301006 59392
rect 300306 59200 300362 59256
rect 302882 59336 302938 59392
rect 304262 59472 304318 59528
rect 305826 59744 305882 59800
rect 309322 59744 309378 59800
rect 310702 59764 310758 59800
rect 310702 59744 310704 59764
rect 310704 59744 310756 59764
rect 310756 59744 310758 59764
rect 305366 59336 305422 59392
rect 305918 59628 305974 59664
rect 305918 59608 305920 59628
rect 305920 59608 305972 59628
rect 305972 59608 305974 59628
rect 306746 59492 306802 59528
rect 306746 59472 306748 59492
rect 306748 59472 306800 59492
rect 306800 59472 306802 59492
rect 307206 59336 307262 59392
rect 311806 59744 311862 59800
rect 309874 59472 309930 59528
rect 310702 59472 310758 59528
rect 309322 59336 309378 59392
rect 313462 59744 313518 59800
rect 314290 59780 314292 59800
rect 314292 59780 314344 59800
rect 314344 59780 314346 59800
rect 314290 59744 314346 59780
rect 315394 59780 315396 59800
rect 315396 59780 315448 59800
rect 315448 59780 315450 59800
rect 315394 59744 315450 59780
rect 316590 59744 316646 59800
rect 311346 59336 311402 59392
rect 311806 59336 311862 59392
rect 312726 59472 312782 59528
rect 314290 59608 314346 59664
rect 313462 59336 313518 59392
rect 313922 59200 313978 59256
rect 316590 59628 316646 59664
rect 316590 59608 316592 59628
rect 316592 59608 316644 59628
rect 316644 59608 316646 59628
rect 316590 59472 316646 59528
rect 315302 59336 315358 59392
rect 318430 59764 318486 59800
rect 318430 59744 318432 59764
rect 318432 59744 318484 59764
rect 318484 59744 318486 59764
rect 319258 59744 319314 59800
rect 320822 59744 320878 59800
rect 325054 59744 325110 59800
rect 325882 59744 325938 59800
rect 326710 59764 326766 59800
rect 326710 59744 326712 59764
rect 326712 59744 326764 59764
rect 326764 59744 326766 59764
rect 319442 59472 319498 59528
rect 319626 59336 319682 59392
rect 321742 59492 321798 59528
rect 321742 59472 321744 59492
rect 321744 59472 321796 59492
rect 321796 59472 321798 59492
rect 321742 59336 321798 59392
rect 324962 59472 325018 59528
rect 330114 59744 330170 59800
rect 326342 59608 326398 59664
rect 325054 59336 325110 59392
rect 325882 59336 325938 59392
rect 328366 59608 328422 59664
rect 327906 59336 327962 59392
rect 328366 59336 328422 59392
rect 329286 59472 329342 59528
rect 330942 59744 330998 59800
rect 337382 59744 337438 59800
rect 337566 59764 337622 59800
rect 337566 59744 337568 59764
rect 337568 59744 337620 59764
rect 337620 59744 337622 59764
rect 330850 59608 330906 59664
rect 330482 59472 330538 59528
rect 330114 59336 330170 59392
rect 331770 59492 331826 59528
rect 331770 59472 331772 59492
rect 331772 59472 331824 59492
rect 331824 59472 331826 59492
rect 331770 59336 331826 59392
rect 335082 59608 335138 59664
rect 333426 59492 333482 59528
rect 333426 59472 333428 59492
rect 333428 59472 333480 59492
rect 333480 59472 333482 59492
rect 336002 59472 336058 59528
rect 334622 59336 334678 59392
rect 335082 59336 335138 59392
rect 341614 59744 341670 59800
rect 345018 59764 345074 59800
rect 345018 59744 345020 59764
rect 345020 59744 345072 59764
rect 345072 59744 345074 59764
rect 337474 59608 337530 59664
rect 339222 59608 339278 59664
rect 337198 59336 337254 59392
rect 337382 59336 337438 59392
rect 340142 59472 340198 59528
rect 338854 59336 338910 59392
rect 339222 59336 339278 59392
rect 341522 59608 341578 59664
rect 350630 59744 350686 59800
rect 351734 59744 351790 59800
rect 356702 59764 356758 59800
rect 356702 59744 356704 59764
rect 356704 59744 356756 59764
rect 356756 59744 356758 59764
rect 342350 59628 342406 59664
rect 342350 59608 342352 59628
rect 342352 59608 342404 59628
rect 342404 59608 342406 59628
rect 343362 59608 343418 59664
rect 341614 59472 341670 59528
rect 345018 59608 345074 59664
rect 344282 59472 344338 59528
rect 341614 59336 341670 59392
rect 342902 59336 342958 59392
rect 343362 59336 343418 59392
rect 345018 59336 345074 59392
rect 347502 59492 347558 59528
rect 347502 59472 347504 59492
rect 347504 59472 347556 59492
rect 347556 59472 347558 59492
rect 349802 59472 349858 59528
rect 348606 59336 348662 59392
rect 348422 59200 348478 59256
rect 350906 59608 350962 59664
rect 357530 59780 357532 59800
rect 357532 59780 357584 59800
rect 357584 59780 357586 59800
rect 357530 59744 357586 59780
rect 353390 59628 353446 59664
rect 353390 59608 353392 59628
rect 353392 59608 353444 59628
rect 353444 59608 353446 59628
rect 354218 59608 354274 59664
rect 354034 59472 354090 59528
rect 352746 58928 352802 58984
rect 357530 59608 357586 59664
rect 354218 59336 354274 59392
rect 356702 59472 356758 59528
rect 356886 59200 356942 59256
rect 360842 59764 360898 59800
rect 360842 59744 360844 59764
rect 360844 59744 360896 59764
rect 360896 59744 360898 59764
rect 361578 59744 361634 59800
rect 360842 59472 360898 59528
rect 360106 59336 360162 59392
rect 369122 59744 369178 59800
rect 369490 59744 369546 59800
rect 361670 59608 361726 59664
rect 361578 59336 361634 59392
rect 362498 59492 362554 59528
rect 362498 59472 362500 59492
rect 362500 59472 362552 59492
rect 362552 59472 362554 59492
rect 363050 59200 363106 59256
rect 369030 59628 369086 59664
rect 369030 59608 369032 59628
rect 369032 59608 369084 59628
rect 369084 59608 369086 59628
rect 364798 59492 364854 59528
rect 364798 59472 364800 59492
rect 364800 59472 364852 59492
rect 364852 59472 364854 59492
rect 366638 59492 366694 59528
rect 366638 59472 366640 59492
rect 366640 59472 366692 59492
rect 366692 59472 366694 59492
rect 368478 59472 368534 59528
rect 364338 59336 364394 59392
rect 367282 59336 367338 59392
rect 367098 59200 367154 59256
rect 369122 59336 369178 59392
rect 376482 59744 376538 59800
rect 376666 59744 376722 59800
rect 379978 59764 380034 59800
rect 379978 59744 379980 59764
rect 379980 59744 380032 59764
rect 380032 59744 380034 59764
rect 372526 59608 372582 59664
rect 373814 59608 373870 59664
rect 369398 3304 369454 3360
rect 372618 59472 372674 59528
rect 372526 59336 372582 59392
rect 371422 59200 371478 59256
rect 374182 59336 374238 59392
rect 372710 59200 372766 59256
rect 375654 59336 375710 59392
rect 376482 59336 376538 59392
rect 381634 59744 381690 59800
rect 389454 59744 389510 59800
rect 398838 59744 398894 59800
rect 376942 59608 376998 59664
rect 376758 59472 376814 59528
rect 379702 59472 379758 59528
rect 378230 59336 378286 59392
rect 380898 59200 380954 59256
rect 383106 59608 383162 59664
rect 384118 59628 384174 59664
rect 384118 59608 384120 59628
rect 384120 59608 384172 59628
rect 384172 59608 384174 59628
rect 387430 59608 387486 59664
rect 383934 59472 383990 59528
rect 382370 59336 382426 59392
rect 383106 59336 383162 59392
rect 381634 59200 381690 59256
rect 383750 59200 383806 59256
rect 385222 59200 385278 59256
rect 385774 59492 385830 59528
rect 385774 59472 385776 59492
rect 385776 59472 385828 59492
rect 385828 59472 385830 59492
rect 387982 59472 388038 59528
rect 386418 59336 386474 59392
rect 387430 59336 387486 59392
rect 389362 59200 389418 59256
rect 393318 59628 393374 59664
rect 393318 59608 393320 59628
rect 393320 59608 393372 59628
rect 393372 59608 393374 59628
rect 390558 59472 390614 59528
rect 393318 59472 393374 59528
rect 389546 59336 389602 59392
rect 392122 59200 392178 59256
rect 394698 59472 394754 59528
rect 393594 59200 393650 59256
rect 397550 59472 397606 59528
rect 396354 59336 396410 59392
rect 396170 59200 396226 59256
rect 400678 59744 400734 59800
rect 400954 59744 401010 59800
rect 401782 59744 401838 59800
rect 406566 59764 406622 59800
rect 406566 59744 406568 59764
rect 406568 59744 406620 59764
rect 406620 59744 406622 59764
rect 400310 59472 400366 59528
rect 401506 59472 401562 59528
rect 398930 59336 398986 59392
rect 399114 59336 399170 59392
rect 400494 59336 400550 59392
rect 401598 59200 401654 59256
rect 409050 59764 409106 59800
rect 409050 59744 409052 59764
rect 409052 59744 409104 59764
rect 409104 59744 409106 59764
rect 412822 59744 412878 59800
rect 417606 59764 417662 59800
rect 422390 59780 422392 59800
rect 422392 59780 422444 59800
rect 422444 59780 422446 59800
rect 417606 59744 417608 59764
rect 417608 59744 417660 59764
rect 417660 59744 417662 59764
rect 405738 59472 405794 59528
rect 402978 59200 403034 59256
rect 404542 59200 404598 59256
rect 405830 59336 405886 59392
rect 407210 59336 407266 59392
rect 408774 59472 408830 59528
rect 409970 59200 410026 59256
rect 411534 59608 411590 59664
rect 412362 59608 412418 59664
rect 412730 59608 412786 59664
rect 412362 59472 412418 59528
rect 411534 59336 411590 59392
rect 411258 59200 411314 59256
rect 422390 59744 422446 59780
rect 414110 59608 414166 59664
rect 414110 59472 414166 59528
rect 412914 59336 412970 59392
rect 417606 59608 417662 59664
rect 417054 59336 417110 59392
rect 416870 59200 416926 59256
rect 418250 59472 418306 59528
rect 419078 59492 419134 59528
rect 419078 59472 419080 59492
rect 419080 59472 419132 59492
rect 419132 59472 419134 59492
rect 420734 59608 420790 59664
rect 422114 59608 422170 59664
rect 422298 59608 422354 59664
rect 421102 59472 421158 59528
rect 420734 59336 420790 59392
rect 419630 3576 419686 3632
rect 425702 59764 425758 59800
rect 425702 59744 425704 59764
rect 425704 59744 425756 59764
rect 425756 59744 425758 59764
rect 428094 59744 428150 59800
rect 429014 59744 429070 59800
rect 429842 59764 429898 59800
rect 429842 59744 429844 59764
rect 429844 59744 429896 59764
rect 429896 59744 429898 59764
rect 425058 59472 425114 59528
rect 425150 59336 425206 59392
rect 426530 59336 426586 59392
rect 435822 59764 435878 59800
rect 435822 59744 435824 59764
rect 435824 59744 435876 59764
rect 435876 59744 435878 59764
rect 438214 59744 438270 59800
rect 429198 59608 429254 59664
rect 430578 59608 430634 59664
rect 428186 59472 428242 59528
rect 429014 59472 429070 59528
rect 428094 59336 428150 59392
rect 430670 59472 430726 59528
rect 431774 59472 431830 59528
rect 429290 59336 429346 59392
rect 430578 59336 430634 59392
rect 432142 59336 432198 59392
rect 438766 59744 438822 59800
rect 440698 59744 440754 59800
rect 441250 59744 441306 59800
rect 442354 59764 442410 59800
rect 442354 59744 442356 59764
rect 442356 59744 442408 59764
rect 442408 59744 442410 59764
rect 433982 59608 434038 59664
rect 433522 59336 433578 59392
rect 434810 59472 434866 59528
rect 438122 59472 438178 59528
rect 433982 59336 434038 59392
rect 436742 59336 436798 59392
rect 436098 59200 436154 59256
rect 439502 59472 439558 59528
rect 440698 59472 440754 59528
rect 438766 59336 438822 59392
rect 445666 59764 445722 59800
rect 445666 59744 445668 59764
rect 445668 59744 445720 59764
rect 445720 59744 445722 59764
rect 450542 59744 450598 59800
rect 454774 59744 454830 59800
rect 455602 59744 455658 59800
rect 456522 59764 456578 59800
rect 456522 59744 456524 59764
rect 456524 59744 456576 59764
rect 456576 59744 456578 59764
rect 442262 59608 442318 59664
rect 444010 59608 444066 59664
rect 441066 59336 441122 59392
rect 441250 59336 441306 59392
rect 442354 59472 442410 59528
rect 445022 59472 445078 59528
rect 443642 59336 443698 59392
rect 444010 59336 444066 59392
rect 445666 59608 445722 59664
rect 446402 59508 446404 59528
rect 446404 59508 446456 59528
rect 446456 59508 446458 59528
rect 446402 59472 446458 59508
rect 446402 59336 446458 59392
rect 448150 59492 448206 59528
rect 448150 59472 448152 59492
rect 448152 59472 448204 59492
rect 448204 59472 448206 59492
rect 450450 59472 450506 59528
rect 449162 59336 449218 59392
rect 450634 59628 450690 59664
rect 450634 59608 450636 59628
rect 450636 59608 450688 59628
rect 450688 59608 450690 59628
rect 450542 59336 450598 59392
rect 451278 59356 451334 59392
rect 451278 59336 451280 59356
rect 451280 59336 451332 59356
rect 451332 59336 451334 59356
rect 452290 59492 452346 59528
rect 452290 59472 452292 59492
rect 452292 59472 452344 59492
rect 452344 59472 452346 59492
rect 454682 59472 454738 59528
rect 453302 59336 453358 59392
rect 461490 59764 461546 59800
rect 461490 59744 461492 59764
rect 461492 59744 461544 59764
rect 461544 59744 461546 59764
rect 467930 59744 467986 59800
rect 456062 59608 456118 59664
rect 455602 59336 455658 59392
rect 458178 59628 458234 59664
rect 458178 59608 458180 59628
rect 458180 59608 458232 59628
rect 458232 59608 458234 59628
rect 457626 59336 457682 59392
rect 458914 59608 458970 59664
rect 460478 59608 460534 59664
rect 459006 59472 459062 59528
rect 458914 59336 458970 59392
rect 461490 59472 461546 59528
rect 460478 59336 460534 59392
rect 461490 59356 461546 59392
rect 461490 59336 461492 59356
rect 461492 59336 461544 59356
rect 461544 59336 461546 59356
rect 461766 59200 461822 59256
rect 464802 59608 464858 59664
rect 467102 59608 467158 59664
rect 463146 59492 463202 59528
rect 463146 59472 463148 59492
rect 463148 59472 463200 59492
rect 463200 59472 463202 59492
rect 465722 59472 465778 59528
rect 464342 59336 464398 59392
rect 464802 59336 464858 59392
rect 467286 59336 467342 59392
rect 472622 59608 472678 59664
rect 471426 59472 471482 59528
rect 471242 59336 471298 59392
rect 470138 59200 470194 59256
rect 471426 3304 471482 3360
rect 583390 3304 583446 3360
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 59494 449326 60076 449386
rect 57605 449306 57671 449309
rect 59494 449306 59554 449326
rect 57605 449304 59554 449306
rect 57605 449248 57610 449304
rect 57666 449248 59554 449304
rect 57605 449246 59554 449248
rect 57605 449243 57671 449246
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 57973 59530 58039 59533
rect 60802 59530 60862 60044
rect 57973 59528 60862 59530
rect 57973 59472 57978 59528
rect 58034 59472 60862 59528
rect 57973 59470 60862 59472
rect 57973 59467 58039 59470
rect 58617 59394 58683 59397
rect 61633 59394 61693 60044
rect 62465 59394 62525 60044
rect 62665 59666 62731 59669
rect 63296 59666 63356 60044
rect 64128 59938 64188 60044
rect 62665 59664 63356 59666
rect 62665 59608 62670 59664
rect 62726 59608 63356 59664
rect 62665 59606 63356 59608
rect 63726 59878 64188 59938
rect 62665 59603 62731 59606
rect 63726 59530 63786 59878
rect 64229 59802 64295 59805
rect 64960 59802 65020 60044
rect 64229 59800 65020 59802
rect 64229 59744 64234 59800
rect 64290 59744 65020 59800
rect 64229 59742 65020 59744
rect 65333 59802 65399 59805
rect 65791 59802 65851 60044
rect 65333 59800 65851 59802
rect 65333 59744 65338 59800
rect 65394 59744 65851 59800
rect 65333 59742 65851 59744
rect 64229 59739 64295 59742
rect 65333 59739 65399 59742
rect 64321 59666 64387 59669
rect 66623 59666 66683 60044
rect 64321 59664 66683 59666
rect 64321 59608 64326 59664
rect 64382 59608 66683 59664
rect 64321 59606 66683 59608
rect 66805 59666 66871 59669
rect 67454 59666 67514 60044
rect 66805 59664 67514 59666
rect 66805 59608 66810 59664
rect 66866 59608 67514 59664
rect 66805 59606 67514 59608
rect 67633 59666 67699 59669
rect 68286 59666 68346 60044
rect 68461 59802 68527 59805
rect 69118 59802 69178 60044
rect 68461 59800 69178 59802
rect 68461 59744 68466 59800
rect 68522 59744 69178 59800
rect 68461 59742 69178 59744
rect 69289 59802 69355 59805
rect 69949 59802 70009 60044
rect 69289 59800 70009 59802
rect 69289 59744 69294 59800
rect 69350 59744 70009 59800
rect 69289 59742 70009 59744
rect 70117 59802 70183 59805
rect 70781 59802 70841 60044
rect 70117 59800 70841 59802
rect 70117 59744 70122 59800
rect 70178 59744 70841 59800
rect 70117 59742 70841 59744
rect 68461 59739 68527 59742
rect 69289 59739 69355 59742
rect 70117 59739 70183 59742
rect 71612 59666 71672 60044
rect 72444 59938 72504 60044
rect 71822 59878 72504 59938
rect 71822 59805 71882 59878
rect 71773 59800 71882 59805
rect 71773 59744 71778 59800
rect 71834 59744 71882 59800
rect 71773 59742 71882 59744
rect 71773 59739 71839 59742
rect 67633 59664 68346 59666
rect 67633 59608 67638 59664
rect 67694 59608 68346 59664
rect 67633 59606 68346 59608
rect 70166 59606 71672 59666
rect 64321 59603 64387 59606
rect 66805 59603 66871 59606
rect 67633 59603 67699 59606
rect 65333 59530 65399 59533
rect 58617 59392 61693 59394
rect 58617 59336 58622 59392
rect 58678 59336 61693 59392
rect 58617 59334 61693 59336
rect 61886 59334 62525 59394
rect 62622 59470 63786 59530
rect 64128 59528 65399 59530
rect 64128 59472 65338 59528
rect 65394 59472 65399 59528
rect 64128 59470 65399 59472
rect 58617 59331 58683 59334
rect 60641 59258 60707 59261
rect 61886 59258 61946 59334
rect 60641 59256 61946 59258
rect 60641 59200 60646 59256
rect 60702 59200 61946 59256
rect 60641 59198 61946 59200
rect 60641 59195 60707 59198
rect 61377 59122 61443 59125
rect 62622 59122 62682 59470
rect 62757 59394 62823 59397
rect 64128 59394 64188 59470
rect 65333 59467 65399 59470
rect 66897 59530 66963 59533
rect 69289 59530 69355 59533
rect 70166 59530 70226 59606
rect 66897 59528 69355 59530
rect 66897 59472 66902 59528
rect 66958 59472 69294 59528
rect 69350 59472 69355 59528
rect 66897 59470 69355 59472
rect 66897 59467 66963 59470
rect 69289 59467 69355 59470
rect 69430 59470 70226 59530
rect 71037 59530 71103 59533
rect 73276 59530 73336 60044
rect 74107 59938 74167 60044
rect 71037 59528 73336 59530
rect 71037 59472 71042 59528
rect 71098 59472 73336 59528
rect 71037 59470 73336 59472
rect 73478 59878 74167 59938
rect 65517 59394 65583 59397
rect 67633 59394 67699 59397
rect 62757 59392 64188 59394
rect 62757 59336 62762 59392
rect 62818 59336 64188 59392
rect 62757 59334 64188 59336
rect 64462 59334 65442 59394
rect 62757 59331 62823 59334
rect 64137 59258 64203 59261
rect 64462 59258 64522 59334
rect 64137 59256 64522 59258
rect 64137 59200 64142 59256
rect 64198 59200 64522 59256
rect 64137 59198 64522 59200
rect 65382 59258 65442 59334
rect 65517 59392 67699 59394
rect 65517 59336 65522 59392
rect 65578 59336 67638 59392
rect 67694 59336 67699 59392
rect 65517 59334 67699 59336
rect 65517 59331 65583 59334
rect 67633 59331 67699 59334
rect 68277 59394 68343 59397
rect 69430 59394 69490 59470
rect 71037 59467 71103 59470
rect 68277 59392 69490 59394
rect 68277 59336 68282 59392
rect 68338 59336 69490 59392
rect 68277 59334 69490 59336
rect 69657 59394 69723 59397
rect 71773 59394 71839 59397
rect 73478 59394 73538 59878
rect 74939 59802 74999 60044
rect 74490 59742 74999 59802
rect 74490 59666 74550 59742
rect 69657 59392 71839 59394
rect 69657 59336 69662 59392
rect 69718 59336 71778 59392
rect 71834 59336 71839 59392
rect 69657 59334 71839 59336
rect 68277 59331 68343 59334
rect 69657 59331 69723 59334
rect 71773 59331 71839 59334
rect 72742 59334 73538 59394
rect 73662 59606 74550 59666
rect 74625 59666 74691 59669
rect 75770 59666 75830 60044
rect 74625 59664 75830 59666
rect 74625 59608 74630 59664
rect 74686 59608 75830 59664
rect 74625 59606 75830 59608
rect 66805 59258 66871 59261
rect 65382 59256 66871 59258
rect 65382 59200 66810 59256
rect 66866 59200 66871 59256
rect 65382 59198 66871 59200
rect 64137 59195 64203 59198
rect 66805 59195 66871 59198
rect 71221 59258 71287 59261
rect 72742 59258 72802 59334
rect 71221 59256 72802 59258
rect 71221 59200 71226 59256
rect 71282 59200 72802 59256
rect 71221 59198 72802 59200
rect 71221 59195 71287 59198
rect 61377 59120 62682 59122
rect 61377 59064 61382 59120
rect 61438 59064 62682 59120
rect 61377 59062 62682 59064
rect 72417 59122 72483 59125
rect 73662 59122 73722 59606
rect 74625 59603 74691 59606
rect 73797 59530 73863 59533
rect 76602 59530 76662 60044
rect 77434 59666 77494 60044
rect 73797 59528 76662 59530
rect 73797 59472 73802 59528
rect 73858 59472 76662 59528
rect 73797 59470 76662 59472
rect 76790 59606 77494 59666
rect 77569 59666 77635 59669
rect 78265 59666 78325 60044
rect 77569 59664 78325 59666
rect 77569 59608 77574 59664
rect 77630 59608 78325 59664
rect 77569 59606 78325 59608
rect 73797 59467 73863 59470
rect 75545 59394 75611 59397
rect 76790 59394 76850 59606
rect 77569 59603 77635 59606
rect 76925 59530 76991 59533
rect 79097 59530 79157 60044
rect 79928 59802 79988 60044
rect 76925 59528 79157 59530
rect 76925 59472 76930 59528
rect 76986 59472 79157 59528
rect 76925 59470 79157 59472
rect 79366 59742 79988 59802
rect 80760 59802 80820 60044
rect 81341 59802 81407 59805
rect 80760 59800 81407 59802
rect 80760 59744 81346 59800
rect 81402 59744 81407 59800
rect 80760 59742 81407 59744
rect 76925 59467 76991 59470
rect 75545 59392 76850 59394
rect 75545 59336 75550 59392
rect 75606 59336 76850 59392
rect 75545 59334 76850 59336
rect 77109 59394 77175 59397
rect 79366 59394 79426 59742
rect 81341 59739 81407 59742
rect 79869 59666 79935 59669
rect 81592 59666 81652 60044
rect 79869 59664 81652 59666
rect 79869 59608 79874 59664
rect 79930 59608 81652 59664
rect 79869 59606 81652 59608
rect 81801 59666 81867 59669
rect 82423 59666 82483 60044
rect 81801 59664 82483 59666
rect 81801 59608 81806 59664
rect 81862 59608 82483 59664
rect 81801 59606 82483 59608
rect 79869 59603 79935 59606
rect 81801 59603 81867 59606
rect 81249 59530 81315 59533
rect 83255 59530 83315 60044
rect 83457 59802 83523 59805
rect 84086 59802 84146 60044
rect 83457 59800 84146 59802
rect 83457 59744 83462 59800
rect 83518 59744 84146 59800
rect 83457 59742 84146 59744
rect 83457 59739 83523 59742
rect 84918 59666 84978 60044
rect 81249 59528 83315 59530
rect 81249 59472 81254 59528
rect 81310 59472 83315 59528
rect 81249 59470 83315 59472
rect 83414 59606 84978 59666
rect 81249 59467 81315 59470
rect 77109 59392 79426 59394
rect 77109 59336 77114 59392
rect 77170 59336 79426 59392
rect 77109 59334 79426 59336
rect 79685 59394 79751 59397
rect 81801 59394 81867 59397
rect 79685 59392 81867 59394
rect 79685 59336 79690 59392
rect 79746 59336 81806 59392
rect 81862 59336 81867 59392
rect 79685 59334 81867 59336
rect 75545 59331 75611 59334
rect 77109 59331 77175 59334
rect 79685 59331 79751 59334
rect 81801 59331 81867 59334
rect 82721 59394 82787 59397
rect 83414 59394 83474 59606
rect 84101 59530 84167 59533
rect 85750 59530 85810 60044
rect 84101 59528 85810 59530
rect 84101 59472 84106 59528
rect 84162 59472 85810 59528
rect 84101 59470 85810 59472
rect 84101 59467 84167 59470
rect 82721 59392 83474 59394
rect 82721 59336 82726 59392
rect 82782 59336 83474 59392
rect 82721 59334 83474 59336
rect 84009 59394 84075 59397
rect 86581 59394 86641 60044
rect 87413 59938 87473 60044
rect 88244 59938 88304 60044
rect 87278 59878 87473 59938
rect 87646 59878 88304 59938
rect 87278 59666 87338 59878
rect 87505 59802 87571 59805
rect 87646 59802 87706 59878
rect 87505 59800 87706 59802
rect 87505 59744 87510 59800
rect 87566 59744 87706 59800
rect 87505 59742 87706 59744
rect 88425 59802 88491 59805
rect 89076 59802 89136 60044
rect 88425 59800 89136 59802
rect 88425 59744 88430 59800
rect 88486 59744 89136 59800
rect 88425 59742 89136 59744
rect 87505 59739 87571 59742
rect 88425 59739 88491 59742
rect 88425 59666 88491 59669
rect 89908 59666 89968 60044
rect 87278 59606 87473 59666
rect 87413 59530 87473 59606
rect 88425 59664 89968 59666
rect 88425 59608 88430 59664
rect 88486 59608 89968 59664
rect 88425 59606 89968 59608
rect 90081 59666 90147 59669
rect 90739 59666 90799 60044
rect 90081 59664 90799 59666
rect 90081 59608 90086 59664
rect 90142 59608 90799 59664
rect 90081 59606 90799 59608
rect 88425 59603 88491 59606
rect 90081 59603 90147 59606
rect 88057 59530 88123 59533
rect 87413 59528 88123 59530
rect 87413 59472 88062 59528
rect 88118 59472 88123 59528
rect 87413 59470 88123 59472
rect 88057 59467 88123 59470
rect 89161 59530 89227 59533
rect 91571 59530 91631 60044
rect 91737 59802 91803 59805
rect 92402 59802 92462 60044
rect 91737 59800 92462 59802
rect 91737 59744 91742 59800
rect 91798 59744 92462 59800
rect 91737 59742 92462 59744
rect 91737 59739 91803 59742
rect 93234 59666 93294 60044
rect 89161 59528 91631 59530
rect 89161 59472 89166 59528
rect 89222 59472 91631 59528
rect 89161 59470 91631 59472
rect 91694 59606 93294 59666
rect 93393 59666 93459 59669
rect 94066 59666 94126 60044
rect 93393 59664 94126 59666
rect 93393 59608 93398 59664
rect 93454 59608 94126 59664
rect 93393 59606 94126 59608
rect 94313 59666 94379 59669
rect 94897 59666 94957 60044
rect 94313 59664 94957 59666
rect 94313 59608 94318 59664
rect 94374 59608 94957 59664
rect 94313 59606 94957 59608
rect 89161 59467 89227 59470
rect 84009 59392 86641 59394
rect 84009 59336 84014 59392
rect 84070 59336 86641 59392
rect 84009 59334 86641 59336
rect 87781 59394 87847 59397
rect 90081 59394 90147 59397
rect 87781 59392 90147 59394
rect 87781 59336 87786 59392
rect 87842 59336 90086 59392
rect 90142 59336 90147 59392
rect 87781 59334 90147 59336
rect 82721 59331 82787 59334
rect 84009 59331 84075 59334
rect 87781 59331 87847 59334
rect 90081 59331 90147 59334
rect 90357 59394 90423 59397
rect 91694 59394 91754 59606
rect 93393 59603 93459 59606
rect 94313 59603 94379 59606
rect 91921 59530 91987 59533
rect 93117 59530 93183 59533
rect 91921 59528 93183 59530
rect 91921 59472 91926 59528
rect 91982 59472 93122 59528
rect 93178 59472 93183 59528
rect 91921 59470 93183 59472
rect 91921 59467 91987 59470
rect 93117 59467 93183 59470
rect 93301 59530 93367 59533
rect 95729 59530 95789 60044
rect 95969 59666 96035 59669
rect 96560 59666 96620 60044
rect 95969 59664 96620 59666
rect 95969 59608 95974 59664
rect 96030 59608 96620 59664
rect 95969 59606 96620 59608
rect 96705 59666 96771 59669
rect 97392 59666 97452 60044
rect 96705 59664 97452 59666
rect 96705 59608 96710 59664
rect 96766 59608 97452 59664
rect 96705 59606 97452 59608
rect 95969 59603 96035 59606
rect 96705 59603 96771 59606
rect 93301 59528 95789 59530
rect 93301 59472 93306 59528
rect 93362 59472 95789 59528
rect 93301 59470 95789 59472
rect 95877 59530 95943 59533
rect 98224 59530 98284 60044
rect 98361 59802 98427 59805
rect 99055 59802 99115 60044
rect 98361 59800 99115 59802
rect 98361 59744 98366 59800
rect 98422 59744 99115 59800
rect 98361 59742 99115 59744
rect 98361 59739 98427 59742
rect 99887 59666 99947 60044
rect 100718 59938 100778 60044
rect 95877 59528 98284 59530
rect 95877 59472 95882 59528
rect 95938 59472 98284 59528
rect 95877 59470 98284 59472
rect 98502 59606 99947 59666
rect 100158 59878 100778 59938
rect 93301 59467 93367 59470
rect 95877 59467 95943 59470
rect 90357 59392 91754 59394
rect 90357 59336 90362 59392
rect 90418 59336 91754 59392
rect 90357 59334 91754 59336
rect 91829 59394 91895 59397
rect 94313 59394 94379 59397
rect 95969 59394 96035 59397
rect 91829 59392 94379 59394
rect 91829 59336 91834 59392
rect 91890 59336 94318 59392
rect 94374 59336 94379 59392
rect 91829 59334 94379 59336
rect 90357 59331 90423 59334
rect 91829 59331 91895 59334
rect 94313 59331 94379 59334
rect 95190 59392 96035 59394
rect 95190 59336 95974 59392
rect 96030 59336 96035 59392
rect 95190 59334 96035 59336
rect 93117 59258 93183 59261
rect 95190 59258 95250 59334
rect 95969 59331 96035 59334
rect 97257 59394 97323 59397
rect 98502 59394 98562 59606
rect 98821 59530 98887 59533
rect 100158 59530 100218 59878
rect 100845 59802 100911 59805
rect 101550 59802 101610 60044
rect 102382 59938 102442 60044
rect 100845 59800 101610 59802
rect 100845 59744 100850 59800
rect 100906 59744 101610 59800
rect 100845 59742 101610 59744
rect 101998 59878 102442 59938
rect 100845 59739 100911 59742
rect 101998 59666 102058 59878
rect 102501 59802 102567 59805
rect 103213 59802 103273 60044
rect 102501 59800 103273 59802
rect 102501 59744 102506 59800
rect 102562 59744 103273 59800
rect 102501 59742 103273 59744
rect 103421 59802 103487 59805
rect 104045 59802 104105 60044
rect 103421 59800 104105 59802
rect 103421 59744 103426 59800
rect 103482 59744 104105 59800
rect 103421 59742 104105 59744
rect 102501 59739 102567 59742
rect 103421 59739 103487 59742
rect 98821 59528 100218 59530
rect 98821 59472 98826 59528
rect 98882 59472 100218 59528
rect 98821 59470 100218 59472
rect 100342 59606 102058 59666
rect 102961 59666 103027 59669
rect 104876 59666 104936 60044
rect 102961 59664 104936 59666
rect 102961 59608 102966 59664
rect 103022 59608 104936 59664
rect 102961 59606 104936 59608
rect 105077 59666 105143 59669
rect 105708 59666 105768 60044
rect 105077 59664 105768 59666
rect 105077 59608 105082 59664
rect 105138 59608 105768 59664
rect 105077 59606 105768 59608
rect 98821 59467 98887 59470
rect 97257 59392 98562 59394
rect 97257 59336 97262 59392
rect 97318 59336 98562 59392
rect 97257 59334 98562 59336
rect 100017 59394 100083 59397
rect 100342 59394 100402 59606
rect 102961 59603 103027 59606
rect 105077 59603 105143 59606
rect 101397 59530 101463 59533
rect 103421 59530 103487 59533
rect 101397 59528 103487 59530
rect 101397 59472 101402 59528
rect 101458 59472 103426 59528
rect 103482 59472 103487 59528
rect 101397 59470 103487 59472
rect 101397 59467 101463 59470
rect 103421 59467 103487 59470
rect 104341 59530 104407 59533
rect 106540 59530 106600 60044
rect 107371 59938 107431 60044
rect 107334 59878 107431 59938
rect 107193 59802 107259 59805
rect 104341 59528 106600 59530
rect 104341 59472 104346 59528
rect 104402 59472 106600 59528
rect 104341 59470 106600 59472
rect 106782 59800 107259 59802
rect 106782 59744 107198 59800
rect 107254 59744 107259 59800
rect 106782 59742 107259 59744
rect 104341 59467 104407 59470
rect 102501 59394 102567 59397
rect 100017 59392 100402 59394
rect 100017 59336 100022 59392
rect 100078 59336 100402 59392
rect 100017 59334 100402 59336
rect 101078 59392 102567 59394
rect 101078 59336 102506 59392
rect 102562 59336 102567 59392
rect 101078 59334 102567 59336
rect 97257 59331 97323 59334
rect 100017 59331 100083 59334
rect 93117 59256 95250 59258
rect 93117 59200 93122 59256
rect 93178 59200 95250 59256
rect 93117 59198 95250 59200
rect 100201 59258 100267 59261
rect 101078 59258 101138 59334
rect 102501 59331 102567 59334
rect 104157 59394 104223 59397
rect 105537 59394 105603 59397
rect 106782 59394 106842 59742
rect 107193 59739 107259 59742
rect 107334 59530 107394 59878
rect 107469 59802 107535 59805
rect 108203 59802 108263 60044
rect 107469 59800 108263 59802
rect 107469 59744 107474 59800
rect 107530 59744 108263 59800
rect 107469 59742 108263 59744
rect 107469 59739 107535 59742
rect 107561 59666 107627 59669
rect 109034 59666 109094 60044
rect 107561 59664 109094 59666
rect 107561 59608 107566 59664
rect 107622 59608 109094 59664
rect 107561 59606 109094 59608
rect 109217 59666 109283 59669
rect 109866 59666 109926 60044
rect 109217 59664 109926 59666
rect 109217 59608 109222 59664
rect 109278 59608 109926 59664
rect 109217 59606 109926 59608
rect 107561 59603 107627 59606
rect 109217 59603 109283 59606
rect 104157 59392 105370 59394
rect 104157 59336 104162 59392
rect 104218 59336 105370 59392
rect 104157 59334 105370 59336
rect 104157 59331 104223 59334
rect 100201 59256 101138 59258
rect 100201 59200 100206 59256
rect 100262 59200 101138 59256
rect 100201 59198 101138 59200
rect 105310 59258 105370 59334
rect 105537 59392 106842 59394
rect 105537 59336 105542 59392
rect 105598 59336 106842 59392
rect 105537 59334 106842 59336
rect 106966 59470 107394 59530
rect 108481 59530 108547 59533
rect 110698 59530 110758 60044
rect 110873 59666 110939 59669
rect 111529 59666 111589 60044
rect 111793 59802 111859 59805
rect 112361 59802 112421 60044
rect 111793 59800 112421 59802
rect 111793 59744 111798 59800
rect 111854 59744 112421 59800
rect 111793 59742 112421 59744
rect 111793 59739 111859 59742
rect 110873 59664 111589 59666
rect 110873 59608 110878 59664
rect 110934 59608 111589 59664
rect 110873 59606 111589 59608
rect 111701 59666 111767 59669
rect 113192 59666 113252 60044
rect 111701 59664 113252 59666
rect 111701 59608 111706 59664
rect 111762 59608 113252 59664
rect 111701 59606 113252 59608
rect 113541 59666 113607 59669
rect 114024 59666 114084 60044
rect 113541 59664 114084 59666
rect 113541 59608 113546 59664
rect 113602 59608 114084 59664
rect 113541 59606 114084 59608
rect 110873 59603 110939 59606
rect 111701 59603 111767 59606
rect 113541 59603 113607 59606
rect 111793 59530 111859 59533
rect 108481 59528 110758 59530
rect 108481 59472 108486 59528
rect 108542 59472 110758 59528
rect 108481 59470 110758 59472
rect 110830 59528 111859 59530
rect 110830 59472 111798 59528
rect 111854 59472 111859 59528
rect 110830 59470 111859 59472
rect 105537 59331 105603 59334
rect 106966 59258 107026 59470
rect 108481 59467 108547 59470
rect 107101 59394 107167 59397
rect 108849 59394 108915 59397
rect 107101 59392 108915 59394
rect 107101 59336 107106 59392
rect 107162 59336 108854 59392
rect 108910 59336 108915 59392
rect 107101 59334 108915 59336
rect 107101 59331 107167 59334
rect 108849 59331 108915 59334
rect 109033 59394 109099 59397
rect 110830 59394 110890 59470
rect 111793 59467 111859 59470
rect 112989 59530 113055 59533
rect 114856 59530 114916 60044
rect 115013 59802 115079 59805
rect 115687 59802 115747 60044
rect 115013 59800 115747 59802
rect 115013 59744 115018 59800
rect 115074 59744 115747 59800
rect 115013 59742 115747 59744
rect 115013 59739 115079 59742
rect 116519 59666 116579 60044
rect 112989 59528 114916 59530
rect 112989 59472 112994 59528
rect 113050 59472 114916 59528
rect 112989 59470 114916 59472
rect 115062 59606 116579 59666
rect 112989 59467 113055 59470
rect 109033 59392 110890 59394
rect 109033 59336 109038 59392
rect 109094 59336 110890 59392
rect 109033 59334 110890 59336
rect 111609 59394 111675 59397
rect 113541 59394 113607 59397
rect 111609 59392 113607 59394
rect 111609 59336 111614 59392
rect 111670 59336 113546 59392
rect 113602 59336 113607 59392
rect 111609 59334 113607 59336
rect 109033 59331 109099 59334
rect 111609 59331 111675 59334
rect 113541 59331 113607 59334
rect 114185 59394 114251 59397
rect 115062 59394 115122 59606
rect 115197 59530 115263 59533
rect 117350 59530 117410 60044
rect 115197 59528 117410 59530
rect 115197 59472 115202 59528
rect 115258 59472 117410 59528
rect 115197 59470 117410 59472
rect 117497 59530 117563 59533
rect 118182 59530 118242 60044
rect 117497 59528 118242 59530
rect 117497 59472 117502 59528
rect 117558 59472 118242 59528
rect 117497 59470 118242 59472
rect 115197 59467 115263 59470
rect 117497 59467 117563 59470
rect 114185 59392 115122 59394
rect 114185 59336 114190 59392
rect 114246 59336 115122 59392
rect 114185 59334 115122 59336
rect 116577 59394 116643 59397
rect 119014 59394 119074 60044
rect 119845 59938 119905 60044
rect 120677 59938 120737 60044
rect 119845 59878 119906 59938
rect 119846 59768 119906 59878
rect 119845 59708 119906 59768
rect 120030 59878 120737 59938
rect 119845 59530 119905 59708
rect 120030 59669 120090 59878
rect 121508 59802 121568 60044
rect 119981 59664 120090 59669
rect 119981 59608 119986 59664
rect 120042 59608 120090 59664
rect 119981 59606 120090 59608
rect 120214 59742 121568 59802
rect 121637 59802 121703 59805
rect 122340 59802 122400 60044
rect 121637 59800 122400 59802
rect 121637 59744 121642 59800
rect 121698 59744 122400 59800
rect 121637 59742 122400 59744
rect 119981 59603 120047 59606
rect 116577 59392 119074 59394
rect 116577 59336 116582 59392
rect 116638 59336 119074 59392
rect 116577 59334 119074 59336
rect 119294 59470 119905 59530
rect 119981 59530 120047 59533
rect 120214 59530 120274 59742
rect 121637 59739 121703 59742
rect 120717 59666 120783 59669
rect 122741 59666 122807 59669
rect 120717 59664 122807 59666
rect 120717 59608 120722 59664
rect 120778 59608 122746 59664
rect 122802 59608 122807 59664
rect 120717 59606 122807 59608
rect 120717 59603 120783 59606
rect 122741 59603 122807 59606
rect 119981 59528 120274 59530
rect 119981 59472 119986 59528
rect 120042 59472 120274 59528
rect 119981 59470 120274 59472
rect 120901 59530 120967 59533
rect 123172 59530 123232 60044
rect 123293 59802 123359 59805
rect 124003 59802 124063 60044
rect 123293 59800 124063 59802
rect 123293 59744 123298 59800
rect 123354 59744 124063 59800
rect 123293 59742 124063 59744
rect 124213 59802 124279 59805
rect 124835 59802 124895 60044
rect 124213 59800 124895 59802
rect 124213 59744 124218 59800
rect 124274 59744 124895 59800
rect 124213 59742 124895 59744
rect 123293 59739 123359 59742
rect 124213 59739 124279 59742
rect 123477 59666 123543 59669
rect 125666 59666 125726 60044
rect 123477 59664 125726 59666
rect 123477 59608 123482 59664
rect 123538 59608 125726 59664
rect 123477 59606 125726 59608
rect 125869 59666 125935 59669
rect 126498 59666 126558 60044
rect 125869 59664 126558 59666
rect 125869 59608 125874 59664
rect 125930 59608 126558 59664
rect 125869 59606 126558 59608
rect 123477 59603 123543 59606
rect 125869 59603 125935 59606
rect 120901 59528 123232 59530
rect 120901 59472 120906 59528
rect 120962 59472 123232 59528
rect 120901 59470 123232 59472
rect 125041 59530 125107 59533
rect 127330 59530 127390 60044
rect 128161 59938 128221 60044
rect 127574 59878 128221 59938
rect 127574 59805 127634 59878
rect 127525 59800 127634 59805
rect 128993 59802 129053 60044
rect 127525 59744 127530 59800
rect 127586 59744 127634 59800
rect 128310 59768 129053 59802
rect 127525 59742 127634 59744
rect 128126 59742 129053 59768
rect 127525 59739 127591 59742
rect 128126 59708 128370 59742
rect 128126 59530 128186 59708
rect 125041 59528 127390 59530
rect 125041 59472 125046 59528
rect 125102 59472 127390 59528
rect 125041 59470 127390 59472
rect 127574 59470 128186 59530
rect 128353 59530 128419 59533
rect 129824 59530 129884 60044
rect 128353 59528 129884 59530
rect 128353 59472 128358 59528
rect 128414 59472 129884 59528
rect 128353 59470 129884 59472
rect 114185 59331 114251 59334
rect 116577 59331 116643 59334
rect 105310 59198 107026 59258
rect 116761 59258 116827 59261
rect 119294 59258 119354 59470
rect 119981 59467 120047 59470
rect 120901 59467 120967 59470
rect 125041 59467 125107 59470
rect 119521 59394 119587 59397
rect 121637 59394 121703 59397
rect 119521 59392 121703 59394
rect 119521 59336 119526 59392
rect 119582 59336 121642 59392
rect 121698 59336 121703 59392
rect 119521 59334 121703 59336
rect 119521 59331 119587 59334
rect 121637 59331 121703 59334
rect 122097 59394 122163 59397
rect 124213 59394 124279 59397
rect 125869 59394 125935 59397
rect 122097 59392 124279 59394
rect 122097 59336 122102 59392
rect 122158 59336 124218 59392
rect 124274 59336 124279 59392
rect 122097 59334 124279 59336
rect 122097 59331 122163 59334
rect 124213 59331 124279 59334
rect 124998 59392 125935 59394
rect 124998 59336 125874 59392
rect 125930 59336 125935 59392
rect 124998 59334 125935 59336
rect 116761 59256 119354 59258
rect 116761 59200 116766 59256
rect 116822 59200 119354 59256
rect 116761 59198 119354 59200
rect 123661 59258 123727 59261
rect 124998 59258 125058 59334
rect 125869 59331 125935 59334
rect 126237 59394 126303 59397
rect 127574 59394 127634 59470
rect 128353 59467 128419 59470
rect 126237 59392 127634 59394
rect 126237 59336 126242 59392
rect 126298 59336 127634 59392
rect 126237 59334 127634 59336
rect 127709 59394 127775 59397
rect 130656 59394 130716 60044
rect 131488 59394 131548 60044
rect 131665 59666 131731 59669
rect 132319 59666 132379 60044
rect 133151 59938 133211 60044
rect 133982 59938 134042 60044
rect 131665 59664 132379 59666
rect 131665 59608 131670 59664
rect 131726 59608 132379 59664
rect 131665 59606 132379 59608
rect 132542 59878 133211 59938
rect 133278 59878 134042 59938
rect 131665 59603 131731 59606
rect 132542 59530 132602 59878
rect 133278 59666 133338 59878
rect 127709 59392 130716 59394
rect 127709 59336 127714 59392
rect 127770 59336 130716 59392
rect 127709 59334 130716 59336
rect 130886 59334 131548 59394
rect 131622 59470 132602 59530
rect 132726 59606 133338 59666
rect 134149 59666 134215 59669
rect 134814 59666 134874 60044
rect 134149 59664 134874 59666
rect 134149 59608 134154 59664
rect 134210 59608 134874 59664
rect 134149 59606 134874 59608
rect 126237 59331 126303 59334
rect 127709 59331 127775 59334
rect 123661 59256 125058 59258
rect 123661 59200 123666 59256
rect 123722 59200 125058 59256
rect 123661 59198 125058 59200
rect 129181 59258 129247 59261
rect 130886 59258 130946 59334
rect 129181 59256 130946 59258
rect 129181 59200 129186 59256
rect 129242 59200 130946 59256
rect 129181 59198 130946 59200
rect 93117 59195 93183 59198
rect 100201 59195 100267 59198
rect 116761 59195 116827 59198
rect 123661 59195 123727 59198
rect 129181 59195 129247 59198
rect 72417 59120 73722 59122
rect 72417 59064 72422 59120
rect 72478 59064 73722 59120
rect 72417 59062 73722 59064
rect 130377 59122 130443 59125
rect 131622 59122 131682 59470
rect 131849 59394 131915 59397
rect 132726 59394 132786 59606
rect 134149 59603 134215 59606
rect 133137 59530 133203 59533
rect 135646 59530 135706 60044
rect 133137 59528 135706 59530
rect 133137 59472 133142 59528
rect 133198 59472 135706 59528
rect 133137 59470 135706 59472
rect 133137 59467 133203 59470
rect 131849 59392 132786 59394
rect 131849 59336 131854 59392
rect 131910 59336 132786 59392
rect 131849 59334 132786 59336
rect 133413 59394 133479 59397
rect 136477 59394 136537 60044
rect 136633 59802 136699 59805
rect 137309 59802 137369 60044
rect 136633 59800 137369 59802
rect 136633 59744 136638 59800
rect 136694 59744 137369 59800
rect 136633 59742 137369 59744
rect 136633 59739 136699 59742
rect 136633 59666 136699 59669
rect 138140 59666 138200 60044
rect 136633 59664 138200 59666
rect 136633 59608 136638 59664
rect 136694 59608 138200 59664
rect 136633 59606 138200 59608
rect 138473 59666 138539 59669
rect 138972 59666 139032 60044
rect 139209 59802 139275 59805
rect 139804 59802 139864 60044
rect 139209 59800 139864 59802
rect 139209 59744 139214 59800
rect 139270 59744 139864 59800
rect 139209 59742 139864 59744
rect 139945 59802 140011 59805
rect 140635 59802 140695 60044
rect 139945 59800 140695 59802
rect 139945 59744 139950 59800
rect 140006 59744 140695 59800
rect 139945 59742 140695 59744
rect 139209 59739 139275 59742
rect 139945 59739 140011 59742
rect 138473 59664 139032 59666
rect 138473 59608 138478 59664
rect 138534 59608 139032 59664
rect 138473 59606 139032 59608
rect 139117 59666 139183 59669
rect 141467 59666 141527 60044
rect 141693 59802 141759 59805
rect 142298 59802 142358 60044
rect 143130 59938 143190 60044
rect 143962 59938 144022 60044
rect 144793 59938 144853 60044
rect 142478 59878 143190 59938
rect 143398 59878 144022 59938
rect 144134 59878 144853 59938
rect 142478 59805 142538 59878
rect 141693 59800 142358 59802
rect 141693 59744 141698 59800
rect 141754 59744 142358 59800
rect 141693 59742 142358 59744
rect 142429 59800 142538 59805
rect 142429 59744 142434 59800
rect 142490 59744 142538 59800
rect 142429 59742 142538 59744
rect 141693 59739 141759 59742
rect 142429 59739 142495 59742
rect 139117 59664 139410 59666
rect 139117 59608 139122 59664
rect 139178 59608 139410 59664
rect 139117 59606 139410 59608
rect 136633 59603 136699 59606
rect 138473 59603 138539 59606
rect 139117 59603 139183 59606
rect 137461 59530 137527 59533
rect 139209 59530 139275 59533
rect 137461 59528 139275 59530
rect 137461 59472 137466 59528
rect 137522 59472 139214 59528
rect 139270 59472 139275 59528
rect 137461 59470 139275 59472
rect 139350 59530 139410 59606
rect 139902 59606 141527 59666
rect 141601 59666 141667 59669
rect 143398 59666 143458 59878
rect 144134 59804 144194 59878
rect 144126 59740 144132 59804
rect 144196 59740 144202 59804
rect 144269 59802 144335 59805
rect 145625 59802 145685 60044
rect 144269 59800 145685 59802
rect 144269 59744 144274 59800
rect 144330 59744 145685 59800
rect 144269 59742 145685 59744
rect 144269 59739 144335 59742
rect 141601 59664 143458 59666
rect 141601 59608 141606 59664
rect 141662 59608 143458 59664
rect 141601 59606 143458 59608
rect 144177 59666 144243 59669
rect 146456 59666 146516 60044
rect 144177 59664 146516 59666
rect 144177 59608 144182 59664
rect 144238 59608 146516 59664
rect 144177 59606 146516 59608
rect 146661 59666 146727 59669
rect 147288 59666 147348 60044
rect 146661 59664 147348 59666
rect 146661 59608 146666 59664
rect 146722 59608 147348 59664
rect 146661 59606 147348 59608
rect 147489 59666 147555 59669
rect 148120 59666 148180 60044
rect 147489 59664 148180 59666
rect 147489 59608 147494 59664
rect 147550 59608 148180 59664
rect 147489 59606 148180 59608
rect 139902 59530 139962 59606
rect 141601 59603 141667 59606
rect 144177 59603 144243 59606
rect 146661 59603 146727 59606
rect 147489 59603 147555 59606
rect 139350 59470 139962 59530
rect 140037 59530 140103 59533
rect 141693 59530 141759 59533
rect 140037 59528 141759 59530
rect 140037 59472 140042 59528
rect 140098 59472 141698 59528
rect 141754 59472 141759 59528
rect 140037 59470 141759 59472
rect 137461 59467 137527 59470
rect 139209 59467 139275 59470
rect 140037 59467 140103 59470
rect 141693 59467 141759 59470
rect 145557 59530 145623 59533
rect 148951 59530 149011 60044
rect 149783 59938 149843 60044
rect 149286 59878 149843 59938
rect 149145 59666 149211 59669
rect 149286 59666 149346 59878
rect 149421 59802 149487 59805
rect 150614 59802 150674 60044
rect 149421 59800 150674 59802
rect 149421 59744 149426 59800
rect 149482 59744 150674 59800
rect 149421 59742 150674 59744
rect 150801 59802 150867 59805
rect 151446 59802 151506 60044
rect 150801 59800 151506 59802
rect 150801 59744 150806 59800
rect 150862 59744 151506 59800
rect 150801 59742 151506 59744
rect 149421 59739 149487 59742
rect 150801 59739 150867 59742
rect 149145 59664 149346 59666
rect 149145 59608 149150 59664
rect 149206 59608 149346 59664
rect 149145 59606 149346 59608
rect 149697 59666 149763 59669
rect 151721 59666 151787 59669
rect 149697 59664 151787 59666
rect 149697 59608 149702 59664
rect 149758 59608 151726 59664
rect 151782 59608 151787 59664
rect 149697 59606 151787 59608
rect 149145 59603 149211 59606
rect 149697 59603 149763 59606
rect 151721 59603 151787 59606
rect 145557 59528 149011 59530
rect 145557 59472 145562 59528
rect 145618 59472 149011 59528
rect 145557 59470 149011 59472
rect 149881 59530 149947 59533
rect 152278 59530 152338 60044
rect 152457 59802 152523 59805
rect 153109 59802 153169 60044
rect 152457 59800 153169 59802
rect 152457 59744 152462 59800
rect 152518 59744 153169 59800
rect 152457 59742 153169 59744
rect 152457 59739 152523 59742
rect 153941 59666 154001 60044
rect 149881 59528 152338 59530
rect 149881 59472 149886 59528
rect 149942 59472 152338 59528
rect 149881 59470 152338 59472
rect 152782 59606 154001 59666
rect 145557 59467 145623 59470
rect 149881 59467 149947 59470
rect 133413 59392 136537 59394
rect 133413 59336 133418 59392
rect 133474 59336 136537 59392
rect 133413 59334 136537 59336
rect 137553 59394 137619 59397
rect 138473 59394 138539 59397
rect 139945 59394 140011 59397
rect 137553 59392 138539 59394
rect 137553 59336 137558 59392
rect 137614 59336 138478 59392
rect 138534 59336 138539 59392
rect 137553 59334 138539 59336
rect 131849 59331 131915 59334
rect 133413 59331 133479 59334
rect 137553 59331 137619 59334
rect 138473 59331 138539 59334
rect 139166 59392 140011 59394
rect 139166 59336 139950 59392
rect 140006 59336 140011 59392
rect 139166 59334 140011 59336
rect 137277 59258 137343 59261
rect 139166 59258 139226 59334
rect 139945 59331 140011 59334
rect 144361 59394 144427 59397
rect 146661 59394 146727 59397
rect 144361 59392 146727 59394
rect 144361 59336 144366 59392
rect 144422 59336 146666 59392
rect 146722 59336 146727 59392
rect 144361 59334 146727 59336
rect 144361 59331 144427 59334
rect 146661 59331 146727 59334
rect 148317 59394 148383 59397
rect 150249 59394 150315 59397
rect 148317 59392 150315 59394
rect 148317 59336 148322 59392
rect 148378 59336 150254 59392
rect 150310 59336 150315 59392
rect 148317 59334 150315 59336
rect 148317 59331 148383 59334
rect 150249 59331 150315 59334
rect 150433 59394 150499 59397
rect 152782 59394 152842 59606
rect 153101 59530 153167 59533
rect 154772 59530 154832 60044
rect 153101 59528 154832 59530
rect 153101 59472 153106 59528
rect 153162 59472 154832 59528
rect 153101 59470 154832 59472
rect 153101 59467 153167 59470
rect 150433 59392 152842 59394
rect 150433 59336 150438 59392
rect 150494 59336 152842 59392
rect 150433 59334 152842 59336
rect 153009 59394 153075 59397
rect 155604 59394 155664 60044
rect 156436 59530 156496 60044
rect 156597 59802 156663 59805
rect 157267 59802 157327 60044
rect 156597 59800 157327 59802
rect 156597 59744 156602 59800
rect 156658 59744 157327 59800
rect 156597 59742 157327 59744
rect 156597 59739 156663 59742
rect 156597 59666 156663 59669
rect 158099 59666 158159 60044
rect 158930 59938 158990 60044
rect 159762 59938 159822 60044
rect 156597 59664 158159 59666
rect 156597 59608 156602 59664
rect 156658 59608 158159 59664
rect 156597 59606 158159 59608
rect 158302 59878 158990 59938
rect 159222 59878 159822 59938
rect 156597 59603 156663 59606
rect 156965 59530 157031 59533
rect 156436 59528 157031 59530
rect 156436 59472 156970 59528
rect 157026 59472 157031 59528
rect 156436 59470 157031 59472
rect 156965 59467 157031 59470
rect 157241 59530 157307 59533
rect 158302 59530 158362 59878
rect 157241 59528 158362 59530
rect 157241 59472 157246 59528
rect 157302 59472 158362 59528
rect 157241 59470 158362 59472
rect 157241 59467 157307 59470
rect 153009 59392 155664 59394
rect 153009 59336 153014 59392
rect 153070 59336 155664 59392
rect 153009 59334 155664 59336
rect 155861 59394 155927 59397
rect 156597 59394 156663 59397
rect 155861 59392 156663 59394
rect 155861 59336 155866 59392
rect 155922 59336 156602 59392
rect 156658 59336 156663 59392
rect 155861 59334 156663 59336
rect 150433 59331 150499 59334
rect 153009 59331 153075 59334
rect 155861 59331 155927 59334
rect 156597 59331 156663 59334
rect 157333 59394 157399 59397
rect 159222 59394 159282 59878
rect 159909 59802 159975 59805
rect 160594 59802 160654 60044
rect 161425 59938 161485 60044
rect 162257 59938 162317 60044
rect 163088 59938 163148 60044
rect 160878 59878 161485 59938
rect 161798 59878 162317 59938
rect 162534 59878 163148 59938
rect 159909 59800 160654 59802
rect 159909 59744 159914 59800
rect 159970 59744 160654 59800
rect 159909 59742 160654 59744
rect 160737 59802 160803 59805
rect 160878 59802 160938 59878
rect 160737 59800 160938 59802
rect 160737 59744 160742 59800
rect 160798 59744 160938 59800
rect 160737 59742 160938 59744
rect 159909 59739 159975 59742
rect 160737 59739 160803 59742
rect 161798 59666 161858 59878
rect 160694 59606 161858 59666
rect 160001 59530 160067 59533
rect 160694 59530 160754 59606
rect 160001 59528 160754 59530
rect 160001 59472 160006 59528
rect 160062 59472 160754 59528
rect 160001 59470 160754 59472
rect 161105 59530 161171 59533
rect 162534 59530 162594 59878
rect 163920 59802 163980 60044
rect 161105 59528 162594 59530
rect 161105 59472 161110 59528
rect 161166 59472 162594 59528
rect 161105 59470 162594 59472
rect 162718 59742 163980 59802
rect 160001 59467 160067 59470
rect 161105 59467 161171 59470
rect 157333 59392 159282 59394
rect 157333 59336 157338 59392
rect 157394 59336 159282 59392
rect 157333 59334 159282 59336
rect 161289 59394 161355 59397
rect 162718 59394 162778 59742
rect 162853 59666 162919 59669
rect 164752 59666 164812 60044
rect 162853 59664 164812 59666
rect 162853 59608 162858 59664
rect 162914 59608 164812 59664
rect 162853 59606 164812 59608
rect 162853 59603 162919 59606
rect 163865 59530 163931 59533
rect 165583 59530 165643 60044
rect 163865 59528 165643 59530
rect 163865 59472 163870 59528
rect 163926 59472 165643 59528
rect 163865 59470 165643 59472
rect 163865 59467 163931 59470
rect 161289 59392 162778 59394
rect 161289 59336 161294 59392
rect 161350 59336 162778 59392
rect 161289 59334 162778 59336
rect 164049 59394 164115 59397
rect 166415 59394 166475 60044
rect 167246 59530 167306 60044
rect 167453 59802 167519 59805
rect 168078 59802 168138 60044
rect 167453 59800 168138 59802
rect 167453 59744 167458 59800
rect 167514 59744 168138 59800
rect 167453 59742 168138 59744
rect 167453 59739 167519 59742
rect 168910 59666 168970 60044
rect 164049 59392 166475 59394
rect 164049 59336 164054 59392
rect 164110 59336 166475 59392
rect 164049 59334 166475 59336
rect 166582 59470 167306 59530
rect 167502 59606 168970 59666
rect 157333 59331 157399 59334
rect 161289 59331 161355 59334
rect 164049 59331 164115 59334
rect 137277 59256 139226 59258
rect 137277 59200 137282 59256
rect 137338 59200 139226 59256
rect 137277 59198 139226 59200
rect 165429 59258 165495 59261
rect 166582 59258 166642 59470
rect 166901 59394 166967 59397
rect 167502 59394 167562 59606
rect 168281 59530 168347 59533
rect 169741 59530 169801 60044
rect 168281 59528 169801 59530
rect 168281 59472 168286 59528
rect 168342 59472 169801 59528
rect 168281 59470 169801 59472
rect 169937 59530 170003 59533
rect 170573 59530 170633 60044
rect 169937 59528 170633 59530
rect 169937 59472 169942 59528
rect 169998 59472 170633 59528
rect 169937 59470 170633 59472
rect 168281 59467 168347 59470
rect 169937 59467 170003 59470
rect 166901 59392 167562 59394
rect 166901 59336 166906 59392
rect 166962 59336 167562 59392
rect 166901 59334 167562 59336
rect 168097 59394 168163 59397
rect 169385 59394 169451 59397
rect 168097 59392 169451 59394
rect 168097 59336 168102 59392
rect 168158 59336 169390 59392
rect 169446 59336 169451 59392
rect 168097 59334 169451 59336
rect 166901 59331 166967 59334
rect 168097 59331 168163 59334
rect 169385 59331 169451 59334
rect 169569 59394 169635 59397
rect 171404 59394 171464 60044
rect 171593 59530 171659 59533
rect 172236 59530 172296 60044
rect 171593 59528 172296 59530
rect 171593 59472 171598 59528
rect 171654 59472 172296 59528
rect 171593 59470 172296 59472
rect 171593 59467 171659 59470
rect 173068 59394 173128 60044
rect 173899 59802 173959 60044
rect 174537 59802 174603 59805
rect 173899 59800 174603 59802
rect 173899 59744 174542 59800
rect 174598 59744 174603 59800
rect 173899 59742 174603 59744
rect 174537 59739 174603 59742
rect 174731 59666 174791 60044
rect 169569 59392 171464 59394
rect 169569 59336 169574 59392
rect 169630 59336 171464 59392
rect 169569 59334 171464 59336
rect 171550 59334 173128 59394
rect 173206 59606 174791 59666
rect 169569 59331 169635 59334
rect 165429 59256 166642 59258
rect 165429 59200 165434 59256
rect 165490 59200 166642 59256
rect 165429 59198 166642 59200
rect 171041 59258 171107 59261
rect 171550 59258 171610 59334
rect 171041 59256 171610 59258
rect 171041 59200 171046 59256
rect 171102 59200 171610 59256
rect 171041 59198 171610 59200
rect 172421 59258 172487 59261
rect 173206 59258 173266 59606
rect 173801 59530 173867 59533
rect 175562 59530 175622 60044
rect 175733 59802 175799 59805
rect 176394 59802 176454 60044
rect 175733 59800 176454 59802
rect 175733 59744 175738 59800
rect 175794 59744 176454 59800
rect 175733 59742 176454 59744
rect 175733 59739 175799 59742
rect 177226 59666 177286 60044
rect 173801 59528 175622 59530
rect 173801 59472 173806 59528
rect 173862 59472 175622 59528
rect 173801 59470 175622 59472
rect 175782 59606 177286 59666
rect 173801 59467 173867 59470
rect 175181 59394 175247 59397
rect 175782 59394 175842 59606
rect 176469 59530 176535 59533
rect 178057 59530 178117 60044
rect 176469 59528 178117 59530
rect 176469 59472 176474 59528
rect 176530 59472 178117 59528
rect 176469 59470 178117 59472
rect 178217 59530 178283 59533
rect 178889 59530 178949 60044
rect 178217 59528 178949 59530
rect 178217 59472 178222 59528
rect 178278 59472 178949 59528
rect 178217 59470 178949 59472
rect 176469 59467 176535 59470
rect 178217 59467 178283 59470
rect 175181 59392 175842 59394
rect 175181 59336 175186 59392
rect 175242 59336 175842 59392
rect 175181 59334 175842 59336
rect 177665 59394 177731 59397
rect 179720 59394 179780 60044
rect 180552 59394 180612 60044
rect 180701 59666 180767 59669
rect 181384 59666 181444 60044
rect 180701 59664 181444 59666
rect 180701 59608 180706 59664
rect 180762 59608 181444 59664
rect 180701 59606 181444 59608
rect 180701 59603 180767 59606
rect 180701 59530 180767 59533
rect 182215 59530 182275 60044
rect 182357 59802 182423 59805
rect 183047 59802 183107 60044
rect 183878 59938 183938 60044
rect 183326 59878 183938 59938
rect 182357 59800 183107 59802
rect 182357 59744 182362 59800
rect 182418 59744 183107 59800
rect 182357 59742 183107 59744
rect 183185 59802 183251 59805
rect 183326 59802 183386 59878
rect 183185 59800 183386 59802
rect 183185 59744 183190 59800
rect 183246 59744 183386 59800
rect 183185 59742 183386 59744
rect 182357 59739 182423 59742
rect 183185 59739 183251 59742
rect 182357 59666 182423 59669
rect 184710 59666 184770 60044
rect 182357 59664 184770 59666
rect 182357 59608 182362 59664
rect 182418 59608 184770 59664
rect 182357 59606 184770 59608
rect 182357 59603 182423 59606
rect 185542 59530 185602 60044
rect 185669 59802 185735 59805
rect 186373 59802 186433 60044
rect 185669 59800 186433 59802
rect 185669 59744 185674 59800
rect 185730 59744 186433 59800
rect 185669 59742 186433 59744
rect 185669 59739 185735 59742
rect 187205 59666 187265 60044
rect 187417 59802 187483 59805
rect 188036 59802 188096 60044
rect 187417 59800 188096 59802
rect 187417 59744 187422 59800
rect 187478 59744 188096 59800
rect 187417 59742 188096 59744
rect 187417 59739 187483 59742
rect 180701 59528 182275 59530
rect 180701 59472 180706 59528
rect 180762 59472 182275 59528
rect 180701 59470 182275 59472
rect 183694 59470 185602 59530
rect 185718 59606 187265 59666
rect 187325 59666 187391 59669
rect 188868 59666 188928 60044
rect 187325 59664 188928 59666
rect 187325 59608 187330 59664
rect 187386 59608 188928 59664
rect 187325 59606 188928 59608
rect 180701 59467 180767 59470
rect 177665 59392 179780 59394
rect 177665 59336 177670 59392
rect 177726 59336 179780 59392
rect 177665 59334 179780 59336
rect 180014 59334 180612 59394
rect 181805 59394 181871 59397
rect 183185 59394 183251 59397
rect 181805 59392 183251 59394
rect 181805 59336 181810 59392
rect 181866 59336 183190 59392
rect 183246 59336 183251 59392
rect 181805 59334 183251 59336
rect 175181 59331 175247 59334
rect 177665 59331 177731 59334
rect 172421 59256 173266 59258
rect 172421 59200 172426 59256
rect 172482 59200 173266 59256
rect 172421 59198 173266 59200
rect 177849 59258 177915 59261
rect 180014 59258 180074 59334
rect 181805 59331 181871 59334
rect 183185 59331 183251 59334
rect 177849 59256 180074 59258
rect 177849 59200 177854 59256
rect 177910 59200 180074 59256
rect 177849 59198 180074 59200
rect 183461 59258 183527 59261
rect 183694 59258 183754 59470
rect 185718 59394 185778 59606
rect 187325 59603 187391 59606
rect 186129 59530 186195 59533
rect 187417 59530 187483 59533
rect 186129 59528 187483 59530
rect 186129 59472 186134 59528
rect 186190 59472 187422 59528
rect 187478 59472 187483 59528
rect 186129 59470 187483 59472
rect 186129 59467 186195 59470
rect 187417 59467 187483 59470
rect 185166 59334 185778 59394
rect 185945 59394 186011 59397
rect 187325 59394 187391 59397
rect 185945 59392 187391 59394
rect 185945 59336 185950 59392
rect 186006 59336 187330 59392
rect 187386 59336 187391 59392
rect 185945 59334 187391 59336
rect 183461 59256 183754 59258
rect 183461 59200 183466 59256
rect 183522 59200 183754 59256
rect 183461 59198 183754 59200
rect 184749 59258 184815 59261
rect 185166 59258 185226 59334
rect 185945 59331 186011 59334
rect 187325 59331 187391 59334
rect 187601 59394 187667 59397
rect 189700 59394 189760 60044
rect 189901 59802 189967 59805
rect 190531 59802 190591 60044
rect 189901 59800 190591 59802
rect 189901 59744 189906 59800
rect 189962 59744 190591 59800
rect 189901 59742 190591 59744
rect 189901 59739 189967 59742
rect 191363 59666 191423 60044
rect 192194 59938 192254 60044
rect 187601 59392 189760 59394
rect 187601 59336 187606 59392
rect 187662 59336 189760 59392
rect 187601 59334 189760 59336
rect 189950 59606 191423 59666
rect 191606 59878 192254 59938
rect 187601 59331 187667 59334
rect 184749 59256 185226 59258
rect 184749 59200 184754 59256
rect 184810 59200 185226 59256
rect 184749 59198 185226 59200
rect 188889 59258 188955 59261
rect 189950 59258 190010 59606
rect 190085 59530 190151 59533
rect 191606 59530 191666 59878
rect 193026 59802 193086 60044
rect 192194 59742 193086 59802
rect 191741 59666 191807 59669
rect 192194 59666 192254 59742
rect 193858 59666 193918 60044
rect 191741 59664 192254 59666
rect 191741 59608 191746 59664
rect 191802 59608 192254 59664
rect 191741 59606 192254 59608
rect 192342 59606 193918 59666
rect 191741 59603 191807 59606
rect 190085 59528 191666 59530
rect 190085 59472 190090 59528
rect 190146 59472 191666 59528
rect 190085 59470 191666 59472
rect 190085 59467 190151 59470
rect 190269 59394 190335 59397
rect 191557 59394 191623 59397
rect 190269 59392 191623 59394
rect 190269 59336 190274 59392
rect 190330 59336 191562 59392
rect 191618 59336 191623 59392
rect 190269 59334 191623 59336
rect 190269 59331 190335 59334
rect 191557 59331 191623 59334
rect 191741 59394 191807 59397
rect 192342 59394 192402 59606
rect 193029 59530 193095 59533
rect 194689 59530 194749 60044
rect 193029 59528 194749 59530
rect 193029 59472 193034 59528
rect 193090 59472 194749 59528
rect 193029 59470 194749 59472
rect 194869 59530 194935 59533
rect 195521 59530 195581 60044
rect 194869 59528 195581 59530
rect 194869 59472 194874 59528
rect 194930 59472 195581 59528
rect 194869 59470 195581 59472
rect 193029 59467 193095 59470
rect 194869 59467 194935 59470
rect 191741 59392 192402 59394
rect 191741 59336 191746 59392
rect 191802 59336 192402 59392
rect 191741 59334 192402 59336
rect 192845 59394 192911 59397
rect 194317 59394 194383 59397
rect 192845 59392 194383 59394
rect 192845 59336 192850 59392
rect 192906 59336 194322 59392
rect 194378 59336 194383 59392
rect 192845 59334 194383 59336
rect 191741 59331 191807 59334
rect 192845 59331 192911 59334
rect 194317 59331 194383 59334
rect 194501 59394 194567 59397
rect 196352 59394 196412 60044
rect 196525 59802 196591 59805
rect 197184 59802 197244 60044
rect 196525 59800 197244 59802
rect 196525 59744 196530 59800
rect 196586 59744 197244 59800
rect 196525 59742 197244 59744
rect 196525 59739 196591 59742
rect 198016 59666 198076 60044
rect 194501 59392 196412 59394
rect 194501 59336 194506 59392
rect 194562 59336 196412 59392
rect 194501 59334 196412 59336
rect 196574 59606 198076 59666
rect 194501 59331 194567 59334
rect 188889 59256 190010 59258
rect 188889 59200 188894 59256
rect 188950 59200 190010 59256
rect 188889 59198 190010 59200
rect 195881 59258 195947 59261
rect 196574 59258 196634 59606
rect 197169 59530 197235 59533
rect 198847 59530 198907 60044
rect 197169 59528 198907 59530
rect 197169 59472 197174 59528
rect 197230 59472 198907 59528
rect 197169 59470 198907 59472
rect 197169 59467 197235 59470
rect 196985 59394 197051 59397
rect 199679 59394 199739 60044
rect 200510 59394 200570 60044
rect 200665 59666 200731 59669
rect 201342 59666 201402 60044
rect 201493 59802 201559 59805
rect 202174 59802 202234 60044
rect 201493 59800 202234 59802
rect 201493 59744 201498 59800
rect 201554 59744 202234 59800
rect 201493 59742 202234 59744
rect 201493 59739 201559 59742
rect 203005 59666 203065 60044
rect 200665 59664 201402 59666
rect 200665 59608 200670 59664
rect 200726 59608 201402 59664
rect 200665 59606 201402 59608
rect 201542 59606 203065 59666
rect 203149 59666 203215 59669
rect 203837 59666 203897 60044
rect 203149 59664 203897 59666
rect 203149 59608 203154 59664
rect 203210 59608 203897 59664
rect 203149 59606 203897 59608
rect 200665 59603 200731 59606
rect 201125 59530 201191 59533
rect 201542 59530 201602 59606
rect 203149 59603 203215 59606
rect 201125 59528 201602 59530
rect 201125 59472 201130 59528
rect 201186 59472 201602 59528
rect 201125 59470 201602 59472
rect 202505 59530 202571 59533
rect 204668 59530 204728 60044
rect 205500 59938 205560 60044
rect 204854 59878 205560 59938
rect 204854 59805 204914 59878
rect 204805 59800 204914 59805
rect 204805 59744 204810 59800
rect 204866 59744 204914 59800
rect 204805 59742 204914 59744
rect 204805 59739 204871 59742
rect 206332 59666 206392 60044
rect 207163 59938 207223 60044
rect 202505 59528 204728 59530
rect 202505 59472 202510 59528
rect 202566 59472 204728 59528
rect 202505 59470 204728 59472
rect 204854 59606 206392 59666
rect 206510 59878 207223 59938
rect 201125 59467 201191 59470
rect 202505 59467 202571 59470
rect 201493 59394 201559 59397
rect 203149 59394 203215 59397
rect 196985 59392 199739 59394
rect 196985 59336 196990 59392
rect 197046 59336 199739 59392
rect 196985 59334 199739 59336
rect 199886 59334 200570 59394
rect 200806 59392 201559 59394
rect 200806 59336 201498 59392
rect 201554 59336 201559 59392
rect 200806 59334 201559 59336
rect 196985 59331 197051 59334
rect 195881 59256 196634 59258
rect 195881 59200 195886 59256
rect 195942 59200 196634 59256
rect 195881 59198 196634 59200
rect 198365 59258 198431 59261
rect 199886 59258 199946 59334
rect 198365 59256 199946 59258
rect 198365 59200 198370 59256
rect 198426 59200 199946 59256
rect 198365 59198 199946 59200
rect 200021 59258 200087 59261
rect 200806 59258 200866 59334
rect 201493 59331 201559 59334
rect 202462 59392 203215 59394
rect 202462 59336 203154 59392
rect 203210 59336 203215 59392
rect 202462 59334 203215 59336
rect 200021 59256 200866 59258
rect 200021 59200 200026 59256
rect 200082 59200 200866 59256
rect 200021 59198 200866 59200
rect 201309 59258 201375 59261
rect 202462 59258 202522 59334
rect 203149 59331 203215 59334
rect 204161 59394 204227 59397
rect 204854 59394 204914 59606
rect 205449 59530 205515 59533
rect 206510 59530 206570 59878
rect 205449 59528 206570 59530
rect 205449 59472 205454 59528
rect 205510 59472 206570 59528
rect 205449 59470 206570 59472
rect 207289 59530 207355 59533
rect 207995 59530 208055 60044
rect 207289 59528 208055 59530
rect 207289 59472 207294 59528
rect 207350 59472 208055 59528
rect 207289 59470 208055 59472
rect 205449 59467 205515 59470
rect 207289 59467 207355 59470
rect 204161 59392 204914 59394
rect 204161 59336 204166 59392
rect 204222 59336 204914 59392
rect 204161 59334 204914 59336
rect 206645 59394 206711 59397
rect 208826 59394 208886 60044
rect 209658 59802 209718 60044
rect 206645 59392 208886 59394
rect 206645 59336 206650 59392
rect 206706 59336 208886 59392
rect 206645 59334 208886 59336
rect 209086 59742 209718 59802
rect 204161 59331 204227 59334
rect 206645 59331 206711 59334
rect 201309 59256 202522 59258
rect 201309 59200 201314 59256
rect 201370 59200 202522 59256
rect 201309 59198 202522 59200
rect 206829 59258 206895 59261
rect 209086 59258 209146 59742
rect 210490 59666 210550 60044
rect 209730 59606 210550 59666
rect 210693 59666 210759 59669
rect 211321 59666 211381 60044
rect 210693 59664 211381 59666
rect 210693 59608 210698 59664
rect 210754 59608 211381 59664
rect 210693 59606 211381 59608
rect 209730 59530 209790 59606
rect 210693 59603 210759 59606
rect 206829 59256 209146 59258
rect 206829 59200 206834 59256
rect 206890 59200 209146 59256
rect 206829 59198 209146 59200
rect 209270 59470 209790 59530
rect 209865 59530 209931 59533
rect 212153 59530 212213 60044
rect 209865 59528 212213 59530
rect 209865 59472 209870 59528
rect 209926 59472 212213 59528
rect 209865 59470 212213 59472
rect 137277 59195 137343 59198
rect 165429 59195 165495 59198
rect 171041 59195 171107 59198
rect 172421 59195 172487 59198
rect 177849 59195 177915 59198
rect 183461 59195 183527 59198
rect 184749 59195 184815 59198
rect 188889 59195 188955 59198
rect 195881 59195 195947 59198
rect 198365 59195 198431 59198
rect 200021 59195 200087 59198
rect 201309 59195 201375 59198
rect 206829 59195 206895 59198
rect 130377 59120 131682 59122
rect 130377 59064 130382 59120
rect 130438 59064 131682 59120
rect 130377 59062 131682 59064
rect 208301 59122 208367 59125
rect 209270 59122 209330 59470
rect 209865 59467 209931 59470
rect 209589 59394 209655 59397
rect 210693 59394 210759 59397
rect 209589 59392 210759 59394
rect 209589 59336 209594 59392
rect 209650 59336 210698 59392
rect 210754 59336 210759 59392
rect 209589 59334 210759 59336
rect 209589 59331 209655 59334
rect 210693 59331 210759 59334
rect 210969 59394 211035 59397
rect 212984 59394 213044 60044
rect 213177 59802 213243 59805
rect 213816 59802 213876 60044
rect 213177 59800 213876 59802
rect 213177 59744 213182 59800
rect 213238 59744 213876 59800
rect 213177 59742 213876 59744
rect 214005 59802 214071 59805
rect 214648 59802 214708 60044
rect 214005 59800 214708 59802
rect 214005 59744 214010 59800
rect 214066 59744 214708 59800
rect 214005 59742 214708 59744
rect 213177 59739 213243 59742
rect 214005 59739 214071 59742
rect 213545 59666 213611 59669
rect 215479 59666 215539 60044
rect 213545 59664 215539 59666
rect 213545 59608 213550 59664
rect 213606 59608 215539 59664
rect 213545 59606 215539 59608
rect 215753 59666 215819 59669
rect 216311 59666 216371 60044
rect 215753 59664 216371 59666
rect 215753 59608 215758 59664
rect 215814 59608 216371 59664
rect 215753 59606 216371 59608
rect 213545 59603 213611 59606
rect 215753 59603 215819 59606
rect 214925 59530 214991 59533
rect 217142 59530 217202 60044
rect 214925 59528 217202 59530
rect 214925 59472 214930 59528
rect 214986 59472 217202 59528
rect 214925 59470 217202 59472
rect 214925 59467 214991 59470
rect 214005 59394 214071 59397
rect 215753 59394 215819 59397
rect 210969 59392 213044 59394
rect 210969 59336 210974 59392
rect 211030 59336 213044 59392
rect 210969 59334 213044 59336
rect 213134 59392 214071 59394
rect 213134 59336 214010 59392
rect 214066 59336 214071 59392
rect 213134 59334 214071 59336
rect 210969 59331 211035 59334
rect 212441 59258 212507 59261
rect 213134 59258 213194 59334
rect 214005 59331 214071 59334
rect 214790 59392 215819 59394
rect 214790 59336 215758 59392
rect 215814 59336 215819 59392
rect 214790 59334 215819 59336
rect 212441 59256 213194 59258
rect 212441 59200 212446 59256
rect 212502 59200 213194 59256
rect 212441 59198 213194 59200
rect 213729 59258 213795 59261
rect 214790 59258 214850 59334
rect 215753 59331 215819 59334
rect 215937 59394 216003 59397
rect 217974 59394 218034 60044
rect 218145 59802 218211 59805
rect 218806 59802 218866 60044
rect 218145 59800 218866 59802
rect 218145 59744 218150 59800
rect 218206 59744 218866 59800
rect 218145 59742 218866 59744
rect 218145 59739 218211 59742
rect 219637 59666 219697 60044
rect 215937 59392 218034 59394
rect 215937 59336 215942 59392
rect 215998 59336 218034 59392
rect 215937 59334 218034 59336
rect 218102 59606 219697 59666
rect 219801 59666 219867 59669
rect 220469 59666 220529 60044
rect 219801 59664 220529 59666
rect 219801 59608 219806 59664
rect 219862 59608 220529 59664
rect 219801 59606 220529 59608
rect 215937 59331 216003 59334
rect 213729 59256 214850 59258
rect 213729 59200 213734 59256
rect 213790 59200 214850 59256
rect 213729 59198 214850 59200
rect 217869 59258 217935 59261
rect 218102 59258 218162 59606
rect 219801 59603 219867 59606
rect 219065 59530 219131 59533
rect 221300 59530 221360 60044
rect 221457 59802 221523 59805
rect 222132 59802 222192 60044
rect 221457 59800 222192 59802
rect 221457 59744 221462 59800
rect 221518 59744 222192 59800
rect 221457 59742 222192 59744
rect 221457 59739 221523 59742
rect 222964 59666 223024 60044
rect 219065 59528 221360 59530
rect 219065 59472 219070 59528
rect 219126 59472 221360 59528
rect 219065 59470 221360 59472
rect 221598 59606 223024 59666
rect 219065 59467 219131 59470
rect 219801 59394 219867 59397
rect 217869 59256 218162 59258
rect 217869 59200 217874 59256
rect 217930 59200 218162 59256
rect 217869 59198 218162 59200
rect 218286 59392 219867 59394
rect 218286 59336 219806 59392
rect 219862 59336 219867 59392
rect 218286 59334 219867 59336
rect 212441 59195 212507 59198
rect 213729 59195 213795 59198
rect 217869 59195 217935 59198
rect 208301 59120 209330 59122
rect 208301 59064 208306 59120
rect 208362 59064 209330 59120
rect 208301 59062 209330 59064
rect 217685 59122 217751 59125
rect 218286 59122 218346 59334
rect 219801 59331 219867 59334
rect 220721 59394 220787 59397
rect 221598 59394 221658 59606
rect 222101 59530 222167 59533
rect 223795 59530 223855 60044
rect 222101 59528 223855 59530
rect 222101 59472 222106 59528
rect 222162 59472 223855 59528
rect 222101 59470 223855 59472
rect 222101 59467 222167 59470
rect 220721 59392 221658 59394
rect 220721 59336 220726 59392
rect 220782 59336 221658 59392
rect 220721 59334 221658 59336
rect 222009 59394 222075 59397
rect 224627 59394 224687 60044
rect 225458 59938 225518 60044
rect 225094 59878 225518 59938
rect 224953 59666 225019 59669
rect 225094 59666 225154 59878
rect 225229 59802 225295 59805
rect 226290 59802 226350 60044
rect 225229 59800 226350 59802
rect 225229 59744 225234 59800
rect 225290 59744 226350 59800
rect 225229 59742 226350 59744
rect 225229 59739 225295 59742
rect 227122 59666 227182 60044
rect 224953 59664 225154 59666
rect 224953 59608 224958 59664
rect 225014 59608 225154 59664
rect 224953 59606 225154 59608
rect 225462 59606 227182 59666
rect 224953 59603 225019 59606
rect 224769 59530 224835 59533
rect 225462 59530 225522 59606
rect 224769 59528 225522 59530
rect 224769 59472 224774 59528
rect 224830 59472 225522 59528
rect 224769 59470 225522 59472
rect 226149 59530 226215 59533
rect 227953 59530 228013 60044
rect 226149 59528 228013 59530
rect 226149 59472 226154 59528
rect 226210 59472 228013 59528
rect 226149 59470 228013 59472
rect 224769 59467 224835 59470
rect 226149 59467 226215 59470
rect 224953 59394 225019 59397
rect 222009 59392 224687 59394
rect 222009 59336 222014 59392
rect 222070 59336 224687 59392
rect 222009 59334 224687 59336
rect 224910 59392 225019 59394
rect 224910 59336 224958 59392
rect 225014 59336 225019 59392
rect 220721 59331 220787 59334
rect 222009 59331 222075 59334
rect 224910 59331 225019 59336
rect 225965 59394 226031 59397
rect 228785 59394 228845 60044
rect 228909 59666 228975 59669
rect 229616 59666 229676 60044
rect 228909 59664 229676 59666
rect 228909 59608 228914 59664
rect 228970 59608 229676 59664
rect 228909 59606 229676 59608
rect 228909 59603 228975 59606
rect 229001 59530 229067 59533
rect 230448 59530 230508 60044
rect 229001 59528 230508 59530
rect 229001 59472 229006 59528
rect 229062 59472 230508 59528
rect 229001 59470 230508 59472
rect 229001 59467 229067 59470
rect 225965 59392 228845 59394
rect 225965 59336 225970 59392
rect 226026 59336 228845 59392
rect 225965 59334 228845 59336
rect 228909 59394 228975 59397
rect 231280 59394 231340 60044
rect 232111 59802 232171 60044
rect 232773 59802 232839 59805
rect 232111 59800 232839 59802
rect 232111 59744 232778 59800
rect 232834 59744 232839 59800
rect 232111 59742 232839 59744
rect 232773 59739 232839 59742
rect 232943 59666 233003 60044
rect 228909 59392 231340 59394
rect 228909 59336 228914 59392
rect 228970 59336 231340 59392
rect 228909 59334 231340 59336
rect 231534 59606 233003 59666
rect 225965 59331 226031 59334
rect 228909 59331 228975 59334
rect 223481 59258 223547 59261
rect 224910 59258 224970 59331
rect 223481 59256 224970 59258
rect 223481 59200 223486 59256
rect 223542 59200 224970 59256
rect 223481 59198 224970 59200
rect 230197 59258 230263 59261
rect 231534 59258 231594 59606
rect 231761 59530 231827 59533
rect 233774 59530 233834 60044
rect 234606 59802 234666 60044
rect 235438 59805 235498 60044
rect 235257 59802 235323 59805
rect 234606 59800 235323 59802
rect 234606 59744 235262 59800
rect 235318 59744 235323 59800
rect 234606 59742 235323 59744
rect 235438 59800 235507 59805
rect 235438 59744 235446 59800
rect 235502 59744 235507 59800
rect 235438 59742 235507 59744
rect 236269 59802 236329 60044
rect 236913 59802 236979 59805
rect 236269 59800 236979 59802
rect 236269 59744 236918 59800
rect 236974 59744 236979 59800
rect 236269 59742 236979 59744
rect 235257 59739 235323 59742
rect 235441 59739 235507 59742
rect 236913 59739 236979 59742
rect 234245 59666 234311 59669
rect 237101 59666 237161 60044
rect 234245 59664 237161 59666
rect 234245 59608 234250 59664
rect 234306 59608 237161 59664
rect 234245 59606 237161 59608
rect 234245 59603 234311 59606
rect 231761 59528 233834 59530
rect 231761 59472 231766 59528
rect 231822 59472 233834 59528
rect 231761 59470 233834 59472
rect 235901 59530 235967 59533
rect 237932 59530 237992 60044
rect 238764 59938 238824 60044
rect 235901 59528 237992 59530
rect 235901 59472 235906 59528
rect 235962 59472 237992 59528
rect 235901 59470 237992 59472
rect 238158 59878 238824 59938
rect 239596 59938 239656 60044
rect 240427 59938 240487 60044
rect 239596 59878 239874 59938
rect 231761 59467 231827 59470
rect 235901 59467 235967 59470
rect 232957 59394 233023 59397
rect 235441 59394 235507 59397
rect 232957 59392 235507 59394
rect 232957 59336 232962 59392
rect 233018 59336 235446 59392
rect 235502 59336 235507 59392
rect 232957 59334 235507 59336
rect 232957 59331 233023 59334
rect 235441 59331 235507 59334
rect 237281 59394 237347 59397
rect 238158 59394 238218 59878
rect 239814 59802 239874 59878
rect 240182 59878 240487 59938
rect 239949 59802 240015 59805
rect 239814 59800 240015 59802
rect 239814 59744 239954 59800
rect 240010 59744 240015 59800
rect 239814 59742 240015 59744
rect 239949 59739 240015 59742
rect 238385 59666 238451 59669
rect 240182 59666 240242 59878
rect 240593 59802 240659 59805
rect 241259 59802 241319 60044
rect 240593 59800 241319 59802
rect 240593 59744 240598 59800
rect 240654 59744 241319 59800
rect 240593 59742 241319 59744
rect 240593 59739 240659 59742
rect 242090 59666 242150 60044
rect 238385 59664 240242 59666
rect 238385 59608 238390 59664
rect 238446 59608 240242 59664
rect 238385 59606 240242 59608
rect 240550 59606 242150 59666
rect 238385 59603 238451 59606
rect 237281 59392 238218 59394
rect 237281 59336 237286 59392
rect 237342 59336 238218 59392
rect 237281 59334 238218 59336
rect 240041 59394 240107 59397
rect 240550 59394 240610 59606
rect 241329 59530 241395 59533
rect 242922 59530 242982 60044
rect 241329 59528 242982 59530
rect 241329 59472 241334 59528
rect 241390 59472 242982 59528
rect 241329 59470 242982 59472
rect 241329 59467 241395 59470
rect 240041 59392 240610 59394
rect 240041 59336 240046 59392
rect 240102 59336 240610 59392
rect 240041 59334 240610 59336
rect 241145 59394 241211 59397
rect 243754 59394 243814 60044
rect 244585 59938 244645 60044
rect 244230 59878 244645 59938
rect 244230 59802 244290 59878
rect 241145 59392 243814 59394
rect 241145 59336 241150 59392
rect 241206 59336 243814 59392
rect 241145 59334 243814 59336
rect 244046 59742 244290 59802
rect 244733 59802 244799 59805
rect 245417 59802 245477 60044
rect 244733 59800 245477 59802
rect 244733 59744 244738 59800
rect 244794 59744 245477 59800
rect 244733 59742 245477 59744
rect 237281 59331 237347 59334
rect 240041 59331 240107 59334
rect 241145 59331 241211 59334
rect 230197 59256 231594 59258
rect 230197 59200 230202 59256
rect 230258 59200 231594 59256
rect 230197 59198 231594 59200
rect 242525 59258 242591 59261
rect 244046 59258 244106 59742
rect 244733 59739 244799 59742
rect 244181 59666 244247 59669
rect 246248 59666 246308 60044
rect 244181 59664 246308 59666
rect 244181 59608 244186 59664
rect 244242 59608 246308 59664
rect 244181 59606 246308 59608
rect 244181 59603 244247 59606
rect 245469 59530 245535 59533
rect 247080 59530 247140 60044
rect 245469 59528 247140 59530
rect 245469 59472 245474 59528
rect 245530 59472 247140 59528
rect 245469 59470 247140 59472
rect 245469 59467 245535 59470
rect 245285 59394 245351 59397
rect 247912 59394 247972 60044
rect 248743 59394 248803 60044
rect 248873 59530 248939 59533
rect 249575 59530 249635 60044
rect 249701 59802 249767 59805
rect 250406 59802 250466 60044
rect 251238 59938 251298 60044
rect 252070 59938 252130 60044
rect 250670 59878 251298 59938
rect 251406 59878 252130 59938
rect 249701 59800 250466 59802
rect 249701 59744 249706 59800
rect 249762 59744 250466 59800
rect 249701 59742 250466 59744
rect 250529 59802 250595 59805
rect 250670 59802 250730 59878
rect 250529 59800 250730 59802
rect 250529 59744 250534 59800
rect 250590 59744 250730 59800
rect 250529 59742 250730 59744
rect 249701 59739 249767 59742
rect 250529 59739 250595 59742
rect 249701 59666 249767 59669
rect 251406 59666 251466 59878
rect 249701 59664 251466 59666
rect 249701 59608 249706 59664
rect 249762 59608 251466 59664
rect 249701 59606 251466 59608
rect 252277 59666 252343 59669
rect 252901 59666 252961 60044
rect 253733 59938 253793 60044
rect 252277 59664 252961 59666
rect 252277 59608 252282 59664
rect 252338 59608 252961 59664
rect 252277 59606 252961 59608
rect 253062 59878 253793 59938
rect 249701 59603 249767 59606
rect 252277 59603 252343 59606
rect 248873 59528 249635 59530
rect 248873 59472 248878 59528
rect 248934 59472 249635 59528
rect 248873 59470 249635 59472
rect 251081 59530 251147 59533
rect 251081 59528 252570 59530
rect 251081 59472 251086 59528
rect 251142 59472 252570 59528
rect 251081 59470 252570 59472
rect 248873 59467 248939 59470
rect 251081 59467 251147 59470
rect 245285 59392 247972 59394
rect 245285 59336 245290 59392
rect 245346 59336 247972 59392
rect 245285 59334 247972 59336
rect 248094 59334 248803 59394
rect 249609 59394 249675 59397
rect 250529 59394 250595 59397
rect 249609 59392 250595 59394
rect 249609 59336 249614 59392
rect 249670 59336 250534 59392
rect 250590 59336 250595 59392
rect 249609 59334 250595 59336
rect 245285 59331 245351 59334
rect 242525 59256 244106 59258
rect 242525 59200 242530 59256
rect 242586 59200 244106 59256
rect 242525 59198 244106 59200
rect 246849 59258 246915 59261
rect 248094 59258 248154 59334
rect 249609 59331 249675 59334
rect 250529 59331 250595 59334
rect 250989 59394 251055 59397
rect 252277 59394 252343 59397
rect 250989 59392 252343 59394
rect 250989 59336 250994 59392
rect 251050 59336 252282 59392
rect 252338 59336 252343 59392
rect 250989 59334 252343 59336
rect 252510 59394 252570 59470
rect 253062 59394 253122 59878
rect 253197 59802 253263 59805
rect 254564 59802 254624 60044
rect 253197 59800 254624 59802
rect 253197 59744 253202 59800
rect 253258 59744 254624 59800
rect 253197 59742 254624 59744
rect 253197 59739 253263 59742
rect 253381 59666 253447 59669
rect 255396 59666 255456 60044
rect 253381 59664 255456 59666
rect 253381 59608 253386 59664
rect 253442 59608 255456 59664
rect 253381 59606 255456 59608
rect 255589 59666 255655 59669
rect 256228 59666 256288 60044
rect 255589 59664 256288 59666
rect 255589 59608 255594 59664
rect 255650 59608 256288 59664
rect 255589 59606 256288 59608
rect 253381 59603 253447 59606
rect 255589 59603 255655 59606
rect 254761 59530 254827 59533
rect 257059 59530 257119 60044
rect 257429 59802 257495 59805
rect 257891 59802 257951 60044
rect 257429 59800 257951 59802
rect 257429 59744 257434 59800
rect 257490 59744 257951 59800
rect 257429 59742 257951 59744
rect 257429 59739 257495 59742
rect 257245 59666 257311 59669
rect 258722 59666 258782 60044
rect 257245 59664 258782 59666
rect 257245 59608 257250 59664
rect 257306 59608 258782 59664
rect 257245 59606 258782 59608
rect 258901 59666 258967 59669
rect 259554 59666 259614 60044
rect 258901 59664 259614 59666
rect 258901 59608 258906 59664
rect 258962 59608 259614 59664
rect 258901 59606 259614 59608
rect 257245 59603 257311 59606
rect 258901 59603 258967 59606
rect 254761 59528 257119 59530
rect 254761 59472 254766 59528
rect 254822 59472 257119 59528
rect 254761 59470 257119 59472
rect 258073 59530 258139 59533
rect 260386 59530 260446 60044
rect 260557 59666 260623 59669
rect 261217 59666 261277 60044
rect 260557 59664 261277 59666
rect 260557 59608 260562 59664
rect 260618 59608 261277 59664
rect 260557 59606 261277 59608
rect 260557 59603 260623 59606
rect 258073 59528 260446 59530
rect 258073 59472 258078 59528
rect 258134 59472 260446 59528
rect 258073 59470 260446 59472
rect 260557 59530 260623 59533
rect 262049 59530 262109 60044
rect 260557 59528 262109 59530
rect 260557 59472 260562 59528
rect 260618 59472 262109 59528
rect 260557 59470 262109 59472
rect 254761 59467 254827 59470
rect 258073 59467 258139 59470
rect 260557 59467 260623 59470
rect 252510 59334 253122 59394
rect 253197 59394 253263 59397
rect 255589 59394 255655 59397
rect 257429 59394 257495 59397
rect 258901 59394 258967 59397
rect 253197 59392 255655 59394
rect 253197 59336 253202 59392
rect 253258 59336 255594 59392
rect 255650 59336 255655 59392
rect 253197 59334 255655 59336
rect 250989 59331 251055 59334
rect 252277 59331 252343 59334
rect 253197 59331 253263 59334
rect 255589 59331 255655 59334
rect 255822 59392 257495 59394
rect 255822 59336 257434 59392
rect 257490 59336 257495 59392
rect 255822 59334 257495 59336
rect 246849 59256 248154 59258
rect 246849 59200 246854 59256
rect 246910 59200 248154 59256
rect 246849 59198 248154 59200
rect 254577 59258 254643 59261
rect 255822 59258 255882 59334
rect 257429 59331 257495 59334
rect 258030 59392 258967 59394
rect 258030 59336 258906 59392
rect 258962 59336 258967 59392
rect 258030 59334 258967 59336
rect 254577 59256 255882 59258
rect 254577 59200 254582 59256
rect 254638 59200 255882 59256
rect 254577 59198 255882 59200
rect 257521 59258 257587 59261
rect 258030 59258 258090 59334
rect 258901 59331 258967 59334
rect 260097 59394 260163 59397
rect 262880 59394 262940 60044
rect 263712 59394 263772 60044
rect 264544 59394 264604 60044
rect 260097 59392 262940 59394
rect 260097 59336 260102 59392
rect 260158 59336 262940 59392
rect 260097 59334 262940 59336
rect 263182 59334 263772 59394
rect 263918 59334 264604 59394
rect 265375 59394 265435 60044
rect 266207 59530 266267 60044
rect 267038 59802 267098 60044
rect 267733 59802 267799 59805
rect 267038 59800 267799 59802
rect 267038 59744 267738 59800
rect 267794 59744 267799 59800
rect 267038 59742 267799 59744
rect 267733 59739 267799 59742
rect 267733 59530 267799 59533
rect 266207 59528 267799 59530
rect 266207 59472 267738 59528
rect 267794 59472 267799 59528
rect 266207 59470 267799 59472
rect 267733 59467 267799 59470
rect 267870 59394 267930 60044
rect 268193 59530 268259 59533
rect 268702 59530 268762 60044
rect 268193 59528 268762 59530
rect 268193 59472 268198 59528
rect 268254 59472 268762 59528
rect 268193 59470 268762 59472
rect 268193 59467 268259 59470
rect 269533 59394 269593 60044
rect 270365 59530 270425 60044
rect 271196 59666 271256 60044
rect 272028 59802 272088 60044
rect 272701 59802 272767 59805
rect 272028 59800 272767 59802
rect 272028 59744 272706 59800
rect 272762 59744 272767 59800
rect 272028 59742 272767 59744
rect 272701 59739 272767 59742
rect 271196 59606 272626 59666
rect 271873 59530 271939 59533
rect 270365 59528 271939 59530
rect 270365 59472 271878 59528
rect 271934 59472 271939 59528
rect 270365 59470 271939 59472
rect 271873 59467 271939 59470
rect 271965 59394 272031 59397
rect 265375 59334 267750 59394
rect 267870 59334 269314 59394
rect 269533 59392 272031 59394
rect 269533 59336 271970 59392
rect 272026 59336 272031 59392
rect 269533 59334 272031 59336
rect 260097 59331 260163 59334
rect 257521 59256 258090 59258
rect 257521 59200 257526 59256
rect 257582 59200 258090 59256
rect 257521 59198 258090 59200
rect 262121 59258 262187 59261
rect 263182 59258 263242 59334
rect 262121 59256 263242 59258
rect 262121 59200 262126 59256
rect 262182 59200 263242 59256
rect 262121 59198 263242 59200
rect 223481 59195 223547 59198
rect 230197 59195 230263 59198
rect 242525 59195 242591 59198
rect 246849 59195 246915 59198
rect 254577 59195 254643 59198
rect 257521 59195 257587 59198
rect 262121 59195 262187 59198
rect 217685 59120 218346 59122
rect 217685 59064 217690 59120
rect 217746 59064 218346 59120
rect 217685 59062 218346 59064
rect 262029 59122 262095 59125
rect 263918 59122 263978 59334
rect 267690 59258 267750 59334
rect 268009 59258 268075 59261
rect 267690 59256 268075 59258
rect 267690 59200 268014 59256
rect 268070 59200 268075 59256
rect 267690 59198 268075 59200
rect 269254 59258 269314 59334
rect 271965 59331 272031 59334
rect 270677 59258 270743 59261
rect 269254 59256 270743 59258
rect 269254 59200 270682 59256
rect 270738 59200 270743 59256
rect 269254 59198 270743 59200
rect 272566 59258 272626 59606
rect 272860 59394 272920 60044
rect 273691 59394 273751 60044
rect 274523 59530 274583 60044
rect 275354 59666 275414 60044
rect 276186 59802 276246 60044
rect 276841 59802 276907 59805
rect 276186 59800 276907 59802
rect 276186 59744 276846 59800
rect 276902 59744 276907 59800
rect 276186 59742 276907 59744
rect 276841 59739 276907 59742
rect 275354 59606 276858 59666
rect 276289 59530 276355 59533
rect 274523 59528 276355 59530
rect 274523 59472 276294 59528
rect 276350 59472 276355 59528
rect 274523 59470 276355 59472
rect 276289 59467 276355 59470
rect 272860 59334 273546 59394
rect 273691 59334 275202 59394
rect 273345 59258 273411 59261
rect 272566 59256 273411 59258
rect 272566 59200 273350 59256
rect 273406 59200 273411 59256
rect 272566 59198 273411 59200
rect 273486 59258 273546 59334
rect 274909 59258 274975 59261
rect 273486 59256 274975 59258
rect 273486 59200 274914 59256
rect 274970 59200 274975 59256
rect 273486 59198 274975 59200
rect 275142 59258 275202 59334
rect 276105 59258 276171 59261
rect 275142 59256 276171 59258
rect 275142 59200 276110 59256
rect 276166 59200 276171 59256
rect 275142 59198 276171 59200
rect 276798 59258 276858 59606
rect 277018 59394 277078 60044
rect 277393 59394 277459 59397
rect 277018 59392 277459 59394
rect 277018 59336 277398 59392
rect 277454 59336 277459 59392
rect 277018 59334 277459 59336
rect 277849 59394 277909 60044
rect 278681 59530 278741 60044
rect 279512 59666 279572 60044
rect 280061 59802 280127 59805
rect 280344 59802 280404 60044
rect 280061 59800 280404 59802
rect 280061 59744 280066 59800
rect 280122 59744 280404 59800
rect 280061 59742 280404 59744
rect 280061 59739 280127 59742
rect 279512 59606 281090 59666
rect 280153 59530 280219 59533
rect 278681 59528 280219 59530
rect 278681 59472 280158 59528
rect 280214 59472 280219 59528
rect 278681 59470 280219 59472
rect 280153 59467 280219 59470
rect 280337 59394 280403 59397
rect 277849 59392 280403 59394
rect 277849 59336 280342 59392
rect 280398 59336 280403 59392
rect 277849 59334 280403 59336
rect 277393 59331 277459 59334
rect 280337 59331 280403 59334
rect 277485 59258 277551 59261
rect 276798 59256 277551 59258
rect 276798 59200 277490 59256
rect 277546 59200 277551 59256
rect 276798 59198 277551 59200
rect 281030 59258 281090 59606
rect 281176 59394 281236 60044
rect 282007 59530 282067 60044
rect 282637 59530 282703 59533
rect 282007 59528 282703 59530
rect 282007 59472 282642 59528
rect 282698 59472 282703 59528
rect 282007 59470 282703 59472
rect 282839 59530 282899 60044
rect 283670 59530 283730 60044
rect 284502 59666 284562 60044
rect 285121 59666 285187 59669
rect 284502 59664 285187 59666
rect 284502 59608 285126 59664
rect 285182 59608 285187 59664
rect 284502 59606 285187 59608
rect 285334 59666 285394 60044
rect 286165 59802 286225 60044
rect 286997 59938 287057 60044
rect 287828 59938 287888 60044
rect 286918 59878 287057 59938
rect 287286 59878 287888 59938
rect 286777 59802 286843 59805
rect 286165 59800 286843 59802
rect 286165 59744 286782 59800
rect 286838 59744 286843 59800
rect 286165 59742 286843 59744
rect 286777 59739 286843 59742
rect 286918 59666 286978 59878
rect 287053 59802 287119 59805
rect 287286 59802 287346 59878
rect 287053 59800 287346 59802
rect 287053 59744 287058 59800
rect 287114 59744 287346 59800
rect 287053 59742 287346 59744
rect 287053 59739 287119 59742
rect 288660 59666 288720 60044
rect 285334 59606 286794 59666
rect 286918 59606 287057 59666
rect 288660 59606 289370 59666
rect 285121 59603 285187 59606
rect 285673 59530 285739 59533
rect 282839 59470 283482 59530
rect 283670 59528 285739 59530
rect 283670 59472 285678 59528
rect 285734 59472 285739 59528
rect 283670 59470 285739 59472
rect 282637 59467 282703 59470
rect 282913 59394 282979 59397
rect 281176 59392 282979 59394
rect 281176 59336 282918 59392
rect 282974 59336 282979 59392
rect 281176 59334 282979 59336
rect 283422 59394 283482 59470
rect 285673 59467 285739 59470
rect 284385 59394 284451 59397
rect 283422 59392 284451 59394
rect 283422 59336 284390 59392
rect 284446 59336 284451 59392
rect 283422 59334 284451 59336
rect 282913 59331 282979 59334
rect 284385 59331 284451 59334
rect 285121 59394 285187 59397
rect 286734 59394 286794 59606
rect 286997 59530 287057 59606
rect 288617 59530 288683 59533
rect 286997 59528 288683 59530
rect 286997 59472 288622 59528
rect 288678 59472 288683 59528
rect 286997 59470 288683 59472
rect 288617 59467 288683 59470
rect 287421 59394 287487 59397
rect 285121 59392 286610 59394
rect 285121 59336 285126 59392
rect 285182 59336 286610 59392
rect 285121 59334 286610 59336
rect 286734 59392 287487 59394
rect 286734 59336 287426 59392
rect 287482 59336 287487 59392
rect 286734 59334 287487 59336
rect 289310 59394 289370 59606
rect 289492 59530 289552 60044
rect 290323 59666 290383 60044
rect 291155 59802 291215 60044
rect 291837 59802 291903 59805
rect 291155 59800 291903 59802
rect 291155 59744 291842 59800
rect 291898 59744 291903 59800
rect 291155 59742 291903 59744
rect 291837 59739 291903 59742
rect 290323 59606 291762 59666
rect 291561 59530 291627 59533
rect 289492 59528 291627 59530
rect 289492 59472 291566 59528
rect 291622 59472 291627 59528
rect 289492 59470 291627 59472
rect 291561 59467 291627 59470
rect 291702 59394 291762 59606
rect 291986 59530 292046 60044
rect 292818 59666 292878 60044
rect 293493 59666 293559 59669
rect 292818 59664 293559 59666
rect 292818 59608 293498 59664
rect 293554 59608 293559 59664
rect 292818 59606 293559 59608
rect 293650 59666 293710 60044
rect 293650 59606 294338 59666
rect 293493 59603 293559 59606
rect 294045 59530 294111 59533
rect 291986 59528 294111 59530
rect 291986 59472 294050 59528
rect 294106 59472 294111 59528
rect 291986 59470 294111 59472
rect 294045 59467 294111 59470
rect 292665 59394 292731 59397
rect 289310 59334 290106 59394
rect 291702 59392 292731 59394
rect 291702 59336 292670 59392
rect 292726 59336 292731 59392
rect 291702 59334 292731 59336
rect 294278 59394 294338 59606
rect 294481 59530 294541 60044
rect 295313 59666 295373 60044
rect 295977 59666 296043 59669
rect 295313 59664 296043 59666
rect 295313 59608 295982 59664
rect 296038 59608 296043 59664
rect 295313 59606 296043 59608
rect 296144 59666 296204 60044
rect 296805 59666 296871 59669
rect 296144 59664 296871 59666
rect 296144 59608 296810 59664
rect 296866 59608 296871 59664
rect 296144 59606 296871 59608
rect 295977 59603 296043 59606
rect 296805 59603 296871 59606
rect 296713 59530 296779 59533
rect 294481 59528 296779 59530
rect 294481 59472 296718 59528
rect 296774 59472 296779 59528
rect 294481 59470 296779 59472
rect 296713 59467 296779 59470
rect 295977 59394 296043 59397
rect 296976 59394 297036 60044
rect 297808 59530 297868 60044
rect 298639 59666 298699 60044
rect 299471 59802 299531 60044
rect 300117 59802 300183 59805
rect 299471 59800 300183 59802
rect 299471 59744 300122 59800
rect 300178 59744 300183 59800
rect 299471 59742 300183 59744
rect 300302 59802 300362 60044
rect 300945 59802 301011 59805
rect 300302 59800 301011 59802
rect 300302 59744 300950 59800
rect 301006 59744 301011 59800
rect 300302 59742 301011 59744
rect 301134 59802 301194 60044
rect 301773 59802 301839 59805
rect 301134 59800 301839 59802
rect 301134 59744 301778 59800
rect 301834 59744 301839 59800
rect 301134 59742 301839 59744
rect 300117 59739 300183 59742
rect 300945 59739 301011 59742
rect 301773 59739 301839 59742
rect 301497 59666 301563 59669
rect 298639 59664 301563 59666
rect 298639 59608 301502 59664
rect 301558 59608 301563 59664
rect 298639 59606 301563 59608
rect 301497 59603 301563 59606
rect 300117 59530 300183 59533
rect 297808 59528 300183 59530
rect 297808 59472 300122 59528
rect 300178 59472 300183 59528
rect 297808 59470 300183 59472
rect 301966 59530 302026 60044
rect 302797 59802 302857 60044
rect 303429 59802 303495 59805
rect 302797 59800 303495 59802
rect 302797 59744 303434 59800
rect 303490 59744 303495 59800
rect 302797 59742 303495 59744
rect 303429 59739 303495 59742
rect 303629 59666 303689 60044
rect 304460 59802 304520 60044
rect 305292 59938 305352 60044
rect 305292 59878 305746 59938
rect 305361 59802 305427 59805
rect 304460 59800 305427 59802
rect 304460 59744 305366 59800
rect 305422 59744 305427 59800
rect 304460 59742 305427 59744
rect 305686 59802 305746 59878
rect 305821 59802 305887 59805
rect 305686 59800 305887 59802
rect 305686 59744 305826 59800
rect 305882 59744 305887 59800
rect 305686 59742 305887 59744
rect 305361 59739 305427 59742
rect 305821 59739 305887 59742
rect 305913 59666 305979 59669
rect 303629 59664 305979 59666
rect 303629 59608 305918 59664
rect 305974 59608 305979 59664
rect 303629 59606 305979 59608
rect 305913 59603 305979 59606
rect 304257 59530 304323 59533
rect 301966 59528 304323 59530
rect 301966 59472 304262 59528
rect 304318 59472 304323 59528
rect 301966 59470 304323 59472
rect 306124 59530 306184 60044
rect 306741 59530 306807 59533
rect 306124 59528 306807 59530
rect 306124 59472 306746 59528
rect 306802 59472 306807 59528
rect 306124 59470 306807 59472
rect 306955 59530 307015 60044
rect 307787 59666 307847 60044
rect 308618 59802 308678 60044
rect 309317 59802 309383 59805
rect 308618 59800 309383 59802
rect 308618 59744 309322 59800
rect 309378 59744 309383 59800
rect 308618 59742 309383 59744
rect 309450 59802 309510 60044
rect 310282 59938 310342 60044
rect 310282 59878 310898 59938
rect 310697 59802 310763 59805
rect 309450 59800 310763 59802
rect 309450 59744 310702 59800
rect 310758 59744 310763 59800
rect 309450 59742 310763 59744
rect 309317 59739 309383 59742
rect 310697 59739 310763 59742
rect 307787 59606 310162 59666
rect 309869 59530 309935 59533
rect 306955 59528 309935 59530
rect 306955 59472 309874 59528
rect 309930 59472 309935 59528
rect 306955 59470 309935 59472
rect 310102 59530 310162 59606
rect 310697 59530 310763 59533
rect 310102 59528 310763 59530
rect 310102 59472 310702 59528
rect 310758 59472 310763 59528
rect 310102 59470 310763 59472
rect 310838 59530 310898 59878
rect 311113 59802 311173 60044
rect 311945 59938 312005 60044
rect 311942 59878 312005 59938
rect 311801 59802 311867 59805
rect 311113 59800 311867 59802
rect 311113 59744 311806 59800
rect 311862 59744 311867 59800
rect 311113 59742 311867 59744
rect 311801 59739 311867 59742
rect 311942 59666 312002 59878
rect 312776 59802 312836 60044
rect 313457 59802 313523 59805
rect 312776 59800 313523 59802
rect 312776 59744 313462 59800
rect 313518 59744 313523 59800
rect 312776 59742 313523 59744
rect 313608 59802 313668 60044
rect 314285 59802 314351 59805
rect 313608 59800 314351 59802
rect 313608 59744 314290 59800
rect 314346 59744 314351 59800
rect 313608 59742 314351 59744
rect 313457 59739 313523 59742
rect 314285 59739 314351 59742
rect 314285 59666 314351 59669
rect 311942 59664 314351 59666
rect 311942 59608 314290 59664
rect 314346 59608 314351 59664
rect 311942 59606 314351 59608
rect 314285 59603 314351 59606
rect 312721 59530 312787 59533
rect 310838 59528 312787 59530
rect 310838 59472 312726 59528
rect 312782 59472 312787 59528
rect 310838 59470 312787 59472
rect 314440 59530 314500 60044
rect 315271 59938 315331 60044
rect 315254 59878 315331 59938
rect 316103 59938 316163 60044
rect 316103 59878 316786 59938
rect 315254 59666 315314 59878
rect 315389 59802 315455 59805
rect 316585 59802 316651 59805
rect 315389 59800 316651 59802
rect 315389 59744 315394 59800
rect 315450 59744 316590 59800
rect 316646 59744 316651 59800
rect 315389 59742 316651 59744
rect 315389 59739 315455 59742
rect 316585 59739 316651 59742
rect 316585 59666 316651 59669
rect 315254 59664 316651 59666
rect 315254 59608 316590 59664
rect 316646 59608 316651 59664
rect 315254 59606 316651 59608
rect 316585 59603 316651 59606
rect 316585 59530 316651 59533
rect 314440 59528 316651 59530
rect 314440 59472 316590 59528
rect 316646 59472 316651 59528
rect 314440 59470 316651 59472
rect 300117 59467 300183 59470
rect 304257 59467 304323 59470
rect 306741 59467 306807 59470
rect 309869 59467 309935 59470
rect 310697 59467 310763 59470
rect 312721 59467 312787 59470
rect 316585 59467 316651 59470
rect 300945 59394 301011 59397
rect 302877 59394 302943 59397
rect 294278 59334 295074 59394
rect 285121 59331 285187 59334
rect 281533 59258 281599 59261
rect 281030 59256 281599 59258
rect 281030 59200 281538 59256
rect 281594 59200 281599 59256
rect 281030 59198 281599 59200
rect 286550 59258 286610 59334
rect 287421 59331 287487 59334
rect 287237 59258 287303 59261
rect 286550 59256 287303 59258
rect 286550 59200 287242 59256
rect 287298 59200 287303 59256
rect 286550 59198 287303 59200
rect 290046 59258 290106 59334
rect 292665 59331 292731 59334
rect 291377 59258 291443 59261
rect 290046 59256 291443 59258
rect 290046 59200 291382 59256
rect 291438 59200 291443 59256
rect 290046 59198 291443 59200
rect 295014 59258 295074 59334
rect 295977 59392 296914 59394
rect 295977 59336 295982 59392
rect 296038 59336 296914 59392
rect 295977 59334 296914 59336
rect 296976 59334 300226 59394
rect 295977 59331 296043 59334
rect 295701 59258 295767 59261
rect 295014 59256 295767 59258
rect 295014 59200 295706 59256
rect 295762 59200 295767 59256
rect 295014 59198 295767 59200
rect 296854 59258 296914 59334
rect 298921 59258 298987 59261
rect 296854 59256 298987 59258
rect 296854 59200 298926 59256
rect 298982 59200 298987 59256
rect 296854 59198 298987 59200
rect 300166 59258 300226 59334
rect 300945 59392 302943 59394
rect 300945 59336 300950 59392
rect 301006 59336 302882 59392
rect 302938 59336 302943 59392
rect 300945 59334 302943 59336
rect 300945 59331 301011 59334
rect 302877 59331 302943 59334
rect 305361 59394 305427 59397
rect 307201 59394 307267 59397
rect 305361 59392 307267 59394
rect 305361 59336 305366 59392
rect 305422 59336 307206 59392
rect 307262 59336 307267 59392
rect 305361 59334 307267 59336
rect 305361 59331 305427 59334
rect 307201 59331 307267 59334
rect 309317 59394 309383 59397
rect 311341 59394 311407 59397
rect 309317 59392 311407 59394
rect 309317 59336 309322 59392
rect 309378 59336 311346 59392
rect 311402 59336 311407 59392
rect 309317 59334 311407 59336
rect 309317 59331 309383 59334
rect 311341 59331 311407 59334
rect 311801 59394 311867 59397
rect 313457 59394 313523 59397
rect 315297 59394 315363 59397
rect 311801 59392 313106 59394
rect 311801 59336 311806 59392
rect 311862 59336 313106 59392
rect 311801 59334 313106 59336
rect 311801 59331 311867 59334
rect 300301 59258 300367 59261
rect 300166 59256 300367 59258
rect 300166 59200 300306 59256
rect 300362 59200 300367 59256
rect 300166 59198 300367 59200
rect 313046 59258 313106 59334
rect 313457 59392 315363 59394
rect 313457 59336 313462 59392
rect 313518 59336 315302 59392
rect 315358 59336 315363 59392
rect 313457 59334 315363 59336
rect 316726 59394 316786 59878
rect 316934 59530 316994 60044
rect 317766 59802 317826 60044
rect 318598 59938 318658 60044
rect 318598 59878 319178 59938
rect 318425 59802 318491 59805
rect 317766 59800 318491 59802
rect 317766 59744 318430 59800
rect 318486 59744 318491 59800
rect 317766 59742 318491 59744
rect 319118 59802 319178 59878
rect 319253 59802 319319 59805
rect 319118 59800 319319 59802
rect 319118 59744 319258 59800
rect 319314 59744 319319 59800
rect 319118 59742 319319 59744
rect 318425 59739 318491 59742
rect 319253 59739 319319 59742
rect 319429 59666 319489 60044
rect 320261 59802 320321 60044
rect 320817 59802 320883 59805
rect 320261 59800 320883 59802
rect 320261 59744 320822 59800
rect 320878 59744 320883 59800
rect 320261 59742 320883 59744
rect 320817 59739 320883 59742
rect 319429 59606 320834 59666
rect 319437 59530 319503 59533
rect 316934 59528 319503 59530
rect 316934 59472 319442 59528
rect 319498 59472 319503 59528
rect 316934 59470 319503 59472
rect 319437 59467 319503 59470
rect 319621 59394 319687 59397
rect 316726 59392 319687 59394
rect 316726 59336 319626 59392
rect 319682 59336 319687 59392
rect 316726 59334 319687 59336
rect 320774 59394 320834 59606
rect 321092 59530 321152 60044
rect 321737 59530 321803 59533
rect 321092 59528 321803 59530
rect 321092 59472 321742 59528
rect 321798 59472 321803 59528
rect 321092 59470 321803 59472
rect 321737 59467 321803 59470
rect 321737 59394 321803 59397
rect 320774 59392 321803 59394
rect 320774 59336 321742 59392
rect 321798 59336 321803 59392
rect 320774 59334 321803 59336
rect 321924 59394 321984 60044
rect 322756 59530 322816 60044
rect 323587 59666 323647 60044
rect 324419 59802 324479 60044
rect 325049 59802 325115 59805
rect 324419 59800 325115 59802
rect 324419 59744 325054 59800
rect 325110 59744 325115 59800
rect 324419 59742 325115 59744
rect 325250 59802 325310 60044
rect 325877 59802 325943 59805
rect 325250 59800 325943 59802
rect 325250 59744 325882 59800
rect 325938 59744 325943 59800
rect 325250 59742 325943 59744
rect 326082 59802 326142 60044
rect 326705 59802 326771 59805
rect 326082 59800 326771 59802
rect 326082 59744 326710 59800
rect 326766 59744 326771 59800
rect 326082 59742 326771 59744
rect 325049 59739 325115 59742
rect 325877 59739 325943 59742
rect 326705 59739 326771 59742
rect 326337 59666 326403 59669
rect 323587 59664 326403 59666
rect 323587 59608 326342 59664
rect 326398 59608 326403 59664
rect 323587 59606 326403 59608
rect 326337 59603 326403 59606
rect 324957 59530 325023 59533
rect 322756 59528 325023 59530
rect 322756 59472 324962 59528
rect 325018 59472 325023 59528
rect 322756 59470 325023 59472
rect 326914 59530 326974 60044
rect 327745 59666 327805 60044
rect 328361 59666 328427 59669
rect 327745 59664 328427 59666
rect 327745 59608 328366 59664
rect 328422 59608 328427 59664
rect 327745 59606 328427 59608
rect 328577 59666 328637 60044
rect 329408 59802 329468 60044
rect 330109 59802 330175 59805
rect 329408 59800 330175 59802
rect 329408 59744 330114 59800
rect 330170 59744 330175 59800
rect 329408 59742 330175 59744
rect 330240 59802 330300 60044
rect 330937 59802 331003 59805
rect 330240 59800 331003 59802
rect 330240 59744 330942 59800
rect 330998 59744 331003 59800
rect 330240 59742 331003 59744
rect 330109 59739 330175 59742
rect 330937 59739 331003 59742
rect 330845 59666 330911 59669
rect 328577 59664 330911 59666
rect 328577 59608 330850 59664
rect 330906 59608 330911 59664
rect 328577 59606 330911 59608
rect 328361 59603 328427 59606
rect 330845 59603 330911 59606
rect 329281 59530 329347 59533
rect 330477 59530 330543 59533
rect 326914 59528 329347 59530
rect 326914 59472 329286 59528
rect 329342 59472 329347 59528
rect 326914 59470 329347 59472
rect 324957 59467 325023 59470
rect 329281 59467 329347 59470
rect 329974 59528 330543 59530
rect 329974 59472 330482 59528
rect 330538 59472 330543 59528
rect 329974 59470 330543 59472
rect 331072 59530 331132 60044
rect 331765 59530 331831 59533
rect 331072 59528 331831 59530
rect 331072 59472 331770 59528
rect 331826 59472 331831 59528
rect 331072 59470 331831 59472
rect 325049 59394 325115 59397
rect 321924 59392 325115 59394
rect 321924 59336 325054 59392
rect 325110 59336 325115 59392
rect 321924 59334 325115 59336
rect 313457 59331 313523 59334
rect 315297 59331 315363 59334
rect 319621 59331 319687 59334
rect 321737 59331 321803 59334
rect 325049 59331 325115 59334
rect 325877 59394 325943 59397
rect 327901 59394 327967 59397
rect 325877 59392 327967 59394
rect 325877 59336 325882 59392
rect 325938 59336 327906 59392
rect 327962 59336 327967 59392
rect 325877 59334 327967 59336
rect 325877 59331 325943 59334
rect 327901 59331 327967 59334
rect 328361 59394 328427 59397
rect 329974 59394 330034 59470
rect 330477 59467 330543 59470
rect 331765 59467 331831 59470
rect 328361 59392 330034 59394
rect 328361 59336 328366 59392
rect 328422 59336 330034 59392
rect 328361 59334 330034 59336
rect 330109 59394 330175 59397
rect 331765 59394 331831 59397
rect 330109 59392 331831 59394
rect 330109 59336 330114 59392
rect 330170 59336 331770 59392
rect 331826 59336 331831 59392
rect 330109 59334 331831 59336
rect 331903 59394 331963 60044
rect 332735 59530 332795 60044
rect 333421 59530 333487 59533
rect 332735 59528 333487 59530
rect 332735 59472 333426 59528
rect 333482 59472 333487 59528
rect 332735 59470 333487 59472
rect 333566 59530 333626 60044
rect 334398 59666 334458 60044
rect 335077 59666 335143 59669
rect 334398 59664 335143 59666
rect 334398 59608 335082 59664
rect 335138 59608 335143 59664
rect 334398 59606 335143 59608
rect 335230 59666 335290 60044
rect 336061 59802 336121 60044
rect 336893 59938 336953 60044
rect 336893 59878 337578 59938
rect 337518 59805 337578 59878
rect 337377 59802 337443 59805
rect 336061 59800 337443 59802
rect 336061 59744 337382 59800
rect 337438 59744 337443 59800
rect 336061 59742 337443 59744
rect 337518 59800 337627 59805
rect 337518 59744 337566 59800
rect 337622 59744 337627 59800
rect 337518 59742 337627 59744
rect 337377 59739 337443 59742
rect 337561 59739 337627 59742
rect 337469 59666 337535 59669
rect 335230 59664 337535 59666
rect 335230 59608 337474 59664
rect 337530 59608 337535 59664
rect 335230 59606 337535 59608
rect 335077 59603 335143 59606
rect 337469 59603 337535 59606
rect 335997 59530 336063 59533
rect 333566 59528 336063 59530
rect 333566 59472 336002 59528
rect 336058 59472 336063 59528
rect 333566 59470 336063 59472
rect 337724 59530 337784 60044
rect 338556 59666 338616 60044
rect 339217 59666 339283 59669
rect 338556 59664 339283 59666
rect 338556 59608 339222 59664
rect 339278 59608 339283 59664
rect 338556 59606 339283 59608
rect 339388 59666 339448 60044
rect 340219 59802 340279 60044
rect 341051 59938 341111 60044
rect 341882 59938 341942 60044
rect 341051 59878 341810 59938
rect 341882 59878 342546 59938
rect 341609 59802 341675 59805
rect 340219 59800 341675 59802
rect 340219 59744 341614 59800
rect 341670 59744 341675 59800
rect 340219 59742 341675 59744
rect 341609 59739 341675 59742
rect 341517 59666 341583 59669
rect 339388 59664 341583 59666
rect 339388 59608 341522 59664
rect 341578 59608 341583 59664
rect 339388 59606 341583 59608
rect 341750 59666 341810 59878
rect 342345 59666 342411 59669
rect 341750 59664 342411 59666
rect 341750 59608 342350 59664
rect 342406 59608 342411 59664
rect 341750 59606 342411 59608
rect 339217 59603 339283 59606
rect 341517 59603 341583 59606
rect 342345 59603 342411 59606
rect 340137 59530 340203 59533
rect 337724 59528 340203 59530
rect 337724 59472 340142 59528
rect 340198 59472 340203 59528
rect 337724 59470 340203 59472
rect 333421 59467 333487 59470
rect 335997 59467 336063 59470
rect 340137 59467 340203 59470
rect 341609 59530 341675 59533
rect 342486 59530 342546 59878
rect 342714 59666 342774 60044
rect 343357 59666 343423 59669
rect 342714 59664 343423 59666
rect 342714 59608 343362 59664
rect 343418 59608 343423 59664
rect 342714 59606 343423 59608
rect 343546 59666 343606 60044
rect 344377 59802 344437 60044
rect 345013 59802 345079 59805
rect 344377 59800 345079 59802
rect 344377 59744 345018 59800
rect 345074 59744 345079 59800
rect 344377 59742 345079 59744
rect 345013 59739 345079 59742
rect 345013 59666 345079 59669
rect 343546 59664 345079 59666
rect 343546 59608 345018 59664
rect 345074 59608 345079 59664
rect 343546 59606 345079 59608
rect 343357 59603 343423 59606
rect 345013 59603 345079 59606
rect 344277 59530 344343 59533
rect 341609 59528 342362 59530
rect 341609 59472 341614 59528
rect 341670 59472 342362 59528
rect 341609 59470 342362 59472
rect 342486 59528 344343 59530
rect 342486 59472 344282 59528
rect 344338 59472 344343 59528
rect 342486 59470 344343 59472
rect 341609 59467 341675 59470
rect 334617 59394 334683 59397
rect 331903 59392 334683 59394
rect 331903 59336 334622 59392
rect 334678 59336 334683 59392
rect 331903 59334 334683 59336
rect 328361 59331 328427 59334
rect 330109 59331 330175 59334
rect 331765 59331 331831 59334
rect 334617 59331 334683 59334
rect 335077 59394 335143 59397
rect 337193 59394 337259 59397
rect 335077 59392 337259 59394
rect 335077 59336 335082 59392
rect 335138 59336 337198 59392
rect 337254 59336 337259 59392
rect 335077 59334 337259 59336
rect 335077 59331 335143 59334
rect 337193 59331 337259 59334
rect 337377 59394 337443 59397
rect 338849 59394 338915 59397
rect 337377 59392 338915 59394
rect 337377 59336 337382 59392
rect 337438 59336 338854 59392
rect 338910 59336 338915 59392
rect 337377 59334 338915 59336
rect 337377 59331 337443 59334
rect 338849 59331 338915 59334
rect 339217 59394 339283 59397
rect 341609 59394 341675 59397
rect 339217 59392 341675 59394
rect 339217 59336 339222 59392
rect 339278 59336 341614 59392
rect 341670 59336 341675 59392
rect 339217 59334 341675 59336
rect 342302 59394 342362 59470
rect 344277 59467 344343 59470
rect 342897 59394 342963 59397
rect 342302 59392 342963 59394
rect 342302 59336 342902 59392
rect 342958 59336 342963 59392
rect 342302 59334 342963 59336
rect 339217 59331 339283 59334
rect 341609 59331 341675 59334
rect 342897 59331 342963 59334
rect 343357 59394 343423 59397
rect 345013 59394 345079 59397
rect 343357 59392 345079 59394
rect 343357 59336 343362 59392
rect 343418 59336 345018 59392
rect 345074 59336 345079 59392
rect 343357 59334 345079 59336
rect 345209 59394 345269 60044
rect 346040 59394 346100 60044
rect 346872 59530 346932 60044
rect 347497 59530 347563 59533
rect 346872 59528 347563 59530
rect 346872 59472 347502 59528
rect 347558 59472 347563 59528
rect 346872 59470 347563 59472
rect 347704 59530 347764 60044
rect 348535 59666 348595 60044
rect 349367 59802 349427 60044
rect 350198 59938 350258 60044
rect 351030 59938 351090 60044
rect 351862 59938 351922 60044
rect 350198 59878 350826 59938
rect 351030 59878 351792 59938
rect 351862 59878 352482 59938
rect 350625 59802 350691 59805
rect 350766 59804 350826 59878
rect 351732 59805 351792 59878
rect 349367 59800 350691 59802
rect 349367 59744 350630 59800
rect 350686 59744 350691 59800
rect 349367 59742 350691 59744
rect 350625 59739 350691 59742
rect 350758 59740 350764 59804
rect 350828 59740 350834 59804
rect 351729 59800 351795 59805
rect 351729 59744 351734 59800
rect 351790 59744 351795 59800
rect 351729 59739 351795 59744
rect 350901 59666 350967 59669
rect 348535 59664 350967 59666
rect 348535 59608 350906 59664
rect 350962 59608 350967 59664
rect 348535 59606 350967 59608
rect 350901 59603 350967 59606
rect 349797 59530 349863 59533
rect 347704 59528 349863 59530
rect 347704 59472 349802 59528
rect 349858 59472 349863 59528
rect 347704 59470 349863 59472
rect 352422 59530 352482 59878
rect 352693 59666 352753 60044
rect 353385 59666 353451 59669
rect 352693 59664 353451 59666
rect 352693 59608 353390 59664
rect 353446 59608 353451 59664
rect 352693 59606 353451 59608
rect 353525 59666 353585 60044
rect 354213 59666 354279 59669
rect 353525 59664 354279 59666
rect 353525 59608 354218 59664
rect 354274 59608 354279 59664
rect 353525 59606 354279 59608
rect 353385 59603 353451 59606
rect 354213 59603 354279 59606
rect 354029 59530 354095 59533
rect 352422 59528 354095 59530
rect 352422 59472 354034 59528
rect 354090 59472 354095 59528
rect 352422 59470 354095 59472
rect 354356 59530 354416 60044
rect 355188 59666 355248 60044
rect 356020 59802 356080 60044
rect 356697 59802 356763 59805
rect 356020 59800 356763 59802
rect 356020 59744 356702 59800
rect 356758 59744 356763 59800
rect 356020 59742 356763 59744
rect 356851 59802 356911 60044
rect 357525 59802 357591 59805
rect 356851 59800 357591 59802
rect 356851 59744 357530 59800
rect 357586 59744 357591 59800
rect 356851 59742 357591 59744
rect 356697 59739 356763 59742
rect 357525 59739 357591 59742
rect 357525 59666 357591 59669
rect 355188 59664 357591 59666
rect 355188 59608 357530 59664
rect 357586 59608 357591 59664
rect 355188 59606 357591 59608
rect 357525 59603 357591 59606
rect 356697 59530 356763 59533
rect 354356 59528 356763 59530
rect 354356 59472 356702 59528
rect 356758 59472 356763 59528
rect 354356 59470 356763 59472
rect 347497 59467 347563 59470
rect 349797 59467 349863 59470
rect 354029 59467 354095 59470
rect 356697 59467 356763 59470
rect 348601 59394 348667 59397
rect 345209 59334 345858 59394
rect 346040 59392 348667 59394
rect 346040 59336 348606 59392
rect 348662 59336 348667 59392
rect 346040 59334 348667 59336
rect 343357 59331 343423 59334
rect 345013 59331 345079 59334
rect 313917 59258 313983 59261
rect 313046 59256 313983 59258
rect 313046 59200 313922 59256
rect 313978 59200 313983 59256
rect 313046 59198 313983 59200
rect 345798 59258 345858 59334
rect 348601 59331 348667 59334
rect 354213 59394 354279 59397
rect 357683 59394 357743 60044
rect 358514 59530 358574 60044
rect 359346 59666 359406 60044
rect 360178 59802 360238 60044
rect 360837 59802 360903 59805
rect 360178 59800 360903 59802
rect 360178 59744 360842 59800
rect 360898 59744 360903 59800
rect 360178 59742 360903 59744
rect 361009 59802 361069 60044
rect 361573 59802 361639 59805
rect 361009 59800 361639 59802
rect 361009 59744 361578 59800
rect 361634 59744 361639 59800
rect 361009 59742 361639 59744
rect 360837 59739 360903 59742
rect 361573 59739 361639 59742
rect 361665 59666 361731 59669
rect 359346 59664 361731 59666
rect 359346 59608 361670 59664
rect 361726 59608 361731 59664
rect 359346 59606 361731 59608
rect 361665 59603 361731 59606
rect 360837 59530 360903 59533
rect 358514 59528 360903 59530
rect 358514 59472 360842 59528
rect 360898 59472 360903 59528
rect 358514 59470 360903 59472
rect 361841 59530 361901 60044
rect 362493 59530 362559 59533
rect 361841 59528 362559 59530
rect 361841 59472 362498 59528
rect 362554 59472 362559 59528
rect 361841 59470 362559 59472
rect 360837 59467 360903 59470
rect 362493 59467 362559 59470
rect 360101 59394 360167 59397
rect 354213 59392 356714 59394
rect 354213 59336 354218 59392
rect 354274 59336 356714 59392
rect 354213 59334 356714 59336
rect 357683 59392 360167 59394
rect 357683 59336 360106 59392
rect 360162 59336 360167 59392
rect 357683 59334 360167 59336
rect 354213 59331 354279 59334
rect 348417 59258 348483 59261
rect 345798 59256 348483 59258
rect 345798 59200 348422 59256
rect 348478 59200 348483 59256
rect 345798 59198 348483 59200
rect 356654 59258 356714 59334
rect 360101 59331 360167 59334
rect 361573 59394 361639 59397
rect 362672 59394 362732 60044
rect 363504 59530 363564 60044
rect 364336 59666 364396 60044
rect 364336 59606 364994 59666
rect 364793 59530 364859 59533
rect 363504 59528 364859 59530
rect 363504 59472 364798 59528
rect 364854 59472 364859 59528
rect 363504 59470 364859 59472
rect 364793 59467 364859 59470
rect 364333 59394 364399 59397
rect 361573 59392 362602 59394
rect 361573 59336 361578 59392
rect 361634 59336 362602 59392
rect 361573 59334 362602 59336
rect 362672 59392 364399 59394
rect 362672 59336 364338 59392
rect 364394 59336 364399 59392
rect 362672 59334 364399 59336
rect 361573 59331 361639 59334
rect 356881 59258 356947 59261
rect 356654 59256 356947 59258
rect 356654 59200 356886 59256
rect 356942 59200 356947 59256
rect 356654 59198 356947 59200
rect 362542 59258 362602 59334
rect 364333 59331 364399 59334
rect 363045 59258 363111 59261
rect 362542 59256 363111 59258
rect 362542 59200 363050 59256
rect 363106 59200 363111 59256
rect 362542 59198 363111 59200
rect 364934 59258 364994 59606
rect 365167 59394 365227 60044
rect 365999 59530 366059 60044
rect 366633 59530 366699 59533
rect 365999 59528 366699 59530
rect 365999 59472 366638 59528
rect 366694 59472 366699 59528
rect 365999 59470 366699 59472
rect 366830 59530 366890 60044
rect 367662 59666 367722 60044
rect 368494 59802 368554 60044
rect 369325 59938 369385 60044
rect 369325 59878 369594 59938
rect 369534 59805 369594 59878
rect 369117 59802 369183 59805
rect 368494 59800 369183 59802
rect 368494 59744 369122 59800
rect 369178 59744 369183 59800
rect 368494 59742 369183 59744
rect 369117 59739 369183 59742
rect 369485 59800 369594 59805
rect 369485 59744 369490 59800
rect 369546 59744 369594 59800
rect 369485 59742 369594 59744
rect 369485 59739 369551 59742
rect 369025 59666 369091 59669
rect 367662 59664 369091 59666
rect 367662 59608 369030 59664
rect 369086 59608 369091 59664
rect 367662 59606 369091 59608
rect 369025 59603 369091 59606
rect 368473 59530 368539 59533
rect 366830 59528 368539 59530
rect 366830 59472 368478 59528
rect 368534 59472 368539 59528
rect 366830 59470 368539 59472
rect 366633 59467 366699 59470
rect 368473 59467 368539 59470
rect 367277 59394 367343 59397
rect 365167 59392 367343 59394
rect 365167 59336 367282 59392
rect 367338 59336 367343 59392
rect 365167 59334 367343 59336
rect 367277 59331 367343 59334
rect 369117 59394 369183 59397
rect 370157 59394 370217 60044
rect 370988 59530 371048 60044
rect 371820 59666 371880 60044
rect 372521 59666 372587 59669
rect 371820 59664 372587 59666
rect 371820 59608 372526 59664
rect 372582 59608 372587 59664
rect 371820 59606 372587 59608
rect 372652 59666 372712 60044
rect 373483 59802 373543 60044
rect 373483 59742 374010 59802
rect 373809 59666 373875 59669
rect 372652 59664 373875 59666
rect 372652 59608 373814 59664
rect 373870 59608 373875 59664
rect 372652 59606 373875 59608
rect 372521 59603 372587 59606
rect 373809 59603 373875 59606
rect 372613 59530 372679 59533
rect 370988 59528 372679 59530
rect 370988 59472 372618 59528
rect 372674 59472 372679 59528
rect 370988 59470 372679 59472
rect 373950 59530 374010 59742
rect 374315 59666 374375 60044
rect 375146 59666 375206 60044
rect 375978 59802 376038 60044
rect 376477 59802 376543 59805
rect 375978 59800 376543 59802
rect 375978 59744 376482 59800
rect 376538 59744 376543 59800
rect 375978 59742 376543 59744
rect 376477 59739 376543 59742
rect 376661 59802 376727 59805
rect 376810 59802 376870 60044
rect 376661 59800 376870 59802
rect 376661 59744 376666 59800
rect 376722 59744 376870 59800
rect 376661 59742 376870 59744
rect 376661 59739 376727 59742
rect 376937 59666 377003 59669
rect 374315 59606 374930 59666
rect 375146 59664 377003 59666
rect 375146 59608 376942 59664
rect 376998 59608 377003 59664
rect 375146 59606 377003 59608
rect 374870 59530 374930 59606
rect 376937 59603 377003 59606
rect 376753 59530 376819 59533
rect 373950 59470 374378 59530
rect 374870 59528 376819 59530
rect 374870 59472 376758 59528
rect 376814 59472 376819 59528
rect 374870 59470 376819 59472
rect 377641 59530 377701 60044
rect 378473 59666 378533 60044
rect 379304 59802 379364 60044
rect 380136 59938 380196 60044
rect 380968 59938 381028 60044
rect 380136 59878 380818 59938
rect 380968 59878 381554 59938
rect 379973 59802 380039 59805
rect 379304 59800 380039 59802
rect 379304 59744 379978 59800
rect 380034 59744 380039 59800
rect 379304 59742 380039 59744
rect 379973 59739 380039 59742
rect 378473 59606 379898 59666
rect 379697 59530 379763 59533
rect 377641 59528 379763 59530
rect 377641 59472 379702 59528
rect 379758 59472 379763 59528
rect 377641 59470 379763 59472
rect 372613 59467 372679 59470
rect 372521 59394 372587 59397
rect 374177 59394 374243 59397
rect 369117 59392 369962 59394
rect 369117 59336 369122 59392
rect 369178 59336 369962 59392
rect 369117 59334 369962 59336
rect 370157 59334 372354 59394
rect 369117 59331 369183 59334
rect 367093 59258 367159 59261
rect 364934 59256 367159 59258
rect 364934 59200 367098 59256
rect 367154 59200 367159 59256
rect 364934 59198 367159 59200
rect 369902 59258 369962 59334
rect 371417 59258 371483 59261
rect 369902 59256 371483 59258
rect 369902 59200 371422 59256
rect 371478 59200 371483 59256
rect 369902 59198 371483 59200
rect 372294 59258 372354 59334
rect 372521 59392 374243 59394
rect 372521 59336 372526 59392
rect 372582 59336 374182 59392
rect 374238 59336 374243 59392
rect 372521 59334 374243 59336
rect 374318 59394 374378 59470
rect 376753 59467 376819 59470
rect 379697 59467 379763 59470
rect 375649 59394 375715 59397
rect 374318 59392 375715 59394
rect 374318 59336 375654 59392
rect 375710 59336 375715 59392
rect 374318 59334 375715 59336
rect 372521 59331 372587 59334
rect 374177 59331 374243 59334
rect 375649 59331 375715 59334
rect 376477 59394 376543 59397
rect 378225 59394 378291 59397
rect 376477 59392 378291 59394
rect 376477 59336 376482 59392
rect 376538 59336 378230 59392
rect 378286 59336 378291 59392
rect 376477 59334 378291 59336
rect 376477 59331 376543 59334
rect 378225 59331 378291 59334
rect 372705 59258 372771 59261
rect 372294 59256 372771 59258
rect 372294 59200 372710 59256
rect 372766 59200 372771 59256
rect 372294 59198 372771 59200
rect 379838 59258 379898 59606
rect 380758 59530 380818 59878
rect 381494 59802 381554 59878
rect 381629 59802 381695 59805
rect 381494 59800 381695 59802
rect 381494 59744 381634 59800
rect 381690 59744 381695 59800
rect 381494 59742 381695 59744
rect 381629 59739 381695 59742
rect 381799 59530 381859 60044
rect 382631 59666 382691 60044
rect 383101 59666 383167 59669
rect 382631 59664 383167 59666
rect 382631 59608 383106 59664
rect 383162 59608 383167 59664
rect 382631 59606 383167 59608
rect 383462 59666 383522 60044
rect 384113 59666 384179 59669
rect 383462 59664 384179 59666
rect 383462 59608 384118 59664
rect 384174 59608 384179 59664
rect 383462 59606 384179 59608
rect 383101 59603 383167 59606
rect 384113 59603 384179 59606
rect 383929 59530 383995 59533
rect 380758 59470 381738 59530
rect 381799 59528 383995 59530
rect 381799 59472 383934 59528
rect 383990 59472 383995 59528
rect 381799 59470 383995 59472
rect 381678 59394 381738 59470
rect 383929 59467 383995 59470
rect 382365 59394 382431 59397
rect 381678 59392 382431 59394
rect 381678 59336 382370 59392
rect 382426 59336 382431 59392
rect 381678 59334 382431 59336
rect 382365 59331 382431 59334
rect 383101 59394 383167 59397
rect 384294 59394 384354 60044
rect 385126 59530 385186 60044
rect 385769 59530 385835 59533
rect 385126 59528 385835 59530
rect 385126 59472 385774 59528
rect 385830 59472 385835 59528
rect 385126 59470 385835 59472
rect 385957 59530 386017 60044
rect 386789 59666 386849 60044
rect 387425 59666 387491 59669
rect 386789 59664 387491 59666
rect 386789 59608 387430 59664
rect 387486 59608 387491 59664
rect 386789 59606 387491 59608
rect 387620 59666 387680 60044
rect 387620 59606 388362 59666
rect 387425 59603 387491 59606
rect 387977 59530 388043 59533
rect 385957 59528 388043 59530
rect 385957 59472 387982 59528
rect 388038 59472 388043 59528
rect 385957 59470 388043 59472
rect 385769 59467 385835 59470
rect 387977 59467 388043 59470
rect 386413 59394 386479 59397
rect 383101 59392 384130 59394
rect 383101 59336 383106 59392
rect 383162 59336 384130 59392
rect 383101 59334 384130 59336
rect 384294 59392 386479 59394
rect 384294 59336 386418 59392
rect 386474 59336 386479 59392
rect 384294 59334 386479 59336
rect 383101 59331 383167 59334
rect 380893 59258 380959 59261
rect 379838 59256 380959 59258
rect 379838 59200 380898 59256
rect 380954 59200 380959 59256
rect 379838 59198 380959 59200
rect 268009 59195 268075 59198
rect 270677 59195 270743 59198
rect 273345 59195 273411 59198
rect 274909 59195 274975 59198
rect 276105 59195 276171 59198
rect 277485 59195 277551 59198
rect 281533 59195 281599 59198
rect 287237 59195 287303 59198
rect 291377 59195 291443 59198
rect 295701 59195 295767 59198
rect 298921 59195 298987 59198
rect 300301 59195 300367 59198
rect 313917 59195 313983 59198
rect 348417 59195 348483 59198
rect 356881 59195 356947 59198
rect 363045 59195 363111 59198
rect 367093 59195 367159 59198
rect 371417 59195 371483 59198
rect 372705 59195 372771 59198
rect 380893 59195 380959 59198
rect 381629 59258 381695 59261
rect 383745 59258 383811 59261
rect 381629 59256 383811 59258
rect 381629 59200 381634 59256
rect 381690 59200 383750 59256
rect 383806 59200 383811 59256
rect 381629 59198 383811 59200
rect 384070 59258 384130 59334
rect 386413 59331 386479 59334
rect 387425 59394 387491 59397
rect 388302 59394 388362 59606
rect 388452 59530 388512 60044
rect 389284 59666 389344 60044
rect 389449 59802 389515 59805
rect 390115 59802 390175 60044
rect 389449 59800 390175 59802
rect 389449 59744 389454 59800
rect 389510 59744 390175 59800
rect 389449 59742 390175 59744
rect 389449 59739 389515 59742
rect 389284 59606 390754 59666
rect 390553 59530 390619 59533
rect 388452 59528 390619 59530
rect 388452 59472 390558 59528
rect 390614 59472 390619 59528
rect 388452 59470 390619 59472
rect 390553 59467 390619 59470
rect 389541 59394 389607 59397
rect 387425 59392 388178 59394
rect 387425 59336 387430 59392
rect 387486 59336 388178 59392
rect 387425 59334 388178 59336
rect 388302 59392 389607 59394
rect 388302 59336 389546 59392
rect 389602 59336 389607 59392
rect 388302 59334 389607 59336
rect 387425 59331 387491 59334
rect 385217 59258 385283 59261
rect 384070 59256 385283 59258
rect 384070 59200 385222 59256
rect 385278 59200 385283 59256
rect 384070 59198 385283 59200
rect 388118 59258 388178 59334
rect 389541 59331 389607 59334
rect 389357 59258 389423 59261
rect 388118 59256 389423 59258
rect 388118 59200 389362 59256
rect 389418 59200 389423 59256
rect 388118 59198 389423 59200
rect 390694 59258 390754 59606
rect 390947 59394 391007 60044
rect 391778 59530 391838 60044
rect 392610 59666 392670 60044
rect 393313 59666 393379 59669
rect 392610 59664 393379 59666
rect 392610 59608 393318 59664
rect 393374 59608 393379 59664
rect 392610 59606 393379 59608
rect 393313 59603 393379 59606
rect 393313 59530 393379 59533
rect 391778 59528 393379 59530
rect 391778 59472 393318 59528
rect 393374 59472 393379 59528
rect 391778 59470 393379 59472
rect 393313 59467 393379 59470
rect 393442 59394 393502 60044
rect 394273 59394 394333 60044
rect 394693 59530 394759 59533
rect 395105 59530 395165 60044
rect 394693 59528 395165 59530
rect 394693 59472 394698 59528
rect 394754 59472 395165 59528
rect 394693 59470 395165 59472
rect 395936 59530 395996 60044
rect 396768 59666 396828 60044
rect 397600 59802 397660 60044
rect 398431 59938 398491 60044
rect 398431 59878 399034 59938
rect 398833 59802 398899 59805
rect 397600 59800 398899 59802
rect 397600 59744 398838 59800
rect 398894 59744 398899 59800
rect 397600 59742 398899 59744
rect 398833 59739 398899 59742
rect 396768 59606 398298 59666
rect 397545 59530 397611 59533
rect 395936 59528 397611 59530
rect 395936 59472 397550 59528
rect 397606 59472 397611 59528
rect 395936 59470 397611 59472
rect 394693 59467 394759 59470
rect 397545 59467 397611 59470
rect 396349 59394 396415 59397
rect 390947 59334 393330 59394
rect 393442 59334 394066 59394
rect 394273 59392 396415 59394
rect 394273 59336 396354 59392
rect 396410 59336 396415 59392
rect 394273 59334 396415 59336
rect 398238 59394 398298 59606
rect 398974 59530 399034 59878
rect 399263 59666 399323 60044
rect 400094 59802 400154 60044
rect 400926 59938 400986 60044
rect 400814 59878 400986 59938
rect 401758 59938 401818 60044
rect 401758 59878 401978 59938
rect 400673 59802 400739 59805
rect 400094 59800 400739 59802
rect 400094 59744 400678 59800
rect 400734 59744 400739 59800
rect 400094 59742 400739 59744
rect 400673 59739 400739 59742
rect 400814 59666 400874 59878
rect 400949 59802 401015 59805
rect 401777 59802 401843 59805
rect 400949 59800 401843 59802
rect 400949 59744 400954 59800
rect 401010 59744 401782 59800
rect 401838 59744 401843 59800
rect 400949 59742 401843 59744
rect 400949 59739 401015 59742
rect 401777 59739 401843 59742
rect 401918 59666 401978 59878
rect 399263 59606 400690 59666
rect 400814 59606 400986 59666
rect 400305 59530 400371 59533
rect 398974 59528 400371 59530
rect 398974 59472 400310 59528
rect 400366 59472 400371 59528
rect 398974 59470 400371 59472
rect 400305 59467 400371 59470
rect 398925 59394 398991 59397
rect 398238 59392 398991 59394
rect 398238 59336 398930 59392
rect 398986 59336 398991 59392
rect 398238 59334 398991 59336
rect 392117 59258 392183 59261
rect 390694 59256 392183 59258
rect 390694 59200 392122 59256
rect 392178 59200 392183 59256
rect 390694 59198 392183 59200
rect 393270 59258 393330 59334
rect 393589 59258 393655 59261
rect 393270 59256 393655 59258
rect 393270 59200 393594 59256
rect 393650 59200 393655 59256
rect 393270 59198 393655 59200
rect 394006 59258 394066 59334
rect 396349 59331 396415 59334
rect 398925 59331 398991 59334
rect 399109 59394 399175 59397
rect 400489 59394 400555 59397
rect 399109 59392 400555 59394
rect 399109 59336 399114 59392
rect 399170 59336 400494 59392
rect 400550 59336 400555 59392
rect 399109 59334 400555 59336
rect 399109 59331 399175 59334
rect 400489 59331 400555 59334
rect 396165 59258 396231 59261
rect 394006 59256 396231 59258
rect 394006 59200 396170 59256
rect 396226 59200 396231 59256
rect 394006 59198 396231 59200
rect 400630 59258 400690 59606
rect 400926 59394 400986 59606
rect 401758 59606 401978 59666
rect 401501 59530 401567 59533
rect 401758 59530 401818 59606
rect 401501 59528 401818 59530
rect 401501 59472 401506 59528
rect 401562 59472 401818 59528
rect 401501 59470 401818 59472
rect 401501 59467 401567 59470
rect 402589 59394 402649 60044
rect 403421 59394 403481 60044
rect 404252 59530 404312 60044
rect 405084 59666 405144 60044
rect 405916 59802 405976 60044
rect 406561 59802 406627 59805
rect 405916 59800 406627 59802
rect 405916 59744 406566 59800
rect 406622 59744 406627 59800
rect 405916 59742 406627 59744
rect 406561 59739 406627 59742
rect 405084 59606 406578 59666
rect 405733 59530 405799 59533
rect 404252 59528 405799 59530
rect 404252 59472 405738 59528
rect 405794 59472 405799 59528
rect 404252 59470 405799 59472
rect 405733 59467 405799 59470
rect 405825 59394 405891 59397
rect 400926 59334 402346 59394
rect 402589 59334 403266 59394
rect 403421 59392 405891 59394
rect 403421 59336 405830 59392
rect 405886 59336 405891 59392
rect 403421 59334 405891 59336
rect 406518 59394 406578 59606
rect 406747 59530 406807 60044
rect 407579 59666 407639 60044
rect 408410 59802 408470 60044
rect 409045 59802 409111 59805
rect 408410 59800 409111 59802
rect 408410 59744 409050 59800
rect 409106 59744 409111 59800
rect 408410 59742 409111 59744
rect 409045 59739 409111 59742
rect 407579 59606 409154 59666
rect 408769 59530 408835 59533
rect 406747 59528 408835 59530
rect 406747 59472 408774 59528
rect 408830 59472 408835 59528
rect 406747 59470 408835 59472
rect 408769 59467 408835 59470
rect 407205 59394 407271 59397
rect 406518 59392 407271 59394
rect 406518 59336 407210 59392
rect 407266 59336 407271 59392
rect 406518 59334 407271 59336
rect 401593 59258 401659 59261
rect 400630 59256 401659 59258
rect 400630 59200 401598 59256
rect 401654 59200 401659 59256
rect 400630 59198 401659 59200
rect 402286 59258 402346 59334
rect 402973 59258 403039 59261
rect 402286 59256 403039 59258
rect 402286 59200 402978 59256
rect 403034 59200 403039 59256
rect 402286 59198 403039 59200
rect 403206 59258 403266 59334
rect 405825 59331 405891 59334
rect 407205 59331 407271 59334
rect 404537 59258 404603 59261
rect 403206 59256 404603 59258
rect 403206 59200 404542 59256
rect 404598 59200 404603 59256
rect 403206 59198 404603 59200
rect 409094 59258 409154 59606
rect 409242 59394 409302 60044
rect 410074 59530 410134 60044
rect 410905 59666 410965 60044
rect 411529 59666 411595 59669
rect 410905 59664 411595 59666
rect 410905 59608 411534 59664
rect 411590 59608 411595 59664
rect 410905 59606 411595 59608
rect 411737 59666 411797 60044
rect 412357 59666 412423 59669
rect 411737 59664 412423 59666
rect 411737 59608 412362 59664
rect 412418 59608 412423 59664
rect 411737 59606 412423 59608
rect 411529 59603 411595 59606
rect 412357 59603 412423 59606
rect 412357 59530 412423 59533
rect 410074 59528 412423 59530
rect 410074 59472 412362 59528
rect 412418 59472 412423 59528
rect 410074 59470 412423 59472
rect 412568 59530 412628 60044
rect 412817 59802 412883 59805
rect 413400 59802 413460 60044
rect 412817 59800 413460 59802
rect 412817 59744 412822 59800
rect 412878 59744 413460 59800
rect 412817 59742 413460 59744
rect 412817 59739 412883 59742
rect 412725 59666 412791 59669
rect 414105 59666 414171 59669
rect 412725 59664 414171 59666
rect 412725 59608 412730 59664
rect 412786 59608 414110 59664
rect 414166 59608 414171 59664
rect 412725 59606 414171 59608
rect 412725 59603 412791 59606
rect 414105 59603 414171 59606
rect 414105 59530 414171 59533
rect 412568 59528 414171 59530
rect 412568 59472 414110 59528
rect 414166 59472 414171 59528
rect 412568 59470 414171 59472
rect 412357 59467 412423 59470
rect 414105 59467 414171 59470
rect 411529 59394 411595 59397
rect 412909 59394 412975 59397
rect 409242 59334 410810 59394
rect 409965 59258 410031 59261
rect 409094 59256 410031 59258
rect 409094 59200 409970 59256
rect 410026 59200 410031 59256
rect 409094 59198 410031 59200
rect 410750 59258 410810 59334
rect 411529 59392 412975 59394
rect 411529 59336 411534 59392
rect 411590 59336 412914 59392
rect 412970 59336 412975 59392
rect 411529 59334 412975 59336
rect 414232 59394 414292 60044
rect 415063 59394 415123 60044
rect 415895 59530 415955 60044
rect 416726 59666 416786 60044
rect 417558 59805 417618 60044
rect 417558 59800 417667 59805
rect 417558 59744 417606 59800
rect 417662 59744 417667 59800
rect 417558 59742 417667 59744
rect 417601 59739 417667 59742
rect 417601 59666 417667 59669
rect 416726 59664 417667 59666
rect 416726 59608 417606 59664
rect 417662 59608 417667 59664
rect 416726 59606 417667 59608
rect 417601 59603 417667 59606
rect 418245 59530 418311 59533
rect 415895 59470 417434 59530
rect 417049 59394 417115 59397
rect 414232 59334 414858 59394
rect 415063 59392 417115 59394
rect 415063 59336 417054 59392
rect 417110 59336 417115 59392
rect 415063 59334 417115 59336
rect 417374 59394 417434 59470
rect 417742 59528 418311 59530
rect 417742 59472 418250 59528
rect 418306 59472 418311 59528
rect 417742 59470 418311 59472
rect 418390 59530 418450 60044
rect 419073 59530 419139 59533
rect 418390 59528 419139 59530
rect 418390 59472 419078 59528
rect 419134 59472 419139 59528
rect 418390 59470 419139 59472
rect 419221 59530 419281 60044
rect 420053 59666 420113 60044
rect 420729 59666 420795 59669
rect 420053 59664 420795 59666
rect 420053 59608 420734 59664
rect 420790 59608 420795 59664
rect 420053 59606 420795 59608
rect 420884 59666 420944 60044
rect 421716 59802 421776 60044
rect 422385 59802 422451 59805
rect 421716 59800 422451 59802
rect 421716 59744 422390 59800
rect 422446 59744 422451 59800
rect 421716 59742 422451 59744
rect 422385 59739 422451 59742
rect 422109 59666 422175 59669
rect 422293 59666 422359 59669
rect 420884 59664 422175 59666
rect 420884 59608 422114 59664
rect 422170 59608 422175 59664
rect 420884 59606 422175 59608
rect 420729 59603 420795 59606
rect 422109 59603 422175 59606
rect 422250 59664 422359 59666
rect 422250 59608 422298 59664
rect 422354 59608 422359 59664
rect 422250 59603 422359 59608
rect 421097 59530 421163 59533
rect 419221 59528 421163 59530
rect 419221 59472 421102 59528
rect 421158 59472 421163 59528
rect 419221 59470 421163 59472
rect 417742 59394 417802 59470
rect 418245 59467 418311 59470
rect 419073 59467 419139 59470
rect 421097 59467 421163 59470
rect 417374 59334 417802 59394
rect 420729 59394 420795 59397
rect 422250 59394 422310 59603
rect 420729 59392 422310 59394
rect 420729 59336 420734 59392
rect 420790 59336 422310 59392
rect 420729 59334 422310 59336
rect 422548 59394 422608 60044
rect 423379 59530 423439 60044
rect 424211 59666 424271 60044
rect 425042 59802 425102 60044
rect 425697 59802 425763 59805
rect 425042 59800 425763 59802
rect 425042 59744 425702 59800
rect 425758 59744 425763 59800
rect 425042 59742 425763 59744
rect 425697 59739 425763 59742
rect 424211 59606 425714 59666
rect 425053 59530 425119 59533
rect 423379 59528 425119 59530
rect 423379 59472 425058 59528
rect 425114 59472 425119 59528
rect 423379 59470 425119 59472
rect 425053 59467 425119 59470
rect 425145 59394 425211 59397
rect 422548 59392 425211 59394
rect 422548 59336 425150 59392
rect 425206 59336 425211 59392
rect 422548 59334 425211 59336
rect 425654 59394 425714 59606
rect 425874 59530 425934 60044
rect 426706 59666 426766 60044
rect 427537 59802 427597 60044
rect 428089 59802 428155 59805
rect 427537 59800 428155 59802
rect 427537 59744 428094 59800
rect 428150 59744 428155 59800
rect 427537 59742 428155 59744
rect 428369 59802 428429 60044
rect 429009 59802 429075 59805
rect 428369 59800 429075 59802
rect 428369 59744 429014 59800
rect 429070 59744 429075 59800
rect 428369 59742 429075 59744
rect 429200 59802 429260 60044
rect 429837 59802 429903 59805
rect 429200 59800 429903 59802
rect 429200 59744 429842 59800
rect 429898 59744 429903 59800
rect 429200 59742 429903 59744
rect 428089 59739 428155 59742
rect 429009 59739 429075 59742
rect 429837 59739 429903 59742
rect 429193 59666 429259 59669
rect 426706 59664 429259 59666
rect 426706 59608 429198 59664
rect 429254 59608 429259 59664
rect 426706 59606 429259 59608
rect 430032 59666 430092 60044
rect 430573 59666 430639 59669
rect 430032 59664 430639 59666
rect 430032 59608 430578 59664
rect 430634 59608 430639 59664
rect 430032 59606 430639 59608
rect 429193 59603 429259 59606
rect 430573 59603 430639 59606
rect 428181 59530 428247 59533
rect 425874 59528 428247 59530
rect 425874 59472 428186 59528
rect 428242 59472 428247 59528
rect 425874 59470 428247 59472
rect 428181 59467 428247 59470
rect 429009 59530 429075 59533
rect 430665 59530 430731 59533
rect 429009 59528 430731 59530
rect 429009 59472 429014 59528
rect 429070 59472 430670 59528
rect 430726 59472 430731 59528
rect 429009 59470 430731 59472
rect 430864 59530 430924 60044
rect 431695 59666 431755 60044
rect 431695 59606 432338 59666
rect 431769 59530 431835 59533
rect 430864 59528 431835 59530
rect 430864 59472 431774 59528
rect 431830 59472 431835 59528
rect 430864 59470 431835 59472
rect 429009 59467 429075 59470
rect 430665 59467 430731 59470
rect 431769 59467 431835 59470
rect 426525 59394 426591 59397
rect 425654 59392 426591 59394
rect 425654 59336 426530 59392
rect 426586 59336 426591 59392
rect 425654 59334 426591 59336
rect 411529 59331 411595 59334
rect 412909 59331 412975 59334
rect 411253 59258 411319 59261
rect 410750 59256 411319 59258
rect 410750 59200 411258 59256
rect 411314 59200 411319 59256
rect 410750 59198 411319 59200
rect 414798 59258 414858 59334
rect 417049 59331 417115 59334
rect 420729 59331 420795 59334
rect 425145 59331 425211 59334
rect 426525 59331 426591 59334
rect 428089 59394 428155 59397
rect 429285 59394 429351 59397
rect 428089 59392 429351 59394
rect 428089 59336 428094 59392
rect 428150 59336 429290 59392
rect 429346 59336 429351 59392
rect 428089 59334 429351 59336
rect 428089 59331 428155 59334
rect 429285 59331 429351 59334
rect 430573 59394 430639 59397
rect 432137 59394 432203 59397
rect 430573 59392 432203 59394
rect 430573 59336 430578 59392
rect 430634 59336 432142 59392
rect 432198 59336 432203 59392
rect 430573 59334 432203 59336
rect 432278 59394 432338 59606
rect 432527 59530 432587 60044
rect 433358 59666 433418 60044
rect 433977 59666 434043 59669
rect 433358 59664 434043 59666
rect 433358 59608 433982 59664
rect 434038 59608 434043 59664
rect 433358 59606 434043 59608
rect 434190 59666 434250 60044
rect 435022 59802 435082 60044
rect 435853 59938 435913 60044
rect 436685 59938 436745 60044
rect 435853 59878 436570 59938
rect 436685 59878 437122 59938
rect 435817 59802 435883 59805
rect 435022 59800 435883 59802
rect 435022 59744 435822 59800
rect 435878 59744 435883 59800
rect 435022 59742 435883 59744
rect 435817 59739 435883 59742
rect 434190 59606 435650 59666
rect 433977 59603 434043 59606
rect 434805 59530 434871 59533
rect 432527 59528 434871 59530
rect 432527 59472 434810 59528
rect 434866 59472 434871 59528
rect 432527 59470 434871 59472
rect 434805 59467 434871 59470
rect 433517 59394 433583 59397
rect 432278 59392 433583 59394
rect 432278 59336 433522 59392
rect 433578 59336 433583 59392
rect 432278 59334 433583 59336
rect 430573 59331 430639 59334
rect 432137 59331 432203 59334
rect 433517 59331 433583 59334
rect 433977 59394 434043 59397
rect 435590 59394 435650 59606
rect 436510 59530 436570 59878
rect 437062 59666 437122 59878
rect 437516 59802 437576 60044
rect 438209 59802 438275 59805
rect 437516 59800 438275 59802
rect 437516 59744 438214 59800
rect 438270 59744 438275 59800
rect 437516 59742 438275 59744
rect 438348 59802 438408 60044
rect 438761 59802 438827 59805
rect 438348 59800 438827 59802
rect 438348 59744 438766 59800
rect 438822 59744 438827 59800
rect 438348 59742 438827 59744
rect 438209 59739 438275 59742
rect 438761 59739 438827 59742
rect 439180 59666 439240 60044
rect 440011 59802 440071 60044
rect 440693 59802 440759 59805
rect 440011 59800 440759 59802
rect 440011 59744 440698 59800
rect 440754 59744 440759 59800
rect 440011 59742 440759 59744
rect 440843 59802 440903 60044
rect 441245 59802 441311 59805
rect 440843 59800 441311 59802
rect 440843 59744 441250 59800
rect 441306 59744 441311 59800
rect 440843 59742 441311 59744
rect 441674 59802 441734 60044
rect 442349 59802 442415 59805
rect 441674 59800 442415 59802
rect 441674 59744 442354 59800
rect 442410 59744 442415 59800
rect 441674 59742 442415 59744
rect 440693 59739 440759 59742
rect 441245 59739 441311 59742
rect 442349 59739 442415 59742
rect 442257 59666 442323 59669
rect 437062 59606 438962 59666
rect 439180 59606 439882 59666
rect 438117 59530 438183 59533
rect 436510 59528 438183 59530
rect 436510 59472 438122 59528
rect 438178 59472 438183 59528
rect 436510 59470 438183 59472
rect 438902 59530 438962 59606
rect 439497 59530 439563 59533
rect 438902 59528 439563 59530
rect 438902 59472 439502 59528
rect 439558 59472 439563 59528
rect 438902 59470 439563 59472
rect 439822 59530 439882 59606
rect 440374 59664 442323 59666
rect 440374 59608 442262 59664
rect 442318 59608 442323 59664
rect 440374 59606 442323 59608
rect 440374 59530 440434 59606
rect 442257 59603 442323 59606
rect 439822 59470 440434 59530
rect 440693 59530 440759 59533
rect 442349 59530 442415 59533
rect 440693 59528 442415 59530
rect 440693 59472 440698 59528
rect 440754 59472 442354 59528
rect 442410 59472 442415 59528
rect 440693 59470 442415 59472
rect 442506 59530 442566 60044
rect 443338 59666 443398 60044
rect 444005 59666 444071 59669
rect 443338 59664 444071 59666
rect 443338 59608 444010 59664
rect 444066 59608 444071 59664
rect 443338 59606 444071 59608
rect 444169 59666 444229 60044
rect 445001 59802 445061 60044
rect 445661 59802 445727 59805
rect 445001 59800 445727 59802
rect 445001 59744 445666 59800
rect 445722 59744 445727 59800
rect 445001 59742 445727 59744
rect 445661 59739 445727 59742
rect 445661 59666 445727 59669
rect 444169 59664 445727 59666
rect 444169 59608 445666 59664
rect 445722 59608 445727 59664
rect 444169 59606 445727 59608
rect 444005 59603 444071 59606
rect 445661 59603 445727 59606
rect 445017 59530 445083 59533
rect 442506 59528 445083 59530
rect 442506 59472 445022 59528
rect 445078 59472 445083 59528
rect 442506 59470 445083 59472
rect 445832 59530 445892 60044
rect 446397 59530 446463 59533
rect 445832 59528 446463 59530
rect 445832 59472 446402 59528
rect 446458 59472 446463 59528
rect 445832 59470 446463 59472
rect 438117 59467 438183 59470
rect 439497 59467 439563 59470
rect 440693 59467 440759 59470
rect 442349 59467 442415 59470
rect 445017 59467 445083 59470
rect 446397 59467 446463 59470
rect 436737 59394 436803 59397
rect 433977 59392 435466 59394
rect 433977 59336 433982 59392
rect 434038 59336 435466 59392
rect 433977 59334 435466 59336
rect 435590 59392 436803 59394
rect 435590 59336 436742 59392
rect 436798 59336 436803 59392
rect 435590 59334 436803 59336
rect 433977 59331 434043 59334
rect 416865 59258 416931 59261
rect 414798 59256 416931 59258
rect 414798 59200 416870 59256
rect 416926 59200 416931 59256
rect 414798 59198 416931 59200
rect 435406 59258 435466 59334
rect 436737 59331 436803 59334
rect 438761 59394 438827 59397
rect 441061 59394 441127 59397
rect 438761 59392 441127 59394
rect 438761 59336 438766 59392
rect 438822 59336 441066 59392
rect 441122 59336 441127 59392
rect 438761 59334 441127 59336
rect 438761 59331 438827 59334
rect 441061 59331 441127 59334
rect 441245 59394 441311 59397
rect 443637 59394 443703 59397
rect 441245 59392 443703 59394
rect 441245 59336 441250 59392
rect 441306 59336 443642 59392
rect 443698 59336 443703 59392
rect 441245 59334 443703 59336
rect 441245 59331 441311 59334
rect 443637 59331 443703 59334
rect 444005 59394 444071 59397
rect 446397 59394 446463 59397
rect 444005 59392 446463 59394
rect 444005 59336 444010 59392
rect 444066 59336 446402 59392
rect 446458 59336 446463 59392
rect 444005 59334 446463 59336
rect 446664 59394 446724 60044
rect 447496 59530 447556 60044
rect 448145 59530 448211 59533
rect 447496 59528 448211 59530
rect 447496 59472 448150 59528
rect 448206 59472 448211 59528
rect 447496 59470 448211 59472
rect 448327 59530 448387 60044
rect 449159 59666 449219 60044
rect 449990 59802 450050 60044
rect 450537 59802 450603 59805
rect 449990 59800 450603 59802
rect 449990 59744 450542 59800
rect 450598 59744 450603 59800
rect 449990 59742 450603 59744
rect 450537 59739 450603 59742
rect 450629 59666 450695 59669
rect 449159 59664 450695 59666
rect 449159 59608 450634 59664
rect 450690 59608 450695 59664
rect 449159 59606 450695 59608
rect 450629 59603 450695 59606
rect 450445 59530 450511 59533
rect 448327 59528 450511 59530
rect 448327 59472 450450 59528
rect 450506 59472 450511 59528
rect 448327 59470 450511 59472
rect 448145 59467 448211 59470
rect 450445 59467 450511 59470
rect 449157 59394 449223 59397
rect 446664 59392 449223 59394
rect 446664 59336 449162 59392
rect 449218 59336 449223 59392
rect 446664 59334 449223 59336
rect 444005 59331 444071 59334
rect 446397 59331 446463 59334
rect 449157 59331 449223 59334
rect 450537 59394 450603 59397
rect 450822 59394 450882 60044
rect 451654 59530 451714 60044
rect 452285 59530 452351 59533
rect 451654 59528 452351 59530
rect 451654 59472 452290 59528
rect 452346 59472 452351 59528
rect 451654 59470 452351 59472
rect 452485 59530 452545 60044
rect 453317 59666 453377 60044
rect 454148 59802 454208 60044
rect 454769 59802 454835 59805
rect 454148 59800 454835 59802
rect 454148 59744 454774 59800
rect 454830 59744 454835 59800
rect 454148 59742 454835 59744
rect 454980 59802 455040 60044
rect 455597 59802 455663 59805
rect 454980 59800 455663 59802
rect 454980 59744 455602 59800
rect 455658 59744 455663 59800
rect 454980 59742 455663 59744
rect 455812 59802 455872 60044
rect 456517 59802 456583 59805
rect 455812 59800 456583 59802
rect 455812 59744 456522 59800
rect 456578 59744 456583 59800
rect 455812 59742 456583 59744
rect 454769 59739 454835 59742
rect 455597 59739 455663 59742
rect 456517 59739 456583 59742
rect 456057 59666 456123 59669
rect 453317 59664 456123 59666
rect 453317 59608 456062 59664
rect 456118 59608 456123 59664
rect 453317 59606 456123 59608
rect 456057 59603 456123 59606
rect 454677 59530 454743 59533
rect 452485 59528 454743 59530
rect 452485 59472 454682 59528
rect 454738 59472 454743 59528
rect 452485 59470 454743 59472
rect 456643 59530 456703 60044
rect 457475 59666 457535 60044
rect 458173 59666 458239 59669
rect 457475 59664 458239 59666
rect 457475 59608 458178 59664
rect 458234 59608 458239 59664
rect 457475 59606 458239 59608
rect 458306 59666 458366 60044
rect 458909 59666 458975 59669
rect 458306 59664 458975 59666
rect 458306 59608 458914 59664
rect 458970 59608 458975 59664
rect 458306 59606 458975 59608
rect 458173 59603 458239 59606
rect 458909 59603 458975 59606
rect 459001 59530 459067 59533
rect 456643 59528 459067 59530
rect 456643 59472 459006 59528
rect 459062 59472 459067 59528
rect 456643 59470 459067 59472
rect 459138 59530 459198 60044
rect 459970 59666 460030 60044
rect 460801 59802 460861 60044
rect 461485 59802 461551 59805
rect 460801 59800 461551 59802
rect 460801 59744 461490 59800
rect 461546 59744 461551 59800
rect 460801 59742 461551 59744
rect 461485 59739 461551 59742
rect 460473 59666 460539 59669
rect 459970 59664 460539 59666
rect 459970 59608 460478 59664
rect 460534 59608 460539 59664
rect 459970 59606 460539 59608
rect 460473 59603 460539 59606
rect 461485 59530 461551 59533
rect 459138 59528 461551 59530
rect 459138 59472 461490 59528
rect 461546 59472 461551 59528
rect 459138 59470 461551 59472
rect 452285 59467 452351 59470
rect 454677 59467 454743 59470
rect 459001 59467 459067 59470
rect 461485 59467 461551 59470
rect 451273 59394 451339 59397
rect 453297 59394 453363 59397
rect 450537 59392 450738 59394
rect 450537 59336 450542 59392
rect 450598 59336 450738 59392
rect 450537 59334 450738 59336
rect 450822 59392 451339 59394
rect 450822 59336 451278 59392
rect 451334 59336 451339 59392
rect 450822 59334 451339 59336
rect 450537 59331 450603 59334
rect 436093 59258 436159 59261
rect 435406 59256 436159 59258
rect 435406 59200 436098 59256
rect 436154 59200 436159 59256
rect 435406 59198 436159 59200
rect 381629 59195 381695 59198
rect 383745 59195 383811 59198
rect 385217 59195 385283 59198
rect 389357 59195 389423 59198
rect 392117 59195 392183 59198
rect 393589 59195 393655 59198
rect 396165 59195 396231 59198
rect 401593 59195 401659 59198
rect 402973 59195 403039 59198
rect 404537 59195 404603 59198
rect 409965 59195 410031 59198
rect 411253 59195 411319 59198
rect 416865 59195 416931 59198
rect 436093 59195 436159 59198
rect 262029 59120 263978 59122
rect 262029 59064 262034 59120
rect 262090 59064 263978 59120
rect 262029 59062 263978 59064
rect 450678 59122 450738 59334
rect 451273 59331 451339 59334
rect 451414 59392 453363 59394
rect 451414 59336 453302 59392
rect 453358 59336 453363 59392
rect 451414 59334 453363 59336
rect 451414 59122 451474 59334
rect 453297 59331 453363 59334
rect 455597 59394 455663 59397
rect 457621 59394 457687 59397
rect 455597 59392 457687 59394
rect 455597 59336 455602 59392
rect 455658 59336 457626 59392
rect 457682 59336 457687 59392
rect 455597 59334 457687 59336
rect 455597 59331 455663 59334
rect 457621 59331 457687 59334
rect 458909 59394 458975 59397
rect 460473 59394 460539 59397
rect 461485 59394 461551 59397
rect 458909 59392 459754 59394
rect 458909 59336 458914 59392
rect 458970 59336 459754 59392
rect 458909 59334 459754 59336
rect 458909 59331 458975 59334
rect 459694 59258 459754 59334
rect 460473 59392 461551 59394
rect 460473 59336 460478 59392
rect 460534 59336 461490 59392
rect 461546 59336 461551 59392
rect 460473 59334 461551 59336
rect 461633 59394 461693 60044
rect 462464 59530 462524 60044
rect 463141 59530 463207 59533
rect 462464 59528 463207 59530
rect 462464 59472 463146 59528
rect 463202 59472 463207 59528
rect 462464 59470 463207 59472
rect 463296 59530 463356 60044
rect 464128 59666 464188 60044
rect 464797 59666 464863 59669
rect 464128 59664 464863 59666
rect 464128 59608 464802 59664
rect 464858 59608 464863 59664
rect 464128 59606 464863 59608
rect 464959 59666 465019 60044
rect 465791 59802 465851 60044
rect 466622 59938 466682 60044
rect 466622 59878 468218 59938
rect 467925 59802 467991 59805
rect 465791 59800 467991 59802
rect 465791 59744 467930 59800
rect 467986 59744 467991 59800
rect 465791 59742 467991 59744
rect 467925 59739 467991 59742
rect 467097 59666 467163 59669
rect 464959 59664 467163 59666
rect 464959 59608 467102 59664
rect 467158 59608 467163 59664
rect 464959 59606 467163 59608
rect 464797 59603 464863 59606
rect 467097 59603 467163 59606
rect 465717 59530 465783 59533
rect 463296 59528 465783 59530
rect 463296 59472 465722 59528
rect 465778 59472 465783 59528
rect 463296 59470 465783 59472
rect 463141 59467 463207 59470
rect 465717 59467 465783 59470
rect 464337 59394 464403 59397
rect 461633 59392 464403 59394
rect 461633 59336 464342 59392
rect 464398 59336 464403 59392
rect 461633 59334 464403 59336
rect 460473 59331 460539 59334
rect 461485 59331 461551 59334
rect 464337 59331 464403 59334
rect 464797 59394 464863 59397
rect 467281 59394 467347 59397
rect 464797 59392 467347 59394
rect 464797 59336 464802 59392
rect 464858 59336 467286 59392
rect 467342 59336 467347 59392
rect 464797 59334 467347 59336
rect 464797 59331 464863 59334
rect 467281 59331 467347 59334
rect 461761 59258 461827 59261
rect 459694 59256 461827 59258
rect 459694 59200 461766 59256
rect 461822 59200 461827 59256
rect 459694 59198 461827 59200
rect 468158 59258 468218 59878
rect 468286 59394 468346 60044
rect 469117 59530 469177 60044
rect 469600 59666 469660 60044
rect 472617 59666 472683 59669
rect 469600 59664 472683 59666
rect 469600 59608 472622 59664
rect 472678 59608 472683 59664
rect 469600 59606 472683 59608
rect 472617 59603 472683 59606
rect 471421 59530 471487 59533
rect 469117 59528 471487 59530
rect 469117 59472 471426 59528
rect 471482 59472 471487 59528
rect 583520 59516 584960 59756
rect 469117 59470 471487 59472
rect 471421 59467 471487 59470
rect 471237 59394 471303 59397
rect 468286 59392 471303 59394
rect 468286 59336 471242 59392
rect 471298 59336 471303 59392
rect 468286 59334 471303 59336
rect 471237 59331 471303 59334
rect 470133 59258 470199 59261
rect 468158 59256 470199 59258
rect 468158 59200 470138 59256
rect 470194 59200 470199 59256
rect 468158 59198 470199 59200
rect 461761 59195 461827 59198
rect 470133 59195 470199 59198
rect 450678 59062 451474 59122
rect 61377 59059 61443 59062
rect 72417 59059 72483 59062
rect 130377 59059 130443 59062
rect 208301 59059 208367 59062
rect 217685 59059 217751 59062
rect 262029 59059 262095 59062
rect 141601 58986 141667 58989
rect 144126 58986 144132 58988
rect 141601 58984 144132 58986
rect 141601 58928 141606 58984
rect 141662 58928 144132 58984
rect 141601 58926 144132 58928
rect 141601 58923 141667 58926
rect 144126 58924 144132 58926
rect 144196 58924 144202 58988
rect 350758 58924 350764 58988
rect 350828 58986 350834 58988
rect 352741 58986 352807 58989
rect 350828 58984 352807 58986
rect 350828 58928 352746 58984
rect 352802 58928 352807 58984
rect 350828 58926 352807 58928
rect 350828 58924 350834 58926
rect 352741 58923 352807 58926
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
rect 419625 3634 419691 3637
rect 412590 3632 419691 3634
rect 412590 3576 419630 3632
rect 419686 3576 419691 3632
rect 412590 3574 419691 3576
rect 5257 3362 5323 3365
rect 144177 3362 144243 3365
rect 5257 3360 144243 3362
rect 5257 3304 5262 3360
rect 5318 3304 144182 3360
rect 144238 3304 144243 3360
rect 5257 3302 144243 3304
rect 5257 3299 5323 3302
rect 144177 3299 144243 3302
rect 369393 3362 369459 3365
rect 412590 3362 412650 3574
rect 419625 3571 419691 3574
rect 369393 3360 412650 3362
rect 369393 3304 369398 3360
rect 369454 3304 412650 3360
rect 369393 3302 412650 3304
rect 471421 3362 471487 3365
rect 583385 3362 583451 3365
rect 471421 3360 583451 3362
rect 471421 3304 471426 3360
rect 471482 3304 583390 3360
rect 583446 3304 583451 3360
rect 471421 3302 583451 3304
rect 369393 3299 369459 3302
rect 471421 3299 471487 3302
rect 583385 3299 583451 3302
<< via3 >>
rect 144132 59740 144196 59804
rect 350764 59740 350828 59804
rect 144132 58924 144196 58988
rect 350764 58924 350828 58988
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 451980 60134 456618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 451980 63854 460338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 451980 67574 464058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 451980 74414 470898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 451980 78134 474618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 451980 81854 478338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 451980 85574 482058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 451980 92414 452898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 451980 96134 456618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 451980 99854 460338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 451980 103574 464058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 451980 110414 470898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 451980 114134 474618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 451980 117854 478338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 451980 121574 482058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 451980 128414 452898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 451980 132134 456618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 451980 135854 460338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 451980 139574 464058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 451980 146414 470898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 451980 150134 474618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 451980 153854 478338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 451980 157574 482058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 451980 164414 452898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 451980 168134 456618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 451980 171854 460338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 451980 175574 464058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 451980 182414 470898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 451980 186134 474618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 451980 189854 478338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 451980 193574 482058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 451980 200414 452898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 451980 204134 456618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 451980 207854 460338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 451980 211574 464058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 451980 218414 470898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 451980 222134 474618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 451980 225854 478338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 451980 229574 482058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 451980 236414 452898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 451980 240134 456618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 451980 243854 460338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 451980 247574 464058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 451980 254414 470898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 451980 258134 474618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 451980 261854 478338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 451980 265574 482058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 451980 272414 452898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 451980 276134 456618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 451980 279854 460338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 451980 283574 464058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 451980 290414 470898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 451980 294134 474618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 451980 297854 478338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 451980 301574 482058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 451980 308414 452898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 451980 312134 456618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 451980 315854 460338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 451980 319574 464058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 451980 326414 470898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 451980 330134 474618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 451980 333854 478338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 451980 337574 482058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 451980 344414 452898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 451980 348134 456618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 451980 351854 460338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 451980 355574 464058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 451980 362414 470898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 451980 366134 474618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 451980 369854 478338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 451980 373574 482058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 451980 380414 452898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 451980 384134 456618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 451980 387854 460338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 451980 391574 464058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 451980 398414 470898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 451980 402134 474618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 451980 405854 478338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 451980 409574 482058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 451980 416414 452898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 451980 420134 456618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 451980 423854 460338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 451980 427574 464058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 451980 434414 470898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 451980 438134 474618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 451980 441854 478338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 451980 445574 482058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 451980 452414 452898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 451980 456134 456618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 451980 459854 460338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 451980 463574 464058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 451980 470414 470898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 144131 59804 144197 59805
rect 144131 59740 144132 59804
rect 144196 59740 144197 59804
rect 144131 59739 144197 59740
rect 350763 59804 350829 59805
rect 350763 59740 350764 59804
rect 350828 59740 350829 59804
rect 350763 59739 350829 59740
rect 144134 58989 144194 59739
rect 350766 58989 350826 59739
rect 144131 58988 144197 58989
rect 144131 58924 144132 58988
rect 144196 58924 144197 58988
rect 144131 58923 144197 58924
rect 350763 58988 350829 58989
rect 350763 58924 350764 58988
rect 350828 58924 350829 58988
rect 350763 58923 350829 58924
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 58000
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 28894 63854 58000
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 32614 67574 58000
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 39454 74414 58000
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 43174 78134 58000
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 46894 81854 58000
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 50614 85574 58000
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 58000
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 58000
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 28894 99854 58000
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 32614 103574 58000
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 39454 110414 58000
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 43174 114134 58000
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 46894 117854 58000
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 50614 121574 58000
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 58000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 58000
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 28894 135854 58000
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 32614 139574 58000
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 39454 146414 58000
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 43174 150134 58000
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 46894 153854 58000
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 50614 157574 58000
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 57454 164414 58000
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 25174 168134 58000
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 28894 171854 58000
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 32614 175574 58000
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 39454 182414 58000
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 43174 186134 58000
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 46894 189854 58000
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 50614 193574 58000
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 57454 200414 58000
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 58000
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 28894 207854 58000
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 32614 211574 58000
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 39454 218414 58000
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 43174 222134 58000
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 46894 225854 58000
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 50614 229574 58000
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 57454 236414 58000
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 58000
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 28894 243854 58000
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 32614 247574 58000
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 39454 254414 58000
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 43174 258134 58000
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 46894 261854 58000
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 50614 265574 58000
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 57454 272414 58000
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 25174 276134 58000
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 28894 279854 58000
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 32614 283574 58000
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 39454 290414 58000
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 43174 294134 58000
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 46894 297854 58000
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 50614 301574 58000
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 57454 308414 58000
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 25174 312134 58000
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 28894 315854 58000
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 32614 319574 58000
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 39454 326414 58000
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 43174 330134 58000
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 46894 333854 58000
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 50614 337574 58000
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 57454 344414 58000
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 25174 348134 58000
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 28894 351854 58000
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 32614 355574 58000
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 39454 362414 58000
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 43174 366134 58000
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 46894 369854 58000
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 50614 373574 58000
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 57454 380414 58000
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 25174 384134 58000
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 28894 387854 58000
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 32614 391574 58000
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 39454 398414 58000
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 43174 402134 58000
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 46894 405854 58000
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 50614 409574 58000
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 57454 416414 58000
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 25174 420134 58000
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 28894 423854 58000
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 32614 427574 58000
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 39454 434414 58000
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 43174 438134 58000
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 46894 441854 58000
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 50614 445574 58000
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 57454 452414 58000
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 25174 456134 58000
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 28894 459854 58000
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 32614 463574 58000
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 39454 470414 58000
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 58000 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 58000 446614
rect -8726 446294 58000 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 58000 446294
rect -8726 446026 58000 446058
rect 472044 446614 592650 446646
rect 472044 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect 472044 446294 592650 446378
rect 472044 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect 472044 446026 592650 446058
rect -6806 442894 58000 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 58000 442894
rect -6806 442574 58000 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 58000 442574
rect -6806 442306 58000 442338
rect 472044 442894 590730 442926
rect 472044 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect 472044 442574 590730 442658
rect 472044 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect 472044 442306 590730 442338
rect -4886 439174 58000 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 58000 439174
rect -4886 438854 58000 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 58000 438854
rect -4886 438586 58000 438618
rect 472044 439174 588810 439206
rect 472044 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect 472044 438854 588810 438938
rect 472044 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect 472044 438586 588810 438618
rect -2966 435454 58000 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 58000 435454
rect -2966 435134 58000 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 58000 435134
rect -2966 434866 58000 434898
rect 472044 435454 586890 435486
rect 472044 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect 472044 435134 586890 435218
rect 472044 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect 472044 434866 586890 434898
rect -8726 428614 58000 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 58000 428614
rect -8726 428294 58000 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 58000 428294
rect -8726 428026 58000 428058
rect 472044 428614 592650 428646
rect 472044 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 472044 428294 592650 428378
rect 472044 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 472044 428026 592650 428058
rect -6806 424894 58000 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 58000 424894
rect -6806 424574 58000 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 58000 424574
rect -6806 424306 58000 424338
rect 472044 424894 590730 424926
rect 472044 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 472044 424574 590730 424658
rect 472044 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 472044 424306 590730 424338
rect -4886 421174 58000 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 58000 421174
rect -4886 420854 58000 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 58000 420854
rect -4886 420586 58000 420618
rect 472044 421174 588810 421206
rect 472044 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 472044 420854 588810 420938
rect 472044 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 472044 420586 588810 420618
rect -2966 417454 58000 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 58000 417454
rect -2966 417134 58000 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 58000 417134
rect -2966 416866 58000 416898
rect 472044 417454 586890 417486
rect 472044 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 472044 417134 586890 417218
rect 472044 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 472044 416866 586890 416898
rect -8726 410614 58000 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 58000 410614
rect -8726 410294 58000 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 58000 410294
rect -8726 410026 58000 410058
rect 472044 410614 592650 410646
rect 472044 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect 472044 410294 592650 410378
rect 472044 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect 472044 410026 592650 410058
rect -6806 406894 58000 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 58000 406894
rect -6806 406574 58000 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 58000 406574
rect -6806 406306 58000 406338
rect 472044 406894 590730 406926
rect 472044 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect 472044 406574 590730 406658
rect 472044 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect 472044 406306 590730 406338
rect -4886 403174 58000 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 58000 403174
rect -4886 402854 58000 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 58000 402854
rect -4886 402586 58000 402618
rect 472044 403174 588810 403206
rect 472044 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect 472044 402854 588810 402938
rect 472044 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect 472044 402586 588810 402618
rect -2966 399454 58000 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 58000 399454
rect -2966 399134 58000 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 58000 399134
rect -2966 398866 58000 398898
rect 472044 399454 586890 399486
rect 472044 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect 472044 399134 586890 399218
rect 472044 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect 472044 398866 586890 398898
rect -8726 392614 58000 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 58000 392614
rect -8726 392294 58000 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 58000 392294
rect -8726 392026 58000 392058
rect 472044 392614 592650 392646
rect 472044 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 472044 392294 592650 392378
rect 472044 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 472044 392026 592650 392058
rect -6806 388894 58000 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 58000 388894
rect -6806 388574 58000 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 58000 388574
rect -6806 388306 58000 388338
rect 472044 388894 590730 388926
rect 472044 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 472044 388574 590730 388658
rect 472044 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 472044 388306 590730 388338
rect -4886 385174 58000 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 58000 385174
rect -4886 384854 58000 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 58000 384854
rect -4886 384586 58000 384618
rect 472044 385174 588810 385206
rect 472044 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 472044 384854 588810 384938
rect 472044 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 472044 384586 588810 384618
rect -2966 381454 58000 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 58000 381454
rect -2966 381134 58000 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 58000 381134
rect -2966 380866 58000 380898
rect 472044 381454 586890 381486
rect 472044 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 472044 381134 586890 381218
rect 472044 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 472044 380866 586890 380898
rect -8726 374614 58000 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 58000 374614
rect -8726 374294 58000 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 58000 374294
rect -8726 374026 58000 374058
rect 472044 374614 592650 374646
rect 472044 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect 472044 374294 592650 374378
rect 472044 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect 472044 374026 592650 374058
rect -6806 370894 58000 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 58000 370894
rect -6806 370574 58000 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 58000 370574
rect -6806 370306 58000 370338
rect 472044 370894 590730 370926
rect 472044 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect 472044 370574 590730 370658
rect 472044 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect 472044 370306 590730 370338
rect -4886 367174 58000 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 58000 367174
rect -4886 366854 58000 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 58000 366854
rect -4886 366586 58000 366618
rect 472044 367174 588810 367206
rect 472044 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect 472044 366854 588810 366938
rect 472044 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect 472044 366586 588810 366618
rect -2966 363454 58000 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 58000 363454
rect -2966 363134 58000 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 58000 363134
rect -2966 362866 58000 362898
rect 472044 363454 586890 363486
rect 472044 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect 472044 363134 586890 363218
rect 472044 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect 472044 362866 586890 362898
rect -8726 356614 58000 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 58000 356614
rect -8726 356294 58000 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 58000 356294
rect -8726 356026 58000 356058
rect 472044 356614 592650 356646
rect 472044 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 472044 356294 592650 356378
rect 472044 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 472044 356026 592650 356058
rect -6806 352894 58000 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 58000 352894
rect -6806 352574 58000 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 58000 352574
rect -6806 352306 58000 352338
rect 472044 352894 590730 352926
rect 472044 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 472044 352574 590730 352658
rect 472044 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 472044 352306 590730 352338
rect -4886 349174 58000 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 58000 349174
rect -4886 348854 58000 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 58000 348854
rect -4886 348586 58000 348618
rect 472044 349174 588810 349206
rect 472044 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 472044 348854 588810 348938
rect 472044 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 472044 348586 588810 348618
rect -2966 345454 58000 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 58000 345454
rect -2966 345134 58000 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 58000 345134
rect -2966 344866 58000 344898
rect 472044 345454 586890 345486
rect 472044 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 472044 345134 586890 345218
rect 472044 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 472044 344866 586890 344898
rect -8726 338614 58000 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 58000 338614
rect -8726 338294 58000 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 58000 338294
rect -8726 338026 58000 338058
rect 472044 338614 592650 338646
rect 472044 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect 472044 338294 592650 338378
rect 472044 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect 472044 338026 592650 338058
rect -6806 334894 58000 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 58000 334894
rect -6806 334574 58000 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 58000 334574
rect -6806 334306 58000 334338
rect 472044 334894 590730 334926
rect 472044 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect 472044 334574 590730 334658
rect 472044 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect 472044 334306 590730 334338
rect -4886 331174 58000 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 58000 331174
rect -4886 330854 58000 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 58000 330854
rect -4886 330586 58000 330618
rect 472044 331174 588810 331206
rect 472044 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect 472044 330854 588810 330938
rect 472044 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect 472044 330586 588810 330618
rect -2966 327454 58000 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 58000 327454
rect -2966 327134 58000 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 58000 327134
rect -2966 326866 58000 326898
rect 472044 327454 586890 327486
rect 472044 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect 472044 327134 586890 327218
rect 472044 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect 472044 326866 586890 326898
rect -8726 320614 58000 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 58000 320614
rect -8726 320294 58000 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 58000 320294
rect -8726 320026 58000 320058
rect 472044 320614 592650 320646
rect 472044 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 472044 320294 592650 320378
rect 472044 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 472044 320026 592650 320058
rect -6806 316894 58000 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 58000 316894
rect -6806 316574 58000 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 58000 316574
rect -6806 316306 58000 316338
rect 472044 316894 590730 316926
rect 472044 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 472044 316574 590730 316658
rect 472044 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 472044 316306 590730 316338
rect -4886 313174 58000 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 58000 313174
rect -4886 312854 58000 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 58000 312854
rect -4886 312586 58000 312618
rect 472044 313174 588810 313206
rect 472044 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 472044 312854 588810 312938
rect 472044 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 472044 312586 588810 312618
rect -2966 309454 58000 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 58000 309454
rect -2966 309134 58000 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 58000 309134
rect -2966 308866 58000 308898
rect 472044 309454 586890 309486
rect 472044 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 472044 309134 586890 309218
rect 472044 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 472044 308866 586890 308898
rect -8726 302614 58000 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 58000 302614
rect -8726 302294 58000 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 58000 302294
rect -8726 302026 58000 302058
rect 472044 302614 592650 302646
rect 472044 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect 472044 302294 592650 302378
rect 472044 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect 472044 302026 592650 302058
rect -6806 298894 58000 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 58000 298894
rect -6806 298574 58000 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 58000 298574
rect -6806 298306 58000 298338
rect 472044 298894 590730 298926
rect 472044 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect 472044 298574 590730 298658
rect 472044 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect 472044 298306 590730 298338
rect -4886 295174 58000 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 58000 295174
rect -4886 294854 58000 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 58000 294854
rect -4886 294586 58000 294618
rect 472044 295174 588810 295206
rect 472044 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect 472044 294854 588810 294938
rect 472044 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect 472044 294586 588810 294618
rect -2966 291454 58000 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 58000 291454
rect -2966 291134 58000 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 58000 291134
rect -2966 290866 58000 290898
rect 472044 291454 586890 291486
rect 472044 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect 472044 291134 586890 291218
rect 472044 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect 472044 290866 586890 290898
rect -8726 284614 58000 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 58000 284614
rect -8726 284294 58000 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 58000 284294
rect -8726 284026 58000 284058
rect 472044 284614 592650 284646
rect 472044 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 472044 284294 592650 284378
rect 472044 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 472044 284026 592650 284058
rect -6806 280894 58000 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 58000 280894
rect -6806 280574 58000 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 58000 280574
rect -6806 280306 58000 280338
rect 472044 280894 590730 280926
rect 472044 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 472044 280574 590730 280658
rect 472044 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 472044 280306 590730 280338
rect -4886 277174 58000 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 58000 277174
rect -4886 276854 58000 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 58000 276854
rect -4886 276586 58000 276618
rect 472044 277174 588810 277206
rect 472044 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 472044 276854 588810 276938
rect 472044 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 472044 276586 588810 276618
rect -2966 273454 58000 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 58000 273454
rect -2966 273134 58000 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 58000 273134
rect -2966 272866 58000 272898
rect 472044 273454 586890 273486
rect 472044 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 472044 273134 586890 273218
rect 472044 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 472044 272866 586890 272898
rect -8726 266614 58000 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 58000 266614
rect -8726 266294 58000 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 58000 266294
rect -8726 266026 58000 266058
rect 472044 266614 592650 266646
rect 472044 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect 472044 266294 592650 266378
rect 472044 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect 472044 266026 592650 266058
rect -6806 262894 58000 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 58000 262894
rect -6806 262574 58000 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 58000 262574
rect -6806 262306 58000 262338
rect 472044 262894 590730 262926
rect 472044 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect 472044 262574 590730 262658
rect 472044 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect 472044 262306 590730 262338
rect -4886 259174 58000 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 58000 259174
rect -4886 258854 58000 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 58000 258854
rect -4886 258586 58000 258618
rect 472044 259174 588810 259206
rect 472044 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect 472044 258854 588810 258938
rect 472044 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect 472044 258586 588810 258618
rect -2966 255454 58000 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 58000 255454
rect -2966 255134 58000 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 58000 255134
rect -2966 254866 58000 254898
rect 472044 255454 586890 255486
rect 472044 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect 472044 255134 586890 255218
rect 472044 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect 472044 254866 586890 254898
rect -8726 248614 58000 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 58000 248614
rect -8726 248294 58000 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 58000 248294
rect -8726 248026 58000 248058
rect 472044 248614 592650 248646
rect 472044 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 472044 248294 592650 248378
rect 472044 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 472044 248026 592650 248058
rect -6806 244894 58000 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 58000 244894
rect -6806 244574 58000 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 58000 244574
rect -6806 244306 58000 244338
rect 472044 244894 590730 244926
rect 472044 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 472044 244574 590730 244658
rect 472044 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 472044 244306 590730 244338
rect -4886 241174 58000 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 58000 241174
rect -4886 240854 58000 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 58000 240854
rect -4886 240586 58000 240618
rect 472044 241174 588810 241206
rect 472044 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 472044 240854 588810 240938
rect 472044 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 472044 240586 588810 240618
rect -2966 237454 58000 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 58000 237454
rect -2966 237134 58000 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 58000 237134
rect -2966 236866 58000 236898
rect 472044 237454 586890 237486
rect 472044 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 472044 237134 586890 237218
rect 472044 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 472044 236866 586890 236898
rect -8726 230614 58000 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 58000 230614
rect -8726 230294 58000 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 58000 230294
rect -8726 230026 58000 230058
rect 472044 230614 592650 230646
rect 472044 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect 472044 230294 592650 230378
rect 472044 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect 472044 230026 592650 230058
rect -6806 226894 58000 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 58000 226894
rect -6806 226574 58000 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 58000 226574
rect -6806 226306 58000 226338
rect 472044 226894 590730 226926
rect 472044 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect 472044 226574 590730 226658
rect 472044 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect 472044 226306 590730 226338
rect -4886 223174 58000 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 58000 223174
rect -4886 222854 58000 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 58000 222854
rect -4886 222586 58000 222618
rect 472044 223174 588810 223206
rect 472044 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect 472044 222854 588810 222938
rect 472044 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect 472044 222586 588810 222618
rect -2966 219454 58000 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 58000 219454
rect -2966 219134 58000 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 58000 219134
rect -2966 218866 58000 218898
rect 472044 219454 586890 219486
rect 472044 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect 472044 219134 586890 219218
rect 472044 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect 472044 218866 586890 218898
rect -8726 212614 58000 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 58000 212614
rect -8726 212294 58000 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 58000 212294
rect -8726 212026 58000 212058
rect 472044 212614 592650 212646
rect 472044 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 472044 212294 592650 212378
rect 472044 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 472044 212026 592650 212058
rect -6806 208894 58000 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 58000 208894
rect -6806 208574 58000 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 58000 208574
rect -6806 208306 58000 208338
rect 472044 208894 590730 208926
rect 472044 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 472044 208574 590730 208658
rect 472044 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 472044 208306 590730 208338
rect -4886 205174 58000 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 58000 205174
rect -4886 204854 58000 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 58000 204854
rect -4886 204586 58000 204618
rect 472044 205174 588810 205206
rect 472044 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 472044 204854 588810 204938
rect 472044 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 472044 204586 588810 204618
rect -2966 201454 58000 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 58000 201454
rect -2966 201134 58000 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 58000 201134
rect -2966 200866 58000 200898
rect 472044 201454 586890 201486
rect 472044 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 472044 201134 586890 201218
rect 472044 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 472044 200866 586890 200898
rect -8726 194614 58000 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 58000 194614
rect -8726 194294 58000 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 58000 194294
rect -8726 194026 58000 194058
rect 472044 194614 592650 194646
rect 472044 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect 472044 194294 592650 194378
rect 472044 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect 472044 194026 592650 194058
rect -6806 190894 58000 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 58000 190894
rect -6806 190574 58000 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 58000 190574
rect -6806 190306 58000 190338
rect 472044 190894 590730 190926
rect 472044 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect 472044 190574 590730 190658
rect 472044 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect 472044 190306 590730 190338
rect -4886 187174 58000 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 58000 187174
rect -4886 186854 58000 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 58000 186854
rect -4886 186586 58000 186618
rect 472044 187174 588810 187206
rect 472044 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect 472044 186854 588810 186938
rect 472044 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect 472044 186586 588810 186618
rect -2966 183454 58000 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 58000 183454
rect -2966 183134 58000 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 58000 183134
rect -2966 182866 58000 182898
rect 472044 183454 586890 183486
rect 472044 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect 472044 183134 586890 183218
rect 472044 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect 472044 182866 586890 182898
rect -8726 176614 58000 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 58000 176614
rect -8726 176294 58000 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 58000 176294
rect -8726 176026 58000 176058
rect 472044 176614 592650 176646
rect 472044 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 472044 176294 592650 176378
rect 472044 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 472044 176026 592650 176058
rect -6806 172894 58000 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 58000 172894
rect -6806 172574 58000 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 58000 172574
rect -6806 172306 58000 172338
rect 472044 172894 590730 172926
rect 472044 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 472044 172574 590730 172658
rect 472044 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 472044 172306 590730 172338
rect -4886 169174 58000 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 58000 169174
rect -4886 168854 58000 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 58000 168854
rect -4886 168586 58000 168618
rect 472044 169174 588810 169206
rect 472044 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 472044 168854 588810 168938
rect 472044 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 472044 168586 588810 168618
rect -2966 165454 58000 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 58000 165454
rect -2966 165134 58000 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 58000 165134
rect -2966 164866 58000 164898
rect 472044 165454 586890 165486
rect 472044 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 472044 165134 586890 165218
rect 472044 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 472044 164866 586890 164898
rect -8726 158614 58000 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 58000 158614
rect -8726 158294 58000 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 58000 158294
rect -8726 158026 58000 158058
rect 472044 158614 592650 158646
rect 472044 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect 472044 158294 592650 158378
rect 472044 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect 472044 158026 592650 158058
rect -6806 154894 58000 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 58000 154894
rect -6806 154574 58000 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 58000 154574
rect -6806 154306 58000 154338
rect 472044 154894 590730 154926
rect 472044 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect 472044 154574 590730 154658
rect 472044 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect 472044 154306 590730 154338
rect -4886 151174 58000 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 58000 151174
rect -4886 150854 58000 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 58000 150854
rect -4886 150586 58000 150618
rect 472044 151174 588810 151206
rect 472044 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect 472044 150854 588810 150938
rect 472044 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect 472044 150586 588810 150618
rect -2966 147454 58000 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 58000 147454
rect -2966 147134 58000 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 58000 147134
rect -2966 146866 58000 146898
rect 472044 147454 586890 147486
rect 472044 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect 472044 147134 586890 147218
rect 472044 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect 472044 146866 586890 146898
rect -8726 140614 58000 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 58000 140614
rect -8726 140294 58000 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 58000 140294
rect -8726 140026 58000 140058
rect 472044 140614 592650 140646
rect 472044 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 472044 140294 592650 140378
rect 472044 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 472044 140026 592650 140058
rect -6806 136894 58000 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 58000 136894
rect -6806 136574 58000 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 58000 136574
rect -6806 136306 58000 136338
rect 472044 136894 590730 136926
rect 472044 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 472044 136574 590730 136658
rect 472044 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 472044 136306 590730 136338
rect -4886 133174 58000 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 58000 133174
rect -4886 132854 58000 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 58000 132854
rect -4886 132586 58000 132618
rect 472044 133174 588810 133206
rect 472044 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 472044 132854 588810 132938
rect 472044 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 472044 132586 588810 132618
rect -2966 129454 58000 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 58000 129454
rect -2966 129134 58000 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 58000 129134
rect -2966 128866 58000 128898
rect 472044 129454 586890 129486
rect 472044 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 472044 129134 586890 129218
rect 472044 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 472044 128866 586890 128898
rect -8726 122614 58000 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 58000 122614
rect -8726 122294 58000 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 58000 122294
rect -8726 122026 58000 122058
rect 472044 122614 592650 122646
rect 472044 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect 472044 122294 592650 122378
rect 472044 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect 472044 122026 592650 122058
rect -6806 118894 58000 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 58000 118894
rect -6806 118574 58000 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 58000 118574
rect -6806 118306 58000 118338
rect 472044 118894 590730 118926
rect 472044 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect 472044 118574 590730 118658
rect 472044 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect 472044 118306 590730 118338
rect -4886 115174 58000 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 58000 115174
rect -4886 114854 58000 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 58000 114854
rect -4886 114586 58000 114618
rect 472044 115174 588810 115206
rect 472044 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect 472044 114854 588810 114938
rect 472044 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect 472044 114586 588810 114618
rect -2966 111454 58000 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 58000 111454
rect -2966 111134 58000 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 58000 111134
rect -2966 110866 58000 110898
rect 472044 111454 586890 111486
rect 472044 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect 472044 111134 586890 111218
rect 472044 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect 472044 110866 586890 110898
rect -8726 104614 58000 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 58000 104614
rect -8726 104294 58000 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 58000 104294
rect -8726 104026 58000 104058
rect 472044 104614 592650 104646
rect 472044 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 472044 104294 592650 104378
rect 472044 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 472044 104026 592650 104058
rect -6806 100894 58000 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 58000 100894
rect -6806 100574 58000 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 58000 100574
rect -6806 100306 58000 100338
rect 472044 100894 590730 100926
rect 472044 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 472044 100574 590730 100658
rect 472044 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 472044 100306 590730 100338
rect -4886 97174 58000 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 58000 97174
rect -4886 96854 58000 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 58000 96854
rect -4886 96586 58000 96618
rect 472044 97174 588810 97206
rect 472044 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 472044 96854 588810 96938
rect 472044 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 472044 96586 588810 96618
rect -2966 93454 58000 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 58000 93454
rect -2966 93134 58000 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 58000 93134
rect -2966 92866 58000 92898
rect 472044 93454 586890 93486
rect 472044 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 472044 93134 586890 93218
rect 472044 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 472044 92866 586890 92898
rect -8726 86614 58000 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 58000 86614
rect -8726 86294 58000 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 58000 86294
rect -8726 86026 58000 86058
rect 472044 86614 592650 86646
rect 472044 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect 472044 86294 592650 86378
rect 472044 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect 472044 86026 592650 86058
rect -6806 82894 58000 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 58000 82894
rect -6806 82574 58000 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 58000 82574
rect -6806 82306 58000 82338
rect 472044 82894 590730 82926
rect 472044 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect 472044 82574 590730 82658
rect 472044 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect 472044 82306 590730 82338
rect -4886 79174 58000 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 58000 79174
rect -4886 78854 58000 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 58000 78854
rect -4886 78586 58000 78618
rect 472044 79174 588810 79206
rect 472044 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect 472044 78854 588810 78938
rect 472044 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect 472044 78586 588810 78618
rect -2966 75454 58000 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 58000 75454
rect -2966 75134 58000 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 58000 75134
rect -2966 74866 58000 74898
rect 472044 75454 586890 75486
rect 472044 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect 472044 75134 586890 75218
rect 472044 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect 472044 74866 586890 74898
rect -8726 68614 58000 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 58000 68614
rect -8726 68294 58000 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 58000 68294
rect -8726 68026 58000 68058
rect 472044 68614 592650 68646
rect 472044 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 472044 68294 592650 68378
rect 472044 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 472044 68026 592650 68058
rect -6806 64894 58000 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 58000 64894
rect -6806 64574 58000 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 58000 64574
rect -6806 64306 58000 64338
rect 472044 64894 590730 64926
rect 472044 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 472044 64574 590730 64658
rect 472044 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 472044 64306 590730 64338
rect -4886 61174 58000 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 58000 61174
rect -4886 60854 58000 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 58000 60854
rect -4886 60586 58000 60618
rect 472044 61174 588810 61206
rect 472044 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 472044 60854 588810 60938
rect 472044 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 472044 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use azadi_soc_top_caravel  mprj
timestamp 0
transform 1 0 60000 0 1 60000
box 0 0 410044 389980
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 58000 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s 472044 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 58000 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s 472044 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 58000 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s 472044 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 58000 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s 472044 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 58000 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s 472044 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 58000 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s 472044 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 58000 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s 472044 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 58000 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s 472044 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 58000 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s 472044 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 58000 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s 472044 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 58000 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s 472044 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 451980 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 451980 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 451980 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 451980 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 451980 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 451980 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 451980 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 451980 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 451980 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 451980 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 451980 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 451980 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 58000 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s 472044 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 58000 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s 472044 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 58000 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s 472044 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 58000 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s 472044 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 58000 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s 472044 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 58000 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s 472044 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 58000 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s 472044 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 58000 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s 472044 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 58000 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s 472044 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 58000 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s 472044 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 58000 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s 472044 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 451980 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 451980 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 451980 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 451980 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 451980 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 451980 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 451980 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 451980 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 451980 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 451980 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 451980 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 58000 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s 472044 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 58000 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s 472044 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 58000 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s 472044 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 58000 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s 472044 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 58000 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s 472044 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 58000 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s 472044 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 58000 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s 472044 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 58000 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s 472044 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 58000 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s 472044 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 58000 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s 472044 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 58000 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s 472044 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 451980 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 451980 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 451980 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 451980 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 451980 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 451980 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 451980 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 451980 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 451980 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 451980 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 451980 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 58000 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s 472044 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 58000 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s 472044 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 58000 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s 472044 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 58000 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s 472044 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 58000 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s 472044 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 58000 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s 472044 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 58000 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s 472044 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 58000 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s 472044 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 58000 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s 472044 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 58000 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s 472044 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 58000 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s 472044 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 451980 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 451980 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 451980 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 451980 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 451980 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 451980 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 451980 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 451980 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 451980 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 451980 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 451980 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 58000 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 472044 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 58000 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 472044 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 58000 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 472044 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 58000 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 472044 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 58000 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 472044 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 58000 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 472044 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 58000 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 472044 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 58000 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 472044 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 58000 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 472044 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 58000 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 472044 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 58000 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 472044 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 451980 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 451980 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 451980 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 451980 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 451980 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 451980 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 451980 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 451980 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 451980 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 451980 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 451980 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 451980 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 58000 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 472044 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 58000 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 472044 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 58000 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 472044 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 58000 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 472044 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 58000 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 472044 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 58000 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 472044 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 58000 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 472044 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 58000 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 472044 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 58000 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 472044 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 58000 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 472044 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 58000 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 472044 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 451980 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 451980 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 451980 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 451980 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 451980 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 451980 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 451980 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 451980 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 451980 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 451980 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 451980 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 451980 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 58000 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 472044 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 58000 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 472044 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 58000 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 472044 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 58000 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 472044 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 58000 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 472044 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 58000 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 472044 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 58000 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 472044 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 58000 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 472044 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 58000 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 472044 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 58000 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 472044 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 451980 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 451980 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 451980 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 451980 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 451980 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 451980 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 451980 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 451980 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 451980 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 451980 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 451980 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 58000 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 472044 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 58000 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 472044 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 58000 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 472044 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 58000 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 472044 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 58000 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 472044 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 58000 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 472044 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 58000 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 472044 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 58000 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 472044 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 58000 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 472044 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 58000 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 472044 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 58000 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 472044 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 451980 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 451980 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 451980 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 451980 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 451980 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 451980 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 451980 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 451980 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 451980 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 451980 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 451980 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 451980 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
