magic
tech sky130A
magscale 1 2
timestamp 1654247864
<< metal1 >>
rect 1394 444388 1400 444440
rect 1452 444428 1458 444440
rect 57606 444428 57612 444440
rect 1452 444400 57612 444428
rect 1452 444388 1458 444400
rect 57606 444388 57612 444400
rect 57664 444388 57670 444440
rect 105630 59820 105636 59832
rect 103486 59792 105636 59820
rect 63310 59712 63316 59764
rect 63368 59752 63374 59764
rect 64322 59752 64328 59764
rect 63368 59724 64328 59752
rect 63368 59712 63374 59724
rect 64322 59712 64328 59724
rect 64380 59712 64386 59764
rect 72786 59712 72792 59764
rect 72844 59752 72850 59764
rect 75086 59752 75092 59764
rect 72844 59724 75092 59752
rect 72844 59712 72850 59724
rect 75086 59712 75092 59724
rect 75144 59712 75150 59764
rect 78582 59712 78588 59764
rect 78640 59752 78646 59764
rect 79962 59752 79968 59764
rect 78640 59724 79968 59752
rect 78640 59712 78646 59724
rect 79962 59712 79968 59724
rect 80020 59712 80026 59764
rect 92382 59712 92388 59764
rect 92440 59752 92446 59764
rect 93854 59752 93860 59764
rect 92440 59724 93860 59752
rect 92440 59712 92446 59724
rect 93854 59712 93860 59724
rect 93912 59712 93918 59764
rect 98638 59712 98644 59764
rect 98696 59752 98702 59764
rect 101398 59752 101404 59764
rect 98696 59724 101404 59752
rect 98696 59712 98702 59724
rect 101398 59712 101404 59724
rect 101456 59712 101462 59764
rect 102778 59712 102784 59764
rect 102836 59752 102842 59764
rect 103486 59752 103514 59792
rect 105630 59780 105636 59792
rect 105688 59780 105694 59832
rect 110322 59780 110328 59832
rect 110380 59820 110386 59832
rect 111334 59820 111340 59832
rect 110380 59792 111340 59820
rect 110380 59780 110386 59792
rect 111334 59780 111340 59792
rect 111392 59780 111398 59832
rect 229462 59780 229468 59832
rect 229520 59820 229526 59832
rect 230658 59820 230664 59832
rect 229520 59792 230664 59820
rect 229520 59780 229526 59792
rect 230658 59780 230664 59792
rect 230716 59780 230722 59832
rect 240502 59820 240508 59832
rect 238726 59792 240508 59820
rect 102836 59724 103514 59752
rect 102836 59712 102842 59724
rect 105538 59712 105544 59764
rect 105596 59752 105602 59764
rect 108022 59752 108028 59764
rect 105596 59724 108028 59752
rect 105596 59712 105602 59724
rect 108022 59712 108028 59724
rect 108080 59712 108086 59764
rect 111058 59712 111064 59764
rect 111116 59752 111122 59764
rect 113726 59752 113732 59764
rect 111116 59724 113732 59752
rect 111116 59712 111122 59724
rect 113726 59712 113732 59724
rect 113784 59712 113790 59764
rect 114002 59712 114008 59764
rect 114060 59752 114066 59764
rect 116210 59752 116216 59764
rect 114060 59724 116216 59752
rect 114060 59712 114066 59724
rect 116210 59712 116216 59724
rect 116268 59712 116274 59764
rect 119522 59712 119528 59764
rect 119580 59752 119586 59764
rect 122006 59752 122012 59764
rect 119580 59724 122012 59752
rect 119580 59712 119586 59724
rect 122006 59712 122012 59724
rect 122064 59712 122070 59764
rect 124858 59712 124864 59764
rect 124916 59752 124922 59764
rect 126422 59752 126428 59764
rect 124916 59724 126428 59752
rect 124916 59712 124922 59724
rect 126422 59712 126428 59724
rect 126480 59712 126486 59764
rect 127618 59712 127624 59764
rect 127676 59752 127682 59764
rect 130194 59752 130200 59764
rect 127676 59724 130200 59752
rect 127676 59712 127682 59724
rect 130194 59712 130200 59724
rect 130252 59712 130258 59764
rect 140682 59712 140688 59764
rect 140740 59752 140746 59764
rect 141694 59752 141700 59764
rect 140740 59724 141700 59752
rect 140740 59712 140746 59724
rect 141694 59712 141700 59724
rect 141752 59712 141758 59764
rect 150066 59712 150072 59764
rect 150124 59752 150130 59764
rect 151906 59752 151912 59764
rect 150124 59724 151912 59752
rect 150124 59712 150130 59724
rect 151906 59712 151912 59724
rect 151964 59712 151970 59764
rect 157150 59712 157156 59764
rect 157208 59752 157214 59764
rect 158162 59752 158168 59764
rect 157208 59724 158168 59752
rect 157208 59712 157214 59724
rect 158162 59712 158168 59724
rect 158220 59712 158226 59764
rect 172422 59712 172428 59764
rect 172480 59752 172486 59764
rect 173342 59752 173348 59764
rect 172480 59724 173348 59752
rect 172480 59712 172486 59724
rect 173342 59712 173348 59724
rect 173400 59712 173406 59764
rect 182082 59712 182088 59764
rect 182140 59752 182146 59764
rect 183738 59752 183744 59764
rect 182140 59724 183744 59752
rect 182140 59712 182146 59724
rect 183738 59712 183744 59724
rect 183796 59712 183802 59764
rect 192846 59712 192852 59764
rect 192904 59752 192910 59764
rect 194410 59752 194416 59764
rect 192904 59724 194416 59752
rect 192904 59712 192910 59724
rect 194410 59712 194416 59724
rect 194468 59712 194474 59764
rect 199838 59712 199844 59764
rect 199896 59752 199902 59764
rect 200206 59752 200212 59764
rect 199896 59724 200212 59752
rect 199896 59712 199902 59724
rect 200206 59712 200212 59724
rect 200264 59712 200270 59764
rect 201310 59712 201316 59764
rect 201368 59752 201374 59764
rect 202782 59752 202788 59764
rect 201368 59724 202788 59752
rect 201368 59712 201374 59724
rect 202782 59712 202788 59724
rect 202840 59712 202846 59764
rect 208210 59712 208216 59764
rect 208268 59752 208274 59764
rect 209406 59752 209412 59764
rect 208268 59724 209412 59752
rect 208268 59712 208274 59724
rect 209406 59712 209412 59724
rect 209464 59712 209470 59764
rect 213546 59712 213552 59764
rect 213604 59752 213610 59764
rect 215846 59752 215852 59764
rect 213604 59724 215852 59752
rect 213604 59712 213610 59724
rect 215846 59712 215852 59724
rect 215904 59712 215910 59764
rect 232498 59712 232504 59764
rect 232556 59752 232562 59764
rect 234798 59752 234804 59764
rect 232556 59724 234804 59752
rect 232556 59712 232562 59724
rect 234798 59712 234804 59724
rect 234856 59712 234862 59764
rect 238018 59712 238024 59764
rect 238076 59752 238082 59764
rect 238726 59752 238754 59792
rect 240502 59780 240508 59792
rect 240560 59780 240566 59832
rect 296990 59780 296996 59832
rect 297048 59820 297054 59832
rect 298922 59820 298928 59832
rect 297048 59792 298928 59820
rect 297048 59780 297054 59792
rect 298922 59780 298928 59792
rect 298980 59780 298986 59832
rect 380066 59780 380072 59832
rect 380124 59820 380130 59832
rect 382918 59820 382924 59832
rect 380124 59792 382924 59820
rect 380124 59780 380130 59792
rect 382918 59780 382924 59792
rect 382976 59780 382982 59832
rect 238076 59724 238754 59752
rect 238076 59712 238082 59724
rect 239398 59712 239404 59764
rect 239456 59752 239462 59764
rect 242158 59752 242164 59764
rect 239456 59724 242164 59752
rect 239456 59712 239462 59724
rect 242158 59712 242164 59724
rect 242216 59712 242222 59764
rect 244182 59712 244188 59764
rect 244240 59752 244246 59764
rect 245470 59752 245476 59764
rect 244240 59724 245476 59752
rect 244240 59712 244246 59724
rect 245470 59712 245476 59724
rect 245528 59712 245534 59764
rect 249058 59712 249064 59764
rect 249116 59752 249122 59764
rect 251266 59752 251272 59764
rect 249116 59724 251272 59752
rect 249116 59712 249122 59724
rect 251266 59712 251272 59724
rect 251324 59712 251330 59764
rect 267458 59712 267464 59764
rect 267516 59752 267522 59764
rect 269942 59752 269948 59764
rect 267516 59724 269948 59752
rect 267516 59712 267522 59724
rect 269942 59712 269948 59724
rect 270000 59712 270006 59764
rect 270678 59712 270684 59764
rect 270736 59752 270742 59764
rect 271874 59752 271880 59764
rect 270736 59724 271880 59752
rect 270736 59712 270742 59724
rect 271874 59712 271880 59724
rect 271932 59712 271938 59764
rect 277210 59712 277216 59764
rect 277268 59752 277274 59764
rect 277854 59752 277860 59764
rect 277268 59724 277860 59752
rect 277268 59712 277274 59724
rect 277854 59712 277860 59724
rect 277912 59712 277918 59764
rect 283006 59712 283012 59764
rect 283064 59752 283070 59764
rect 284294 59752 284300 59764
rect 283064 59724 284300 59752
rect 283064 59712 283070 59724
rect 284294 59712 284300 59724
rect 284352 59712 284358 59764
rect 287882 59712 287888 59764
rect 287940 59752 287946 59764
rect 290642 59752 290648 59764
rect 287940 59724 290648 59752
rect 287940 59712 287946 59724
rect 290642 59712 290648 59724
rect 290700 59712 290706 59764
rect 293678 59712 293684 59764
rect 293736 59752 293742 59764
rect 295978 59752 295984 59764
rect 293736 59724 295984 59752
rect 293736 59712 293742 59724
rect 295978 59712 295984 59724
rect 296036 59712 296042 59764
rect 296530 59712 296536 59764
rect 296588 59752 296594 59764
rect 298738 59752 298744 59764
rect 296588 59724 298744 59752
rect 296588 59712 296594 59724
rect 298738 59712 298744 59724
rect 298796 59712 298802 59764
rect 301958 59712 301964 59764
rect 302016 59752 302022 59764
rect 304258 59752 304264 59764
rect 302016 59724 304264 59752
rect 302016 59712 302022 59724
rect 304258 59712 304264 59724
rect 304316 59712 304322 59764
rect 314286 59712 314292 59764
rect 314344 59752 314350 59764
rect 316678 59752 316684 59764
rect 314344 59724 316684 59752
rect 314344 59712 314350 59724
rect 316678 59712 316684 59724
rect 316736 59712 316742 59764
rect 320818 59712 320824 59764
rect 320876 59752 320882 59764
rect 323118 59752 323124 59764
rect 320876 59724 323124 59752
rect 320876 59712 320882 59724
rect 323118 59712 323124 59724
rect 323176 59712 323182 59764
rect 324958 59712 324964 59764
rect 325016 59752 325022 59764
rect 327350 59752 327356 59764
rect 325016 59724 327356 59752
rect 325016 59712 325022 59724
rect 327350 59712 327356 59724
rect 327408 59712 327414 59764
rect 334894 59712 334900 59764
rect 334952 59752 334958 59764
rect 336918 59752 336924 59764
rect 334952 59724 336924 59752
rect 334952 59712 334958 59724
rect 336918 59712 336924 59724
rect 336976 59712 336982 59764
rect 339034 59712 339040 59764
rect 339092 59752 339098 59764
rect 341150 59752 341156 59764
rect 339092 59724 341156 59752
rect 339092 59712 339098 59724
rect 341150 59712 341156 59724
rect 341208 59712 341214 59764
rect 341518 59712 341524 59764
rect 341576 59752 341582 59764
rect 342530 59752 342536 59764
rect 341576 59724 342536 59752
rect 341576 59712 341582 59724
rect 342530 59712 342536 59724
rect 342588 59712 342594 59764
rect 343082 59712 343088 59764
rect 343140 59752 343146 59764
rect 345106 59752 345112 59764
rect 343140 59724 345112 59752
rect 343140 59712 343146 59724
rect 345106 59712 345112 59724
rect 345164 59712 345170 59764
rect 359550 59712 359556 59764
rect 359608 59752 359614 59764
rect 361758 59752 361764 59764
rect 359608 59724 361764 59752
rect 359608 59712 359614 59724
rect 361758 59712 361764 59724
rect 361816 59712 361822 59764
rect 363690 59712 363696 59764
rect 363748 59752 363754 59764
rect 366358 59752 366364 59764
rect 363748 59724 366364 59752
rect 363748 59712 363754 59724
rect 366358 59712 366364 59724
rect 366416 59712 366422 59764
rect 367002 59712 367008 59764
rect 367060 59752 367066 59764
rect 369118 59752 369124 59764
rect 367060 59724 369124 59752
rect 367060 59712 367066 59724
rect 369118 59712 369124 59724
rect 369176 59712 369182 59764
rect 369394 59712 369400 59764
rect 369452 59752 369458 59764
rect 369452 59724 369854 59752
rect 369452 59712 369458 59724
rect 24854 59644 24860 59696
rect 24912 59684 24918 59696
rect 61010 59684 61016 59696
rect 24912 59656 61016 59684
rect 24912 59644 24918 59656
rect 61010 59644 61016 59656
rect 61068 59644 61074 59696
rect 95878 59644 95884 59696
rect 95936 59684 95942 59696
rect 97350 59684 97356 59696
rect 95936 59656 97356 59684
rect 95936 59644 95942 59656
rect 97350 59644 97356 59656
rect 97408 59644 97414 59696
rect 236638 59644 236644 59696
rect 236696 59684 236702 59696
rect 238846 59684 238852 59696
rect 236696 59656 238852 59684
rect 236696 59644 236702 59656
rect 238846 59644 238852 59656
rect 238904 59644 238910 59696
rect 269850 59644 269856 59696
rect 269908 59684 269914 59696
rect 272518 59684 272524 59696
rect 269908 59656 272524 59684
rect 269908 59644 269914 59656
rect 272518 59644 272524 59656
rect 272576 59644 272582 59696
rect 286318 59644 286324 59696
rect 286376 59684 286382 59696
rect 288434 59684 288440 59696
rect 286376 59656 288440 59684
rect 286376 59644 286382 59656
rect 288434 59644 288440 59656
rect 288492 59644 288498 59696
rect 300302 59644 300308 59696
rect 300360 59684 300366 59696
rect 302878 59684 302884 59696
rect 300360 59656 302884 59684
rect 300360 59644 300366 59656
rect 302878 59644 302884 59656
rect 302936 59644 302942 59696
rect 312538 59644 312544 59696
rect 312596 59684 312602 59696
rect 313918 59684 313924 59696
rect 312596 59656 313924 59684
rect 312596 59644 312602 59656
rect 313918 59644 313924 59656
rect 313976 59644 313982 59696
rect 365162 59644 365168 59696
rect 365220 59684 365226 59696
rect 366542 59684 366548 59696
rect 365220 59656 366548 59684
rect 365220 59644 365226 59656
rect 366542 59644 366548 59656
rect 366600 59644 366606 59696
rect 369826 59684 369854 59724
rect 371050 59712 371056 59764
rect 371108 59752 371114 59764
rect 372614 59752 372620 59764
rect 371108 59724 372620 59752
rect 371108 59712 371114 59724
rect 372614 59712 372620 59724
rect 372672 59712 372678 59764
rect 376018 59712 376024 59764
rect 376076 59752 376082 59764
rect 378962 59752 378968 59764
rect 376076 59724 378968 59752
rect 376076 59712 376082 59724
rect 378962 59712 378968 59724
rect 379020 59712 379026 59764
rect 379422 59712 379428 59764
rect 379480 59752 379486 59764
rect 380158 59752 380164 59764
rect 379480 59724 380164 59752
rect 379480 59712 379486 59724
rect 380158 59712 380164 59724
rect 380216 59712 380222 59764
rect 380986 59712 380992 59764
rect 381044 59752 381050 59764
rect 382274 59752 382280 59764
rect 381044 59724 382280 59752
rect 381044 59712 381050 59724
rect 382274 59712 382280 59724
rect 382332 59712 382338 59764
rect 387518 59712 387524 59764
rect 387576 59752 387582 59764
rect 389818 59752 389824 59764
rect 387576 59724 389824 59752
rect 387576 59712 387582 59724
rect 389818 59712 389824 59724
rect 389876 59712 389882 59764
rect 391658 59712 391664 59764
rect 391716 59752 391722 59764
rect 393958 59752 393964 59764
rect 391716 59724 393964 59752
rect 391716 59712 391722 59724
rect 393958 59712 393964 59724
rect 394016 59712 394022 59764
rect 397454 59712 397460 59764
rect 397512 59752 397518 59764
rect 399478 59752 399484 59764
rect 397512 59724 399484 59752
rect 397512 59712 397518 59724
rect 399478 59712 399484 59724
rect 399536 59712 399542 59764
rect 402330 59712 402336 59764
rect 402388 59752 402394 59764
rect 404446 59752 404452 59764
rect 402388 59724 404452 59752
rect 402388 59712 402394 59724
rect 404446 59712 404452 59724
rect 404504 59712 404510 59764
rect 406470 59712 406476 59764
rect 406528 59752 406534 59764
rect 408494 59752 408500 59764
rect 406528 59724 408500 59752
rect 406528 59712 406534 59724
rect 408494 59712 408500 59724
rect 408552 59712 408558 59764
rect 410610 59712 410616 59764
rect 410668 59752 410674 59764
rect 412818 59752 412824 59764
rect 410668 59724 412824 59752
rect 410668 59712 410674 59724
rect 412818 59712 412824 59724
rect 412876 59712 412882 59764
rect 425514 59712 425520 59764
rect 425572 59752 425578 59764
rect 426526 59752 426532 59764
rect 425572 59724 426532 59752
rect 425572 59712 425578 59724
rect 426526 59712 426532 59724
rect 426584 59712 426590 59764
rect 427078 59712 427084 59764
rect 427136 59752 427142 59764
rect 429562 59752 429568 59764
rect 427136 59724 429568 59752
rect 427136 59712 427142 59724
rect 429562 59712 429568 59724
rect 429620 59712 429626 59764
rect 431218 59712 431224 59764
rect 431276 59752 431282 59764
rect 433610 59752 433616 59764
rect 431276 59724 433616 59752
rect 431276 59712 431282 59724
rect 433610 59712 433616 59724
rect 433668 59712 433674 59764
rect 436922 59712 436928 59764
rect 436980 59752 436986 59764
rect 439222 59752 439228 59764
rect 436980 59724 439228 59752
rect 436980 59712 436986 59724
rect 439222 59712 439228 59724
rect 439280 59712 439286 59764
rect 441890 59712 441896 59764
rect 441948 59752 441954 59764
rect 443178 59752 443184 59764
rect 441948 59724 443184 59752
rect 441948 59712 441954 59724
rect 443178 59712 443184 59724
rect 443236 59712 443242 59764
rect 446858 59712 446864 59764
rect 446916 59752 446922 59764
rect 448790 59752 448796 59764
rect 446916 59724 448796 59752
rect 446916 59712 446922 59724
rect 448790 59712 448796 59724
rect 448848 59712 448854 59764
rect 457530 59712 457536 59764
rect 457588 59752 457594 59764
rect 459922 59752 459928 59764
rect 457588 59724 459928 59752
rect 457588 59712 457594 59724
rect 459922 59712 459928 59724
rect 459980 59712 459986 59764
rect 464154 59712 464160 59764
rect 464212 59752 464218 59764
rect 465350 59752 465356 59764
rect 464212 59724 465356 59752
rect 464212 59712 464218 59724
rect 465350 59712 465356 59724
rect 465408 59712 465414 59764
rect 371326 59684 371332 59696
rect 369826 59656 371332 59684
rect 371326 59644 371332 59656
rect 371384 59644 371390 59696
rect 390002 59644 390008 59696
rect 390060 59684 390066 59696
rect 392578 59684 392584 59696
rect 390060 59656 392584 59684
rect 390060 59644 390066 59656
rect 392578 59644 392584 59656
rect 392636 59644 392642 59696
rect 19334 59576 19340 59628
rect 19392 59616 19398 59628
rect 60458 59616 60464 59628
rect 19392 59588 60464 59616
rect 19392 59576 19398 59588
rect 60458 59576 60464 59588
rect 60516 59576 60522 59628
rect 67450 59576 67456 59628
rect 67508 59616 67514 59628
rect 69290 59616 69296 59628
rect 67508 59588 69296 59616
rect 67508 59576 67514 59588
rect 69290 59576 69296 59588
rect 69348 59576 69354 59628
rect 75362 59576 75368 59628
rect 75420 59616 75426 59628
rect 77478 59616 77484 59628
rect 75420 59588 77484 59616
rect 75420 59576 75426 59588
rect 77478 59576 77484 59588
rect 77536 59576 77542 59628
rect 87598 59576 87604 59628
rect 87656 59616 87662 59628
rect 89070 59616 89076 59628
rect 87656 59588 89076 59616
rect 87656 59576 87662 59588
rect 89070 59576 89076 59588
rect 89128 59576 89134 59628
rect 118142 59576 118148 59628
rect 118200 59616 118206 59628
rect 120350 59616 120356 59628
rect 118200 59588 120356 59616
rect 118200 59576 118206 59588
rect 120350 59576 120356 59588
rect 120408 59576 120414 59628
rect 130562 59576 130568 59628
rect 130620 59616 130626 59628
rect 131942 59616 131948 59628
rect 130620 59588 131948 59616
rect 130620 59576 130626 59588
rect 131942 59576 131948 59588
rect 132000 59576 132006 59628
rect 140038 59576 140044 59628
rect 140096 59616 140102 59628
rect 141694 59616 141700 59628
rect 140096 59588 141700 59616
rect 140096 59576 140102 59588
rect 141694 59576 141700 59588
rect 141752 59576 141758 59628
rect 150250 59576 150256 59628
rect 150308 59616 150314 59628
rect 151630 59616 151636 59628
rect 150308 59588 151636 59616
rect 150308 59576 150314 59588
rect 151630 59576 151636 59588
rect 151688 59576 151694 59628
rect 165430 59576 165436 59628
rect 165488 59616 165494 59628
rect 166442 59616 166448 59628
rect 165488 59588 166448 59616
rect 165488 59576 165494 59588
rect 166442 59576 166448 59588
rect 166500 59576 166506 59628
rect 174906 59576 174912 59628
rect 174964 59616 174970 59628
rect 177114 59616 177120 59628
rect 174964 59588 177120 59616
rect 174964 59576 174970 59588
rect 177114 59576 177120 59588
rect 177172 59576 177178 59628
rect 217686 59576 217692 59628
rect 217744 59616 217750 59628
rect 219158 59616 219164 59628
rect 217744 59588 219164 59616
rect 217744 59576 217750 59588
rect 219158 59576 219164 59588
rect 219216 59576 219222 59628
rect 227622 59576 227628 59628
rect 227680 59616 227686 59628
rect 229002 59616 229008 59628
rect 227680 59588 229008 59616
rect 227680 59576 227686 59588
rect 229002 59576 229008 59588
rect 229060 59576 229066 59628
rect 246482 59576 246488 59628
rect 246540 59616 246546 59628
rect 248874 59616 248880 59628
rect 246540 59588 248880 59616
rect 246540 59576 246546 59588
rect 248874 59576 248880 59588
rect 248932 59576 248938 59628
rect 256326 59576 256332 59628
rect 256384 59616 256390 59628
rect 257798 59616 257804 59628
rect 256384 59588 257804 59616
rect 256384 59576 256390 59588
rect 257798 59576 257804 59588
rect 257856 59576 257862 59628
rect 259086 59576 259092 59628
rect 259144 59616 259150 59628
rect 261110 59616 261116 59628
rect 259144 59588 261116 59616
rect 259144 59576 259150 59588
rect 261110 59576 261116 59588
rect 261168 59576 261174 59628
rect 280338 59576 280344 59628
rect 280396 59616 280402 59628
rect 282178 59616 282184 59628
rect 280396 59588 282184 59616
rect 280396 59576 280402 59588
rect 282178 59576 282184 59588
rect 282236 59576 282242 59628
rect 306006 59576 306012 59628
rect 306064 59616 306070 59628
rect 307202 59616 307208 59628
rect 306064 59588 307208 59616
rect 306064 59576 306070 59588
rect 307202 59576 307208 59588
rect 307260 59576 307266 59628
rect 310146 59576 310152 59628
rect 310204 59616 310210 59628
rect 312722 59616 312728 59628
rect 310204 59588 312728 59616
rect 310204 59576 310210 59588
rect 312722 59576 312728 59588
rect 312780 59576 312786 59628
rect 376018 59576 376024 59628
rect 376076 59616 376082 59628
rect 377398 59616 377404 59628
rect 376076 59588 377404 59616
rect 376076 59576 376082 59588
rect 377398 59576 377404 59588
rect 377456 59576 377462 59628
rect 393314 59576 393320 59628
rect 393372 59616 393378 59628
rect 395338 59616 395344 59628
rect 393372 59588 395344 59616
rect 393372 59576 393378 59588
rect 395338 59576 395344 59588
rect 395396 59576 395402 59628
rect 413094 59576 413100 59628
rect 413152 59616 413158 59628
rect 414106 59616 414112 59628
rect 413152 59588 414112 59616
rect 413152 59576 413158 59588
rect 414106 59576 414112 59588
rect 414164 59576 414170 59628
rect 416406 59576 416412 59628
rect 416464 59616 416470 59628
rect 418246 59616 418252 59628
rect 416464 59588 418252 59616
rect 416464 59576 416470 59588
rect 418246 59576 418252 59588
rect 418304 59576 418310 59628
rect 449250 59576 449256 59628
rect 449308 59616 449314 59628
rect 449894 59616 449900 59628
rect 449308 59588 449900 59616
rect 449308 59576 449314 59588
rect 449894 59576 449900 59588
rect 449952 59576 449958 59628
rect 453390 59576 453396 59628
rect 453448 59616 453454 59628
rect 455690 59616 455696 59628
rect 453448 59588 455696 59616
rect 453448 59576 453454 59588
rect 455690 59576 455696 59588
rect 455748 59576 455754 59628
rect 15194 59508 15200 59560
rect 15252 59548 15258 59560
rect 59354 59548 59360 59560
rect 15252 59520 59360 59548
rect 15252 59508 15258 59520
rect 59354 59508 59360 59520
rect 59412 59508 59418 59560
rect 247862 59508 247868 59560
rect 247920 59548 247926 59560
rect 250530 59548 250536 59560
rect 247920 59520 250536 59548
rect 247920 59508 247926 59520
rect 250530 59508 250536 59520
rect 250588 59508 250594 59560
rect 5534 59440 5540 59492
rect 5592 59480 5598 59492
rect 57606 59480 57612 59492
rect 5592 59452 57612 59480
rect 5592 59440 5598 59452
rect 57606 59440 57612 59452
rect 57664 59440 57670 59492
rect 85022 59440 85028 59492
rect 85080 59480 85086 59492
rect 87414 59480 87420 59492
rect 85080 59452 87420 59480
rect 85080 59440 85086 59452
rect 87414 59440 87420 59452
rect 87472 59440 87478 59492
rect 89530 59440 89536 59492
rect 89588 59480 89594 59492
rect 91554 59480 91560 59492
rect 89588 59452 91560 59480
rect 89588 59440 89594 59452
rect 91554 59440 91560 59452
rect 91612 59440 91618 59492
rect 166626 59440 166632 59492
rect 166684 59480 166690 59492
rect 168926 59480 168932 59492
rect 166684 59452 168932 59480
rect 166684 59440 166690 59452
rect 168926 59440 168932 59452
rect 168984 59440 168990 59492
rect 169386 59440 169392 59492
rect 169444 59480 169450 59492
rect 171410 59480 171416 59492
rect 169444 59452 171416 59480
rect 169444 59440 169450 59452
rect 171410 59440 171416 59452
rect 171468 59440 171474 59492
rect 179322 59440 179328 59492
rect 179380 59480 179386 59492
rect 180426 59480 180432 59492
rect 179380 59452 180432 59480
rect 179380 59440 179386 59452
rect 180426 59440 180432 59452
rect 180484 59440 180490 59492
rect 188890 59440 188896 59492
rect 188948 59480 188954 59492
rect 190270 59480 190276 59492
rect 188948 59452 190276 59480
rect 188948 59440 188954 59452
rect 190270 59440 190276 59452
rect 190328 59440 190334 59492
rect 190546 59480 190552 59492
rect 190426 59452 190552 59480
rect 4154 59372 4160 59424
rect 4212 59412 4218 59424
rect 57974 59412 57980 59424
rect 4212 59384 57980 59412
rect 4212 59372 4218 59384
rect 57974 59372 57980 59384
rect 58032 59372 58038 59424
rect 138106 59372 138112 59424
rect 138164 59412 138170 59424
rect 139302 59412 139308 59424
rect 138164 59384 139308 59412
rect 138164 59372 138170 59384
rect 139302 59372 139308 59384
rect 139360 59372 139366 59424
rect 188706 59372 188712 59424
rect 188764 59412 188770 59424
rect 190426 59412 190454 59452
rect 190546 59440 190552 59452
rect 190604 59440 190610 59492
rect 205266 59440 205272 59492
rect 205324 59480 205330 59492
rect 207566 59480 207572 59492
rect 205324 59452 207572 59480
rect 205324 59440 205330 59452
rect 207566 59440 207572 59452
rect 207624 59440 207630 59492
rect 246298 59440 246304 59492
rect 246356 59480 246362 59492
rect 247954 59480 247960 59492
rect 246356 59452 247960 59480
rect 246356 59440 246362 59452
rect 247954 59440 247960 59452
rect 248012 59440 248018 59492
rect 272242 59440 272248 59492
rect 272300 59480 272306 59492
rect 273254 59480 273260 59492
rect 272300 59452 273260 59480
rect 272300 59440 272306 59452
rect 273254 59440 273260 59452
rect 273312 59440 273318 59492
rect 273898 59440 273904 59492
rect 273956 59480 273962 59492
rect 276658 59480 276664 59492
rect 273956 59452 276664 59480
rect 273956 59440 273962 59452
rect 276658 59440 276664 59452
rect 276716 59440 276722 59492
rect 308490 59440 308496 59492
rect 308548 59480 308554 59492
rect 311158 59480 311164 59492
rect 308548 59452 311164 59480
rect 308548 59440 308554 59452
rect 311158 59440 311164 59452
rect 311216 59440 311222 59492
rect 329098 59440 329104 59492
rect 329156 59480 329162 59492
rect 331306 59480 331312 59492
rect 329156 59452 331312 59480
rect 329156 59440 329162 59452
rect 331306 59440 331312 59452
rect 331364 59440 331370 59492
rect 344738 59440 344744 59492
rect 344796 59480 344802 59492
rect 346486 59480 346492 59492
rect 344796 59452 346492 59480
rect 344796 59440 344802 59452
rect 346486 59440 346492 59452
rect 346544 59440 346550 59492
rect 351362 59440 351368 59492
rect 351420 59480 351426 59492
rect 353570 59480 353576 59492
rect 351420 59452 353576 59480
rect 351420 59440 351426 59452
rect 353570 59440 353576 59452
rect 353628 59440 353634 59492
rect 372706 59440 372712 59492
rect 372764 59480 372770 59492
rect 373994 59480 374000 59492
rect 372764 59452 374000 59480
rect 372764 59440 372770 59452
rect 373994 59440 374000 59452
rect 374052 59440 374058 59492
rect 398098 59440 398104 59492
rect 398156 59480 398162 59492
rect 401042 59480 401048 59492
rect 398156 59452 401048 59480
rect 398156 59440 398162 59452
rect 401042 59440 401048 59452
rect 401100 59440 401106 59492
rect 408126 59440 408132 59492
rect 408184 59480 408190 59492
rect 409874 59480 409880 59492
rect 408184 59452 409880 59480
rect 408184 59440 408190 59452
rect 409874 59440 409880 59452
rect 409932 59440 409938 59492
rect 428734 59440 428740 59492
rect 428792 59480 428798 59492
rect 430666 59480 430672 59492
rect 428792 59452 430672 59480
rect 428792 59440 428798 59452
rect 430666 59440 430672 59452
rect 430724 59440 430730 59492
rect 432046 59440 432052 59492
rect 432104 59480 432110 59492
rect 433426 59480 433432 59492
rect 432104 59452 433432 59480
rect 432104 59440 432110 59452
rect 433426 59440 433432 59452
rect 433484 59440 433490 59492
rect 455046 59440 455052 59492
rect 455104 59480 455110 59492
rect 456978 59480 456984 59492
rect 455104 59452 456984 59480
rect 455104 59440 455110 59452
rect 456978 59440 456984 59452
rect 457036 59440 457042 59492
rect 459186 59440 459192 59492
rect 459244 59480 459250 59492
rect 461210 59480 461216 59492
rect 459244 59452 461216 59480
rect 459244 59440 459250 59452
rect 461210 59440 461216 59452
rect 461268 59440 461274 59492
rect 188764 59384 190454 59412
rect 188764 59372 188770 59384
rect 306834 59304 306840 59356
rect 306892 59344 306898 59356
rect 308398 59344 308404 59356
rect 306892 59316 308404 59344
rect 306892 59304 306898 59316
rect 308398 59304 308404 59316
rect 308456 59304 308462 59356
rect 310514 59304 310520 59356
rect 310572 59344 310578 59356
rect 316954 59344 316960 59356
rect 310572 59316 316960 59344
rect 310572 59304 310578 59316
rect 316954 59304 316960 59316
rect 317012 59304 317018 59356
rect 325786 59304 325792 59356
rect 325844 59344 325850 59356
rect 327166 59344 327172 59356
rect 325844 59316 327172 59344
rect 325844 59304 325850 59316
rect 327166 59304 327172 59316
rect 327224 59304 327230 59356
rect 384114 59304 384120 59356
rect 384172 59344 384178 59356
rect 385678 59344 385684 59356
rect 384172 59316 385684 59344
rect 384172 59304 384178 59316
rect 385678 59304 385684 59316
rect 385736 59304 385742 59356
rect 123478 59236 123484 59288
rect 123536 59276 123542 59288
rect 126146 59276 126152 59288
rect 123536 59248 126152 59276
rect 123536 59236 123542 59248
rect 126146 59236 126152 59248
rect 126204 59236 126210 59288
rect 82078 58964 82084 59016
rect 82136 59004 82142 59016
rect 84194 59004 84200 59016
rect 82136 58976 84200 59004
rect 82136 58964 82142 58976
rect 84194 58964 84200 58976
rect 84252 58964 84258 59016
rect 401594 58964 401600 59016
rect 401652 59004 401658 59016
rect 405734 59004 405740 59016
rect 401652 58976 405740 59004
rect 401652 58964 401658 58976
rect 405734 58964 405740 58976
rect 405792 58964 405798 59016
rect 147582 58896 147588 58948
rect 147640 58936 147646 58948
rect 148686 58936 148692 58948
rect 147640 58908 148692 58936
rect 147640 58896 147646 58908
rect 148686 58896 148692 58908
rect 148744 58896 148750 58948
rect 251174 58896 251180 58948
rect 251232 58936 251238 58948
rect 330294 58936 330300 58948
rect 251232 58908 330300 58936
rect 251232 58896 251238 58908
rect 330294 58896 330300 58908
rect 330352 58896 330358 58948
rect 383654 58896 383660 58948
rect 383712 58936 383718 58948
rect 483014 58936 483020 58948
rect 383712 58908 483020 58936
rect 383712 58896 383718 58908
rect 483014 58896 483020 58908
rect 483072 58896 483078 58948
rect 320174 58828 320180 58880
rect 320232 58868 320238 58880
rect 419534 58868 419540 58880
rect 320232 58840 419540 58868
rect 320232 58828 320238 58840
rect 419534 58828 419540 58840
rect 419592 58828 419598 58880
rect 162854 58760 162860 58812
rect 162912 58800 162918 58812
rect 244182 58800 244188 58812
rect 162912 58772 244188 58800
rect 162912 58760 162918 58772
rect 244182 58760 244188 58772
rect 244240 58760 244246 58812
rect 271874 58760 271880 58812
rect 271932 58800 271938 58812
rect 513374 58800 513380 58812
rect 271932 58772 513380 58800
rect 271932 58760 271938 58772
rect 513374 58760 513380 58772
rect 513432 58760 513438 58812
rect 56594 58692 56600 58744
rect 56652 58732 56658 58744
rect 78582 58732 78588 58744
rect 56652 58704 78588 58732
rect 56652 58692 56658 58704
rect 78582 58692 78588 58704
rect 78640 58692 78646 58744
rect 193214 58692 193220 58744
rect 193272 58732 193278 58744
rect 449710 58732 449716 58744
rect 193272 58704 449716 58732
rect 193272 58692 193278 58704
rect 449710 58692 449716 58704
rect 449768 58692 449774 58744
rect 7558 58624 7564 58676
rect 7616 58664 7622 58676
rect 142062 58664 142068 58676
rect 7616 58636 142068 58664
rect 7616 58624 7622 58636
rect 142062 58624 142068 58636
rect 142120 58624 142126 58676
rect 157242 58624 157248 58676
rect 157300 58664 157306 58676
rect 546494 58664 546500 58676
rect 157300 58636 546500 58664
rect 157300 58624 157306 58636
rect 546494 58624 546500 58636
rect 546552 58624 546558 58676
rect 80882 58488 80888 58540
rect 80940 58528 80946 58540
rect 83274 58528 83280 58540
rect 80940 58500 83280 58528
rect 80940 58488 80946 58500
rect 83274 58488 83280 58500
rect 83332 58488 83338 58540
rect 291746 58488 291752 58540
rect 291804 58528 291810 58540
rect 293218 58528 293224 58540
rect 291804 58500 293224 58528
rect 291804 58488 291810 58500
rect 293218 58488 293224 58500
rect 293276 58488 293282 58540
rect 293402 58488 293408 58540
rect 293460 58528 293466 58540
rect 294782 58528 294788 58540
rect 293460 58500 294788 58528
rect 293460 58488 293466 58500
rect 294782 58488 294788 58500
rect 294840 58488 294846 58540
rect 148686 58352 148692 58404
rect 148744 58392 148750 58404
rect 149974 58392 149980 58404
rect 148744 58364 149980 58392
rect 148744 58352 148750 58364
rect 149974 58352 149980 58364
rect 150032 58352 150038 58404
rect 314654 57536 314660 57588
rect 314712 57576 314718 57588
rect 328454 57576 328460 57588
rect 314712 57548 328460 57576
rect 314712 57536 314718 57548
rect 328454 57536 328460 57548
rect 328512 57536 328518 57588
rect 331214 57536 331220 57588
rect 331272 57576 331278 57588
rect 416866 57576 416872 57588
rect 331272 57548 416872 57576
rect 331272 57536 331278 57548
rect 416866 57536 416872 57548
rect 416924 57536 416930 57588
rect 233234 57468 233240 57520
rect 233292 57508 233298 57520
rect 335354 57508 335360 57520
rect 233292 57480 335360 57508
rect 233292 57468 233298 57480
rect 335354 57468 335360 57480
rect 335412 57468 335418 57520
rect 382274 57468 382280 57520
rect 382332 57508 382338 57520
rect 489914 57508 489920 57520
rect 382332 57480 489920 57508
rect 382332 57468 382338 57480
rect 489914 57468 489920 57480
rect 489972 57468 489978 57520
rect 190362 57400 190368 57452
rect 190420 57440 190426 57452
rect 393314 57440 393320 57452
rect 190420 57412 393320 57440
rect 190420 57400 190426 57412
rect 393314 57400 393320 57412
rect 393372 57400 393378 57452
rect 273254 57332 273260 57384
rect 273312 57372 273318 57384
rect 506474 57372 506480 57384
rect 273312 57344 506480 57372
rect 273312 57332 273318 57344
rect 506474 57332 506480 57344
rect 506532 57332 506538 57384
rect 34514 57264 34520 57316
rect 34572 57304 34578 57316
rect 110322 57304 110328 57316
rect 34572 57276 110328 57304
rect 34572 57264 34578 57276
rect 110322 57264 110328 57276
rect 110380 57264 110386 57316
rect 195974 57264 195980 57316
rect 196032 57304 196038 57316
rect 451274 57304 451280 57316
rect 196032 57276 451280 57304
rect 196032 57264 196038 57276
rect 451274 57264 451280 57276
rect 451332 57264 451338 57316
rect 51074 57196 51080 57248
rect 51132 57236 51138 57248
rect 131114 57236 131120 57248
rect 51132 57208 131120 57236
rect 51132 57196 51138 57208
rect 131114 57196 131120 57208
rect 131172 57196 131178 57248
rect 164050 57196 164056 57248
rect 164108 57236 164114 57248
rect 517514 57236 517520 57248
rect 164108 57208 517520 57236
rect 164108 57196 164114 57208
rect 517514 57196 517520 57208
rect 517572 57196 517578 57248
rect 349154 56176 349160 56228
rect 349212 56216 349218 56228
rect 412910 56216 412916 56228
rect 349212 56188 412916 56216
rect 349212 56176 349218 56188
rect 412910 56176 412916 56188
rect 412968 56176 412974 56228
rect 172514 56108 172520 56160
rect 172572 56148 172578 56160
rect 348418 56148 348424 56160
rect 172572 56120 348424 56148
rect 172572 56108 172578 56120
rect 348418 56108 348424 56120
rect 348476 56108 348482 56160
rect 380802 56108 380808 56160
rect 380860 56148 380866 56160
rect 500954 56148 500960 56160
rect 380860 56120 500960 56148
rect 380860 56108 380866 56120
rect 500954 56108 500960 56120
rect 501012 56108 501018 56160
rect 194410 56040 194416 56092
rect 194468 56080 194474 56092
rect 386414 56080 386420 56092
rect 194468 56052 386420 56080
rect 194468 56040 194474 56052
rect 386414 56040 386420 56052
rect 386472 56040 386478 56092
rect 274634 55972 274640 56024
rect 274692 56012 274698 56024
rect 502334 56012 502340 56024
rect 274692 55984 502340 56012
rect 274692 55972 274698 55984
rect 502334 55972 502340 55984
rect 502392 55972 502398 56024
rect 209774 55904 209780 55956
rect 209832 55944 209838 55956
rect 447134 55944 447140 55956
rect 209832 55916 447140 55944
rect 209832 55904 209838 55916
rect 447134 55904 447140 55916
rect 447192 55904 447198 55956
rect 53834 55836 53840 55888
rect 53892 55876 53898 55888
rect 132034 55876 132040 55888
rect 53892 55848 132040 55876
rect 53892 55836 53898 55848
rect 132034 55836 132040 55848
rect 132092 55836 132098 55888
rect 162762 55836 162768 55888
rect 162820 55876 162826 55888
rect 524414 55876 524420 55888
rect 162820 55848 524420 55876
rect 162820 55836 162826 55848
rect 524414 55836 524420 55848
rect 524472 55836 524478 55888
rect 205450 54748 205456 54800
rect 205508 54788 205514 54800
rect 329834 54788 329840 54800
rect 205508 54760 329840 54788
rect 205508 54748 205514 54760
rect 329834 54748 329840 54760
rect 329892 54748 329898 54800
rect 376754 54748 376760 54800
rect 376812 54788 376818 54800
rect 408678 54788 408684 54800
rect 376812 54760 408684 54788
rect 376812 54748 376818 54760
rect 408678 54748 408684 54760
rect 408736 54748 408742 54800
rect 284294 54680 284300 54732
rect 284352 54720 284358 54732
rect 459554 54720 459560 54732
rect 284352 54692 459560 54720
rect 284352 54680 284358 54692
rect 459554 54680 459560 54692
rect 459612 54680 459618 54732
rect 226150 54612 226156 54664
rect 226208 54652 226214 54664
rect 241514 54652 241520 54664
rect 226208 54624 241520 54652
rect 226208 54612 226214 54624
rect 241514 54612 241520 54624
rect 241572 54612 241578 54664
rect 252554 54612 252560 54664
rect 252612 54652 252618 54664
rect 437474 54652 437480 54664
rect 252612 54624 437480 54652
rect 252612 54612 252618 54624
rect 437474 54612 437480 54624
rect 437532 54612 437538 54664
rect 110506 54544 110512 54596
rect 110564 54584 110570 54596
rect 118142 54584 118148 54596
rect 110564 54556 118148 54584
rect 110564 54544 110570 54556
rect 118142 54544 118148 54556
rect 118200 54544 118206 54596
rect 126974 54544 126980 54596
rect 127032 54584 127038 54596
rect 361574 54584 361580 54596
rect 127032 54556 361580 54584
rect 127032 54544 127038 54556
rect 361574 54544 361580 54556
rect 361632 54544 361638 54596
rect 373994 54544 374000 54596
rect 374052 54584 374058 54596
rect 525794 54584 525800 54596
rect 374052 54556 525800 54584
rect 374052 54544 374058 54556
rect 525794 54544 525800 54556
rect 525852 54544 525858 54596
rect 33134 54476 33140 54528
rect 33192 54516 33198 54528
rect 136082 54516 136088 54528
rect 33192 54488 136088 54516
rect 33192 54476 33198 54488
rect 136082 54476 136088 54488
rect 136140 54476 136146 54528
rect 180794 54476 180800 54528
rect 180852 54516 180858 54528
rect 239582 54516 239588 54528
rect 180852 54488 239588 54516
rect 180852 54476 180858 54488
rect 239582 54476 239588 54488
rect 239640 54476 239646 54528
rect 253842 54476 253848 54528
rect 253900 54516 253906 54528
rect 572714 54516 572720 54528
rect 253900 54488 572720 54516
rect 253900 54476 253906 54488
rect 572714 54476 572720 54488
rect 572772 54476 572778 54528
rect 308582 53388 308588 53440
rect 308640 53428 308646 53440
rect 360194 53428 360200 53440
rect 308640 53400 360200 53428
rect 308640 53388 308646 53400
rect 360194 53388 360200 53400
rect 360252 53388 360258 53440
rect 225966 53320 225972 53372
rect 226024 53360 226030 53372
rect 237374 53360 237380 53372
rect 226024 53332 237380 53360
rect 226024 53320 226030 53332
rect 237374 53320 237380 53332
rect 237432 53320 237438 53372
rect 258074 53320 258080 53372
rect 258132 53360 258138 53372
rect 331490 53360 331496 53372
rect 258132 53332 331496 53360
rect 258132 53320 258138 53332
rect 331490 53320 331496 53332
rect 331548 53320 331554 53372
rect 205634 53252 205640 53304
rect 205692 53292 205698 53304
rect 234062 53292 234068 53304
rect 205692 53264 234068 53292
rect 205692 53252 205698 53264
rect 234062 53252 234068 53264
rect 234120 53252 234126 53304
rect 288434 53252 288440 53304
rect 288492 53292 288498 53304
rect 445754 53292 445760 53304
rect 288492 53264 445760 53292
rect 288492 53252 288498 53264
rect 445754 53252 445760 53264
rect 445812 53252 445818 53304
rect 197078 53184 197084 53236
rect 197136 53224 197142 53236
rect 365714 53224 365720 53236
rect 197136 53196 365720 53224
rect 197136 53184 197142 53196
rect 365714 53184 365720 53196
rect 365772 53184 365778 53236
rect 372614 53184 372620 53236
rect 372672 53224 372678 53236
rect 532694 53224 532700 53236
rect 372672 53196 532700 53224
rect 372672 53184 372678 53196
rect 532694 53184 532700 53196
rect 532752 53184 532758 53236
rect 222010 53116 222016 53168
rect 222068 53156 222074 53168
rect 255314 53156 255320 53168
rect 222068 53128 255320 53156
rect 222068 53116 222074 53128
rect 255314 53116 255320 53128
rect 255372 53116 255378 53168
rect 259454 53116 259460 53168
rect 259512 53156 259518 53168
rect 436186 53156 436192 53168
rect 259512 53128 436192 53156
rect 259512 53116 259518 53128
rect 436186 53116 436192 53128
rect 436244 53116 436250 53168
rect 57974 53048 57980 53100
rect 58032 53088 58038 53100
rect 130562 53088 130568 53100
rect 58032 53060 130568 53088
rect 58032 53048 58038 53060
rect 130562 53048 130568 53060
rect 130620 53048 130626 53100
rect 146294 53048 146300 53100
rect 146352 53088 146358 53100
rect 462314 53088 462320 53100
rect 146352 53060 462320 53088
rect 146352 53048 146358 53060
rect 462314 53048 462320 53060
rect 462372 53048 462378 53100
rect 298922 52028 298928 52080
rect 298980 52068 298986 52080
rect 398834 52068 398840 52080
rect 298980 52040 398840 52068
rect 298980 52028 298986 52040
rect 398834 52028 398840 52040
rect 398892 52028 398898 52080
rect 235994 51960 236000 52012
rect 236052 52000 236058 52012
rect 336918 52000 336924 52012
rect 236052 51972 336924 52000
rect 236052 51960 236058 51972
rect 336918 51960 336924 51972
rect 336976 51960 336982 52012
rect 371326 51960 371332 52012
rect 371384 52000 371390 52012
rect 539594 52000 539600 52012
rect 371384 51972 539600 52000
rect 371384 51960 371390 51972
rect 539594 51960 539600 51972
rect 539652 51960 539658 52012
rect 263594 51892 263600 51944
rect 263652 51932 263658 51944
rect 434714 51932 434720 51944
rect 263652 51904 434720 51932
rect 263652 51892 263658 51904
rect 434714 51892 434720 51904
rect 434772 51892 434778 51944
rect 183370 51824 183376 51876
rect 183428 51864 183434 51876
rect 422294 51864 422300 51876
rect 183428 51836 422300 51864
rect 183428 51824 183434 51836
rect 422294 51824 422300 51836
rect 422352 51824 422358 51876
rect 143534 51756 143540 51808
rect 143592 51796 143598 51808
rect 463786 51796 463792 51808
rect 143592 51768 463792 51796
rect 143592 51756 143598 51768
rect 463786 51756 463792 51768
rect 463844 51756 463850 51808
rect 16574 51688 16580 51740
rect 16632 51728 16638 51740
rect 140682 51728 140688 51740
rect 16632 51700 140688 51728
rect 16632 51688 16638 51700
rect 140682 51688 140688 51700
rect 140740 51688 140746 51740
rect 158622 51688 158628 51740
rect 158680 51728 158686 51740
rect 528554 51728 528560 51740
rect 158680 51700 528560 51728
rect 158680 51688 158686 51700
rect 528554 51688 528560 51700
rect 528612 51688 528618 51740
rect 203978 50600 203984 50652
rect 204036 50640 204042 50652
rect 332594 50640 332600 50652
rect 204036 50612 332600 50640
rect 204036 50600 204042 50612
rect 332594 50600 332600 50612
rect 332652 50600 332658 50652
rect 380894 50600 380900 50652
rect 380952 50640 380958 50652
rect 408494 50640 408500 50652
rect 380952 50612 408500 50640
rect 380952 50600 380958 50612
rect 408494 50600 408500 50612
rect 408552 50600 408558 50652
rect 286502 50532 286508 50584
rect 286560 50572 286566 50584
rect 457070 50572 457076 50584
rect 286560 50544 457076 50572
rect 286560 50532 286566 50544
rect 457070 50532 457076 50544
rect 457128 50532 457134 50584
rect 204254 50464 204260 50516
rect 204312 50504 204318 50516
rect 343634 50504 343640 50516
rect 204312 50476 343640 50504
rect 204312 50464 204318 50476
rect 343634 50464 343640 50476
rect 343692 50464 343698 50516
rect 370682 50464 370688 50516
rect 370740 50504 370746 50516
rect 543734 50504 543740 50516
rect 370740 50476 543740 50504
rect 370740 50464 370746 50476
rect 543734 50464 543740 50476
rect 543792 50464 543798 50516
rect 20714 50396 20720 50448
rect 20772 50436 20778 50448
rect 138842 50436 138848 50448
rect 20772 50408 138848 50436
rect 20772 50396 20778 50408
rect 138842 50396 138848 50408
rect 138900 50396 138906 50448
rect 146938 50396 146944 50448
rect 146996 50436 147002 50448
rect 247862 50436 247868 50448
rect 146996 50408 247868 50436
rect 146996 50396 147002 50408
rect 247862 50396 247868 50408
rect 247920 50396 247926 50448
rect 278130 50396 278136 50448
rect 278188 50436 278194 50448
rect 488534 50436 488540 50448
rect 278188 50408 488540 50436
rect 278188 50396 278194 50408
rect 488534 50396 488540 50408
rect 488592 50396 488598 50448
rect 137278 50328 137284 50380
rect 137336 50368 137342 50380
rect 465074 50368 465080 50380
rect 137336 50340 465080 50368
rect 137336 50328 137342 50340
rect 465074 50328 465080 50340
rect 465132 50328 465138 50380
rect 208210 49308 208216 49360
rect 208268 49348 208274 49360
rect 316034 49348 316040 49360
rect 208268 49320 316040 49348
rect 208268 49308 208274 49320
rect 316034 49308 316040 49320
rect 316092 49308 316098 49360
rect 394694 49308 394700 49360
rect 394752 49348 394758 49360
rect 404354 49348 404360 49360
rect 394752 49320 404360 49348
rect 394752 49308 394758 49320
rect 404354 49308 404360 49320
rect 404412 49308 404418 49360
rect 290642 49240 290648 49292
rect 290700 49280 290706 49292
rect 438854 49280 438860 49292
rect 290700 49252 438860 49280
rect 290700 49240 290706 49252
rect 438854 49240 438860 49252
rect 438912 49240 438918 49292
rect 256694 49172 256700 49224
rect 256752 49212 256758 49224
rect 436370 49212 436376 49224
rect 256752 49184 436376 49212
rect 256752 49172 256758 49184
rect 436370 49172 436376 49184
rect 436428 49172 436434 49224
rect 136634 49104 136640 49156
rect 136692 49144 136698 49156
rect 358906 49144 358912 49156
rect 136692 49116 358912 49144
rect 136692 49104 136698 49116
rect 358906 49104 358912 49116
rect 358964 49104 358970 49156
rect 369118 49104 369124 49156
rect 369176 49144 369182 49156
rect 550634 49144 550640 49156
rect 369176 49116 550640 49144
rect 369176 49104 369182 49116
rect 550634 49104 550640 49116
rect 550692 49104 550698 49156
rect 186130 49036 186136 49088
rect 186188 49076 186194 49088
rect 411254 49076 411260 49088
rect 186188 49048 411260 49076
rect 186188 49036 186194 49048
rect 411254 49036 411260 49048
rect 411312 49036 411318 49088
rect 28994 48968 29000 49020
rect 29052 49008 29058 49020
rect 137370 49008 137376 49020
rect 29052 48980 137376 49008
rect 29052 48968 29058 48980
rect 137370 48968 137376 48980
rect 137428 48968 137434 49020
rect 150434 48968 150440 49020
rect 150492 49008 150498 49020
rect 461026 49008 461032 49020
rect 150492 48980 461032 49008
rect 150492 48968 150498 48980
rect 461026 48968 461032 48980
rect 461084 48968 461090 49020
rect 204162 47880 204168 47932
rect 204220 47920 204226 47932
rect 336734 47920 336740 47932
rect 204220 47892 336740 47920
rect 204220 47880 204226 47892
rect 336734 47880 336740 47892
rect 336792 47880 336798 47932
rect 168374 47812 168380 47864
rect 168432 47852 168438 47864
rect 351914 47852 351920 47864
rect 168432 47824 351920 47852
rect 168432 47812 168438 47824
rect 351914 47812 351920 47824
rect 351972 47812 351978 47864
rect 398282 47812 398288 47864
rect 398340 47852 398346 47864
rect 423674 47852 423680 47864
rect 398340 47824 423680 47852
rect 398340 47812 398346 47824
rect 423674 47812 423680 47824
rect 423732 47812 423738 47864
rect 242894 47744 242900 47796
rect 242952 47784 242958 47796
rect 440234 47784 440240 47796
rect 242952 47756 440240 47784
rect 242952 47744 242958 47756
rect 440234 47744 440240 47756
rect 440292 47744 440298 47796
rect 154574 47676 154580 47728
rect 154632 47716 154638 47728
rect 354858 47716 354864 47728
rect 154632 47688 354864 47716
rect 154632 47676 154638 47688
rect 354858 47676 354864 47688
rect 354916 47676 354922 47728
rect 367922 47676 367928 47728
rect 367980 47716 367986 47728
rect 554774 47716 554780 47728
rect 367980 47688 554780 47716
rect 367980 47676 367986 47688
rect 554774 47676 554780 47688
rect 554832 47676 554838 47728
rect 279418 47608 279424 47660
rect 279476 47648 279482 47660
rect 484394 47648 484400 47660
rect 279476 47620 484400 47648
rect 279476 47608 279482 47620
rect 484394 47608 484400 47620
rect 484452 47608 484458 47660
rect 26234 47540 26240 47592
rect 26292 47580 26298 47592
rect 138658 47580 138664 47592
rect 26292 47552 138664 47580
rect 26292 47540 26298 47552
rect 138658 47540 138664 47552
rect 138716 47540 138722 47592
rect 185946 47540 185952 47592
rect 186004 47580 186010 47592
rect 415394 47580 415400 47592
rect 186004 47552 415400 47580
rect 186004 47540 186010 47552
rect 415394 47540 415400 47552
rect 415452 47540 415458 47592
rect 308398 46520 308404 46572
rect 308456 46560 308462 46572
rect 357434 46560 357440 46572
rect 308456 46532 357440 46560
rect 308456 46520 308462 46532
rect 357434 46520 357440 46532
rect 357492 46520 357498 46572
rect 276014 46452 276020 46504
rect 276072 46492 276078 46504
rect 327166 46492 327172 46504
rect 276072 46464 327172 46492
rect 276072 46452 276078 46464
rect 327166 46452 327172 46464
rect 327224 46452 327230 46504
rect 387242 46452 387248 46504
rect 387300 46492 387306 46504
rect 473354 46492 473360 46504
rect 387300 46464 473360 46492
rect 387300 46452 387306 46464
rect 473354 46452 473360 46464
rect 473412 46452 473418 46504
rect 296990 46384 296996 46436
rect 297048 46424 297054 46436
rect 407114 46424 407120 46436
rect 297048 46396 407120 46424
rect 297048 46384 297054 46396
rect 407114 46384 407120 46396
rect 407172 46384 407178 46436
rect 161474 46316 161480 46368
rect 161532 46356 161538 46368
rect 353386 46356 353392 46368
rect 161532 46328 353392 46356
rect 161532 46316 161538 46328
rect 353386 46316 353392 46328
rect 353444 46316 353450 46368
rect 366542 46316 366548 46368
rect 366600 46356 366606 46368
rect 561674 46356 561680 46368
rect 366600 46328 561680 46356
rect 366600 46316 366606 46328
rect 561674 46316 561680 46328
rect 561732 46316 561738 46368
rect 224954 46248 224960 46300
rect 225012 46288 225018 46300
rect 444466 46288 444472 46300
rect 225012 46260 444472 46288
rect 225012 46248 225018 46260
rect 444466 46248 444472 46260
rect 444524 46248 444530 46300
rect 35894 46180 35900 46232
rect 35952 46220 35958 46232
rect 135898 46220 135904 46232
rect 35952 46192 135904 46220
rect 35952 46180 35958 46192
rect 135898 46180 135904 46192
rect 135956 46180 135962 46232
rect 154298 46180 154304 46232
rect 154356 46220 154362 46232
rect 548518 46220 548524 46232
rect 154356 46192 548524 46220
rect 154356 46180 154362 46192
rect 548518 46180 548524 46192
rect 548576 46180 548582 46232
rect 271874 45160 271880 45212
rect 271932 45200 271938 45212
rect 328638 45200 328644 45212
rect 271932 45172 328644 45200
rect 271932 45160 271938 45172
rect 328638 45160 328644 45172
rect 328696 45160 328702 45212
rect 307202 45092 307208 45144
rect 307260 45132 307266 45144
rect 364334 45132 364340 45144
rect 307260 45104 364340 45132
rect 307260 45092 307266 45104
rect 364334 45092 364340 45104
rect 364392 45092 364398 45144
rect 217870 45024 217876 45076
rect 217928 45064 217934 45076
rect 273254 45064 273260 45076
rect 217928 45036 273260 45064
rect 217928 45024 217934 45036
rect 273254 45024 273260 45036
rect 273312 45024 273318 45076
rect 290458 45024 290464 45076
rect 290516 45064 290522 45076
rect 434714 45064 434720 45076
rect 290516 45036 434720 45064
rect 290516 45024 290522 45036
rect 434714 45024 434720 45036
rect 434772 45024 434778 45076
rect 197262 44956 197268 45008
rect 197320 44996 197326 45008
rect 361574 44996 361580 45008
rect 197320 44968 361580 44996
rect 197320 44956 197326 44968
rect 361574 44956 361580 44968
rect 361632 44956 361638 45008
rect 388622 44956 388628 45008
rect 388680 44996 388686 45008
rect 465258 44996 465264 45008
rect 388680 44968 465264 44996
rect 388680 44956 388686 44968
rect 465258 44956 465264 44968
rect 465316 44956 465322 45008
rect 165614 44888 165620 44940
rect 165672 44928 165678 44940
rect 353570 44928 353576 44940
rect 165672 44900 353576 44928
rect 165672 44888 165678 44900
rect 353570 44888 353576 44900
rect 353628 44888 353634 44940
rect 366358 44888 366364 44940
rect 366416 44928 366422 44940
rect 564434 44928 564440 44940
rect 366416 44900 564440 44928
rect 366416 44888 366422 44900
rect 564434 44888 564440 44900
rect 564492 44888 564498 44940
rect 40034 44820 40040 44872
rect 40092 44860 40098 44872
rect 134702 44860 134708 44872
rect 40092 44832 134708 44860
rect 40092 44820 40098 44832
rect 134702 44820 134708 44832
rect 134760 44820 134766 44872
rect 220814 44820 220820 44872
rect 220872 44860 220878 44872
rect 444374 44860 444380 44872
rect 220872 44832 444380 44860
rect 220872 44820 220878 44832
rect 444374 44820 444380 44832
rect 444432 44820 444438 44872
rect 201310 43732 201316 43784
rect 201368 43772 201374 43784
rect 343634 43772 343640 43784
rect 201368 43744 343640 43772
rect 201368 43732 201374 43744
rect 343634 43732 343640 43744
rect 343692 43732 343698 43784
rect 270494 43664 270500 43716
rect 270552 43704 270558 43716
rect 433426 43704 433432 43716
rect 270552 43676 433432 43704
rect 270552 43664 270558 43676
rect 433426 43664 433432 43676
rect 433484 43664 433490 43716
rect 158714 43596 158720 43648
rect 158772 43636 158778 43648
rect 354950 43636 354956 43648
rect 158772 43608 354956 43636
rect 158772 43596 158778 43608
rect 354950 43596 354956 43608
rect 355008 43596 355014 43648
rect 390002 43596 390008 43648
rect 390060 43636 390066 43648
rect 458174 43636 458180 43648
rect 390060 43608 458180 43636
rect 390060 43596 390066 43608
rect 458174 43596 458180 43608
rect 458232 43596 458238 43648
rect 181990 43528 181996 43580
rect 182048 43568 182054 43580
rect 431954 43568 431960 43580
rect 182048 43540 431960 43568
rect 182048 43528 182054 43540
rect 431954 43528 431960 43540
rect 432012 43528 432018 43580
rect 175274 43460 175280 43512
rect 175332 43500 175338 43512
rect 455506 43500 455512 43512
rect 175332 43472 455512 43500
rect 175332 43460 175338 43472
rect 455506 43460 455512 43472
rect 455564 43460 455570 43512
rect 11698 43392 11704 43444
rect 11756 43432 11762 43444
rect 115198 43432 115204 43444
rect 11756 43404 115204 43432
rect 11756 43392 11762 43404
rect 115198 43392 115204 43404
rect 115256 43392 115262 43444
rect 255130 43392 255136 43444
rect 255188 43432 255194 43444
rect 569954 43432 569960 43444
rect 255188 43404 569960 43432
rect 255188 43392 255194 43404
rect 569954 43392 569960 43404
rect 570012 43392 570018 43444
rect 209590 42372 209596 42424
rect 209648 42412 209654 42424
rect 307754 42412 307760 42424
rect 209648 42384 307760 42412
rect 209648 42372 209654 42384
rect 307754 42372 307760 42384
rect 307812 42372 307818 42424
rect 299474 42304 299480 42356
rect 299532 42344 299538 42356
rect 426526 42344 426532 42356
rect 299532 42316 426532 42344
rect 299532 42304 299538 42316
rect 426526 42304 426532 42316
rect 426584 42304 426590 42356
rect 195790 42236 195796 42288
rect 195848 42276 195854 42288
rect 372614 42276 372620 42288
rect 195848 42248 372620 42276
rect 195848 42236 195854 42248
rect 372614 42236 372620 42248
rect 372672 42236 372678 42288
rect 142798 42168 142804 42220
rect 142856 42208 142862 42220
rect 358814 42208 358820 42220
rect 142856 42180 358820 42208
rect 142856 42168 142862 42180
rect 358814 42168 358820 42180
rect 358872 42168 358878 42220
rect 392762 42168 392768 42220
rect 392820 42208 392826 42220
rect 448514 42208 448520 42220
rect 392820 42180 448520 42208
rect 392820 42168 392826 42180
rect 448514 42168 448520 42180
rect 448572 42168 448578 42220
rect 272518 42100 272524 42152
rect 272576 42140 272582 42152
rect 516134 42140 516140 42152
rect 272576 42112 516140 42140
rect 272576 42100 272582 42112
rect 516134 42100 516140 42112
rect 516192 42100 516198 42152
rect 3418 42032 3424 42084
rect 3476 42072 3482 42084
rect 142890 42072 142896 42084
rect 3476 42044 142896 42072
rect 3476 42032 3482 42044
rect 142890 42032 142896 42044
rect 142948 42032 142954 42084
rect 182174 42032 182180 42084
rect 182232 42072 182238 42084
rect 454034 42072 454040 42084
rect 182232 42044 454040 42072
rect 182232 42032 182238 42044
rect 454034 42032 454040 42044
rect 454092 42032 454098 42084
rect 253934 41012 253940 41064
rect 253992 41052 253998 41064
rect 332686 41052 332692 41064
rect 253992 41024 332692 41052
rect 253992 41012 253998 41024
rect 332686 41012 332692 41024
rect 332744 41012 332750 41064
rect 303062 40944 303068 40996
rect 303120 40984 303126 40996
rect 382274 40984 382280 40996
rect 303120 40956 382280 40984
rect 303120 40944 303126 40956
rect 382274 40944 382280 40956
rect 382332 40944 382338 40996
rect 193030 40876 193036 40928
rect 193088 40916 193094 40928
rect 379514 40916 379520 40928
rect 193088 40888 379520 40916
rect 193088 40876 193094 40888
rect 379514 40876 379520 40888
rect 379572 40876 379578 40928
rect 387058 40876 387064 40928
rect 387116 40916 387122 40928
rect 476114 40916 476120 40928
rect 387116 40888 476120 40916
rect 387116 40876 387122 40888
rect 476114 40876 476120 40888
rect 476172 40876 476178 40928
rect 282362 40808 282368 40860
rect 282420 40848 282426 40860
rect 470594 40848 470600 40860
rect 282420 40820 470600 40848
rect 282420 40808 282426 40820
rect 470594 40808 470600 40820
rect 470652 40808 470658 40860
rect 178034 40740 178040 40792
rect 178092 40780 178098 40792
rect 455690 40780 455696 40792
rect 178092 40752 455696 40780
rect 178092 40740 178098 40752
rect 455690 40740 455696 40752
rect 455748 40740 455754 40792
rect 14458 40672 14464 40724
rect 14516 40712 14522 40724
rect 114002 40712 114008 40724
rect 14516 40684 114008 40712
rect 14516 40672 14522 40684
rect 114002 40672 114008 40684
rect 114060 40672 114066 40724
rect 139394 40672 139400 40724
rect 139452 40712 139458 40724
rect 463970 40712 463976 40724
rect 139452 40684 463976 40712
rect 139452 40672 139458 40684
rect 463970 40672 463976 40684
rect 464028 40672 464034 40724
rect 278774 39652 278780 39704
rect 278832 39692 278838 39704
rect 327350 39692 327356 39704
rect 278832 39664 327356 39692
rect 278832 39652 278838 39664
rect 327350 39652 327356 39664
rect 327408 39652 327414 39704
rect 216490 39584 216496 39636
rect 216548 39624 216554 39636
rect 284294 39624 284300 39636
rect 216548 39596 284300 39624
rect 216548 39584 216554 39596
rect 284294 39584 284300 39596
rect 284352 39584 284358 39636
rect 313274 39584 313280 39636
rect 313332 39624 313338 39636
rect 423766 39624 423772 39636
rect 313332 39596 423772 39624
rect 313332 39584 313338 39596
rect 423766 39584 423772 39596
rect 423824 39584 423830 39636
rect 195606 39516 195612 39568
rect 195664 39556 195670 39568
rect 368474 39556 368480 39568
rect 195664 39528 368480 39556
rect 195664 39516 195670 39528
rect 368474 39516 368480 39528
rect 368532 39516 368538 39568
rect 395338 39516 395344 39568
rect 395396 39556 395402 39568
rect 437474 39556 437480 39568
rect 395396 39528 437480 39556
rect 395396 39516 395402 39528
rect 437474 39516 437480 39528
rect 437532 39516 437538 39568
rect 212534 39448 212540 39500
rect 212592 39488 212598 39500
rect 232682 39488 232688 39500
rect 212592 39460 232688 39488
rect 212592 39448 212598 39460
rect 232682 39448 232688 39460
rect 232740 39448 232746 39500
rect 283558 39448 283564 39500
rect 283616 39488 283622 39500
rect 466454 39488 466460 39500
rect 283616 39460 466460 39488
rect 283616 39448 283622 39460
rect 466454 39448 466460 39460
rect 466512 39448 466518 39500
rect 221826 39380 221832 39432
rect 221884 39420 221890 39432
rect 259546 39420 259552 39432
rect 221884 39392 259552 39420
rect 221884 39380 221890 39392
rect 259546 39380 259552 39392
rect 259604 39380 259610 39432
rect 276842 39380 276848 39432
rect 276900 39420 276906 39432
rect 495434 39420 495440 39432
rect 276900 39392 495440 39420
rect 276900 39380 276906 39392
rect 495434 39380 495440 39392
rect 495492 39380 495498 39432
rect 18598 39312 18604 39364
rect 18656 39352 18662 39364
rect 113818 39352 113824 39364
rect 18656 39324 113824 39352
rect 18656 39312 18662 39324
rect 113818 39312 113824 39324
rect 113876 39312 113882 39364
rect 171134 39312 171140 39364
rect 171192 39352 171198 39364
rect 456978 39352 456984 39364
rect 171192 39324 456984 39352
rect 171192 39312 171198 39324
rect 456978 39312 456984 39324
rect 457036 39312 457042 39364
rect 282914 38224 282920 38276
rect 282972 38264 282978 38276
rect 325694 38264 325700 38276
rect 282972 38236 325700 38264
rect 282972 38224 282978 38236
rect 325694 38224 325700 38236
rect 325752 38224 325758 38276
rect 302234 38156 302240 38208
rect 302292 38196 302298 38208
rect 426434 38196 426440 38208
rect 302292 38168 426440 38196
rect 302292 38156 302298 38168
rect 426434 38156 426440 38168
rect 426492 38156 426498 38208
rect 199838 38088 199844 38140
rect 199896 38128 199902 38140
rect 350626 38128 350632 38140
rect 199896 38100 350632 38128
rect 199896 38088 199902 38100
rect 350626 38088 350632 38100
rect 350684 38088 350690 38140
rect 394142 38088 394148 38140
rect 394200 38128 394206 38140
rect 440234 38128 440240 38140
rect 394200 38100 440240 38128
rect 394200 38088 394206 38100
rect 440234 38088 440240 38100
rect 440292 38088 440298 38140
rect 276658 38020 276664 38072
rect 276716 38060 276722 38072
rect 498194 38060 498200 38072
rect 276716 38032 498200 38060
rect 276716 38020 276722 38032
rect 498194 38020 498200 38032
rect 498252 38020 498258 38072
rect 168466 37952 168472 38004
rect 168524 37992 168530 38004
rect 456794 37992 456800 38004
rect 168524 37964 456800 37992
rect 168524 37952 168530 37964
rect 456794 37952 456800 37964
rect 456852 37952 456858 38004
rect 27614 37884 27620 37936
rect 27672 37924 27678 37936
rect 111242 37924 111248 37936
rect 27672 37896 111248 37924
rect 27672 37884 27678 37896
rect 111242 37884 111248 37896
rect 111300 37884 111306 37936
rect 162670 37884 162676 37936
rect 162728 37924 162734 37936
rect 510614 37924 510620 37936
rect 162728 37896 510620 37924
rect 162728 37884 162734 37896
rect 510614 37884 510620 37896
rect 510672 37884 510678 37936
rect 296162 36864 296168 36916
rect 296220 36904 296226 36916
rect 410058 36904 410064 36916
rect 296220 36876 410064 36904
rect 296220 36864 296226 36876
rect 410058 36864 410064 36876
rect 410116 36864 410122 36916
rect 206922 36796 206928 36848
rect 206980 36836 206986 36848
rect 322934 36836 322940 36848
rect 206980 36808 322940 36836
rect 206980 36796 206986 36808
rect 322934 36796 322940 36808
rect 322992 36796 322998 36848
rect 176654 36728 176660 36780
rect 176712 36768 176718 36780
rect 350534 36768 350540 36780
rect 176712 36740 350540 36768
rect 176712 36728 176718 36740
rect 350534 36728 350540 36740
rect 350592 36728 350598 36780
rect 367738 36728 367744 36780
rect 367796 36768 367802 36780
rect 557534 36768 557540 36780
rect 367796 36740 557540 36768
rect 367796 36728 367802 36740
rect 557534 36728 557540 36740
rect 557592 36728 557598 36780
rect 141418 36660 141424 36712
rect 141476 36700 141482 36712
rect 249058 36700 249064 36712
rect 141476 36672 249064 36700
rect 141476 36660 141482 36672
rect 249058 36660 249064 36672
rect 249116 36660 249122 36712
rect 280982 36660 280988 36712
rect 281040 36700 281046 36712
rect 481634 36700 481640 36712
rect 281040 36672 481640 36700
rect 281040 36660 281046 36672
rect 481634 36660 481640 36672
rect 481692 36660 481698 36712
rect 187510 36592 187516 36644
rect 187568 36632 187574 36644
rect 404354 36632 404360 36644
rect 187568 36604 404360 36632
rect 187568 36592 187574 36604
rect 404354 36592 404360 36604
rect 404412 36592 404418 36644
rect 10318 36524 10324 36576
rect 10376 36564 10382 36576
rect 141510 36564 141516 36576
rect 10376 36536 141516 36564
rect 10376 36524 10382 36536
rect 141510 36524 141516 36536
rect 141568 36524 141574 36576
rect 218054 36524 218060 36576
rect 218112 36564 218118 36576
rect 445846 36564 445852 36576
rect 218112 36536 445852 36564
rect 218112 36524 218118 36536
rect 445846 36524 445852 36536
rect 445904 36524 445910 36576
rect 205266 35436 205272 35488
rect 205324 35476 205330 35488
rect 325694 35476 325700 35488
rect 205324 35448 325700 35476
rect 205324 35436 205330 35448
rect 325694 35436 325700 35448
rect 325752 35436 325758 35488
rect 391198 35436 391204 35488
rect 391256 35476 391262 35488
rect 455414 35476 455420 35488
rect 391256 35448 455420 35476
rect 391256 35436 391262 35448
rect 455414 35436 455420 35448
rect 455472 35436 455478 35488
rect 277394 35368 277400 35420
rect 277452 35408 277458 35420
rect 432046 35408 432052 35420
rect 277452 35380 432052 35408
rect 277452 35368 277458 35380
rect 432046 35368 432052 35380
rect 432104 35368 432110 35420
rect 164234 35300 164240 35352
rect 164292 35340 164298 35352
rect 458266 35340 458272 35352
rect 164292 35312 458272 35340
rect 164292 35300 164298 35312
rect 458266 35300 458272 35312
rect 458324 35300 458330 35352
rect 254946 35232 254952 35284
rect 255004 35272 255010 35284
rect 565814 35272 565820 35284
rect 255004 35244 565820 35272
rect 255004 35232 255010 35244
rect 565814 35232 565820 35244
rect 565872 35232 565878 35284
rect 43438 35164 43444 35216
rect 43496 35204 43502 35216
rect 107102 35204 107108 35216
rect 43496 35176 107108 35204
rect 43496 35164 43502 35176
rect 107102 35164 107108 35176
rect 107160 35164 107166 35216
rect 162486 35164 162492 35216
rect 162544 35204 162550 35216
rect 514754 35204 514760 35216
rect 162544 35176 514760 35204
rect 162544 35164 162550 35176
rect 514754 35164 514760 35176
rect 514812 35164 514818 35216
rect 315298 34076 315304 34128
rect 315356 34116 315362 34128
rect 332686 34116 332692 34128
rect 315356 34088 332692 34116
rect 315356 34076 315362 34088
rect 332686 34076 332692 34088
rect 332744 34076 332750 34128
rect 298738 34008 298744 34060
rect 298796 34048 298802 34060
rect 402974 34048 402980 34060
rect 298796 34020 402980 34048
rect 298796 34008 298802 34020
rect 402974 34008 402980 34020
rect 403032 34008 403038 34060
rect 267734 33940 267740 33992
rect 267792 33980 267798 33992
rect 328822 33980 328828 33992
rect 267792 33952 328828 33980
rect 267792 33940 267798 33952
rect 328822 33940 328828 33952
rect 328880 33940 328886 33992
rect 370498 33940 370504 33992
rect 370556 33980 370562 33992
rect 547874 33980 547880 33992
rect 370556 33952 547880 33980
rect 370556 33940 370562 33952
rect 547874 33940 547880 33952
rect 547932 33940 547938 33992
rect 213914 33872 213920 33924
rect 213972 33912 213978 33924
rect 447410 33912 447416 33924
rect 213972 33884 447416 33912
rect 213972 33872 213978 33884
rect 447410 33872 447416 33884
rect 447468 33872 447474 33924
rect 157334 33804 157340 33856
rect 157392 33844 157398 33856
rect 459738 33844 459744 33856
rect 157392 33816 459744 33844
rect 157392 33804 157398 33816
rect 459738 33804 459744 33816
rect 459796 33804 459802 33856
rect 49694 33736 49700 33788
rect 49752 33776 49758 33788
rect 79502 33776 79508 33788
rect 49752 33748 79508 33776
rect 49752 33736 49758 33748
rect 79502 33736 79508 33748
rect 79560 33736 79566 33788
rect 150250 33736 150256 33788
rect 150308 33776 150314 33788
rect 564526 33776 564532 33788
rect 150308 33748 564532 33776
rect 150308 33736 150314 33748
rect 564526 33736 564532 33748
rect 564584 33736 564590 33788
rect 300302 32716 300308 32768
rect 300360 32756 300366 32768
rect 396074 32756 396080 32768
rect 300360 32728 396080 32756
rect 300360 32716 300366 32728
rect 396074 32716 396080 32728
rect 396132 32716 396138 32768
rect 260834 32648 260840 32700
rect 260892 32688 260898 32700
rect 331306 32688 331312 32700
rect 260892 32660 331312 32688
rect 260892 32648 260898 32660
rect 331306 32648 331312 32660
rect 331364 32648 331370 32700
rect 374638 32648 374644 32700
rect 374696 32688 374702 32700
rect 529934 32688 529940 32700
rect 374696 32660 529940 32688
rect 374696 32648 374702 32660
rect 529934 32648 529940 32660
rect 529992 32648 529998 32700
rect 207014 32580 207020 32632
rect 207072 32620 207078 32632
rect 448790 32620 448796 32632
rect 207072 32592 448796 32620
rect 207072 32580 207078 32592
rect 448790 32580 448796 32592
rect 448848 32580 448854 32632
rect 179138 32512 179144 32564
rect 179196 32552 179202 32564
rect 440326 32552 440332 32564
rect 179196 32524 440332 32552
rect 179196 32512 179202 32524
rect 440326 32512 440332 32524
rect 440384 32512 440390 32564
rect 153194 32444 153200 32496
rect 153252 32484 153258 32496
rect 461210 32484 461216 32496
rect 153252 32456 461216 32484
rect 153252 32444 153258 32456
rect 461210 32444 461216 32456
rect 461268 32444 461274 32496
rect 157150 32376 157156 32428
rect 157208 32416 157214 32428
rect 539686 32416 539692 32428
rect 157208 32388 539692 32416
rect 157208 32376 157214 32388
rect 539686 32376 539692 32388
rect 539744 32376 539750 32428
rect 202782 31288 202788 31340
rect 202840 31328 202846 31340
rect 340874 31328 340880 31340
rect 202840 31300 340880 31328
rect 202840 31288 202846 31300
rect 340874 31288 340880 31300
rect 340932 31288 340938 31340
rect 373994 31288 374000 31340
rect 374052 31328 374058 31340
rect 409874 31328 409880 31340
rect 374052 31300 409880 31328
rect 374052 31288 374058 31300
rect 409874 31288 409880 31300
rect 409932 31288 409938 31340
rect 286318 31220 286324 31272
rect 286376 31260 286382 31272
rect 452654 31260 452660 31272
rect 286376 31232 452660 31260
rect 286376 31220 286382 31232
rect 452654 31220 452660 31232
rect 452712 31220 452718 31272
rect 179414 31152 179420 31204
rect 179472 31192 179478 31204
rect 349246 31192 349252 31204
rect 179472 31164 349252 31192
rect 179472 31152 179478 31164
rect 349246 31152 349252 31164
rect 349304 31152 349310 31204
rect 376202 31152 376208 31204
rect 376260 31192 376266 31204
rect 523034 31192 523040 31204
rect 376260 31164 523040 31192
rect 376260 31152 376266 31164
rect 523034 31152 523040 31164
rect 523092 31152 523098 31204
rect 219342 31084 219348 31136
rect 219400 31124 219406 31136
rect 269114 31124 269120 31136
rect 219400 31096 269120 31124
rect 219400 31084 219406 31096
rect 269114 31084 269120 31096
rect 269172 31084 269178 31136
rect 278038 31084 278044 31136
rect 278096 31124 278102 31136
rect 491294 31124 491300 31136
rect 278096 31096 491300 31124
rect 278096 31084 278102 31096
rect 491294 31084 491300 31096
rect 491352 31084 491358 31136
rect 202874 31016 202880 31068
rect 202932 31056 202938 31068
rect 448606 31056 448612 31068
rect 202932 31028 448612 31056
rect 202932 31016 202938 31028
rect 448606 31016 448612 31028
rect 448664 31016 448670 31068
rect 396902 29996 396908 30048
rect 396960 30036 396966 30048
rect 433334 30036 433340 30048
rect 396960 30008 433340 30036
rect 396960 29996 396966 30008
rect 433334 29996 433340 30008
rect 433392 29996 433398 30048
rect 208026 29928 208032 29980
rect 208084 29968 208090 29980
rect 318794 29968 318800 29980
rect 208084 29940 318800 29968
rect 208084 29928 208090 29940
rect 318794 29928 318800 29940
rect 318852 29928 318858 29980
rect 274634 29860 274640 29912
rect 274692 29900 274698 29912
rect 433610 29900 433616 29912
rect 274692 29872 433616 29900
rect 274692 29860 274698 29872
rect 433610 29860 433616 29872
rect 433668 29860 433674 29912
rect 198734 29792 198740 29844
rect 198792 29832 198798 29844
rect 235442 29832 235448 29844
rect 198792 29804 235448 29832
rect 198792 29792 198798 29804
rect 235442 29792 235448 29804
rect 235500 29792 235506 29844
rect 284938 29792 284944 29844
rect 284996 29832 285002 29844
rect 463694 29832 463700 29844
rect 284996 29804 463700 29832
rect 284996 29792 285002 29804
rect 463694 29792 463700 29804
rect 463752 29792 463758 29844
rect 184842 29724 184848 29776
rect 184900 29764 184906 29776
rect 418338 29764 418344 29776
rect 184900 29736 418344 29764
rect 184900 29724 184906 29736
rect 418338 29724 418344 29736
rect 418396 29724 418402 29776
rect 220630 29656 220636 29708
rect 220688 29696 220694 29708
rect 262214 29696 262220 29708
rect 220688 29668 262220 29696
rect 220688 29656 220694 29668
rect 262214 29656 262220 29668
rect 262272 29656 262278 29708
rect 269942 29656 269948 29708
rect 270000 29696 270006 29708
rect 527174 29696 527180 29708
rect 270000 29668 527180 29696
rect 270000 29656 270006 29668
rect 527174 29656 527180 29668
rect 527232 29656 527238 29708
rect 160094 29588 160100 29640
rect 160152 29628 160158 29640
rect 459922 29628 459928 29640
rect 160152 29600 459928 29628
rect 160152 29588 160158 29600
rect 459922 29588 459928 29600
rect 459980 29588 459986 29640
rect 333974 28500 333980 28552
rect 334032 28540 334038 28552
rect 418154 28540 418160 28552
rect 334032 28512 418160 28540
rect 334032 28500 334038 28512
rect 418154 28500 418160 28512
rect 418212 28500 418218 28552
rect 129734 28432 129740 28484
rect 129792 28472 129798 28484
rect 361758 28472 361764 28484
rect 129792 28444 361764 28472
rect 129792 28432 129798 28444
rect 361758 28432 361764 28444
rect 361816 28432 361822 28484
rect 380158 28432 380164 28484
rect 380216 28472 380222 28484
rect 505094 28472 505100 28484
rect 380216 28444 505100 28472
rect 380216 28432 380222 28444
rect 505094 28432 505100 28444
rect 505152 28432 505158 28484
rect 273898 28364 273904 28416
rect 273956 28404 273962 28416
rect 509234 28404 509240 28416
rect 273956 28376 509240 28404
rect 273956 28364 273962 28376
rect 509234 28364 509240 28376
rect 509292 28364 509298 28416
rect 200114 28296 200120 28348
rect 200172 28336 200178 28348
rect 449894 28336 449900 28348
rect 200172 28308 449900 28336
rect 200172 28296 200178 28308
rect 449894 28296 449900 28308
rect 449952 28296 449958 28348
rect 68830 28228 68836 28280
rect 68888 28268 68894 28280
rect 99374 28268 99380 28280
rect 68888 28240 99380 28268
rect 68888 28228 68894 28240
rect 99374 28228 99380 28240
rect 99432 28228 99438 28280
rect 150066 28228 150072 28280
rect 150124 28268 150130 28280
rect 566458 28268 566464 28280
rect 150124 28240 566464 28268
rect 150124 28228 150130 28240
rect 566458 28228 566464 28240
rect 566516 28228 566522 28280
rect 327074 27208 327080 27260
rect 327132 27248 327138 27260
rect 421098 27248 421104 27260
rect 327132 27220 421104 27248
rect 327132 27208 327138 27220
rect 421098 27208 421104 27220
rect 421156 27208 421162 27260
rect 215294 27140 215300 27192
rect 215352 27180 215358 27192
rect 340966 27180 340972 27192
rect 215352 27152 340972 27180
rect 215352 27140 215358 27152
rect 340966 27140 340972 27152
rect 341024 27140 341030 27192
rect 381538 27140 381544 27192
rect 381596 27180 381602 27192
rect 498286 27180 498292 27192
rect 381596 27152 498292 27180
rect 381596 27140 381602 27152
rect 498286 27140 498292 27152
rect 498344 27140 498350 27192
rect 188890 27072 188896 27124
rect 188948 27112 188954 27124
rect 400214 27112 400220 27124
rect 188948 27084 400220 27112
rect 188948 27072 188954 27084
rect 400214 27072 400220 27084
rect 400272 27072 400278 27124
rect 268562 27004 268568 27056
rect 268620 27044 268626 27056
rect 531314 27044 531320 27056
rect 268620 27016 531320 27044
rect 268620 27004 268626 27016
rect 531314 27004 531320 27016
rect 531372 27004 531378 27056
rect 128354 26936 128360 26988
rect 128412 26976 128418 26988
rect 466546 26976 466552 26988
rect 128412 26948 466552 26976
rect 128412 26936 128418 26948
rect 466546 26936 466552 26948
rect 466604 26936 466610 26988
rect 17954 26868 17960 26920
rect 18012 26908 18018 26920
rect 112438 26908 112444 26920
rect 18012 26880 112444 26908
rect 18012 26868 18018 26880
rect 112438 26868 112444 26880
rect 112496 26868 112502 26920
rect 147582 26868 147588 26920
rect 147640 26908 147646 26920
rect 578234 26908 578240 26920
rect 147640 26880 578240 26908
rect 147640 26868 147646 26880
rect 578234 26868 578240 26880
rect 578292 26868 578298 26920
rect 316862 25984 316868 26036
rect 316920 26024 316926 26036
rect 321554 26024 321560 26036
rect 316920 25996 321560 26024
rect 316920 25984 316926 25996
rect 321554 25984 321560 25996
rect 321612 25984 321618 26036
rect 242986 25848 242992 25900
rect 243044 25888 243050 25900
rect 335354 25888 335360 25900
rect 243044 25860 335360 25888
rect 243044 25848 243050 25860
rect 335354 25848 335360 25860
rect 335412 25848 335418 25900
rect 324314 25780 324320 25832
rect 324372 25820 324378 25832
rect 420914 25820 420920 25832
rect 324372 25792 420920 25820
rect 324372 25780 324378 25792
rect 420914 25780 420920 25792
rect 420972 25780 420978 25832
rect 198642 25712 198648 25764
rect 198700 25752 198706 25764
rect 357526 25752 357532 25764
rect 198700 25724 357532 25752
rect 198700 25712 198706 25724
rect 357526 25712 357532 25724
rect 357584 25712 357590 25764
rect 382918 25712 382924 25764
rect 382976 25752 382982 25764
rect 494054 25752 494060 25764
rect 382976 25724 494060 25752
rect 382976 25712 382982 25724
rect 494054 25712 494060 25724
rect 494112 25712 494118 25764
rect 271138 25644 271144 25696
rect 271196 25684 271202 25696
rect 520274 25684 520280 25696
rect 271196 25656 520280 25684
rect 271196 25644 271202 25656
rect 520274 25644 520280 25656
rect 520332 25644 520338 25696
rect 189074 25576 189080 25628
rect 189132 25616 189138 25628
rect 452930 25616 452936 25628
rect 189132 25588 452936 25616
rect 189132 25576 189138 25588
rect 452930 25576 452936 25588
rect 452988 25576 452994 25628
rect 90910 25508 90916 25560
rect 90968 25548 90974 25560
rect 111794 25548 111800 25560
rect 90968 25520 111800 25548
rect 90968 25508 90974 25520
rect 111794 25508 111800 25520
rect 111852 25508 111858 25560
rect 158346 25508 158352 25560
rect 158404 25548 158410 25560
rect 531406 25548 531412 25560
rect 158404 25520 531412 25548
rect 158404 25508 158410 25520
rect 531406 25508 531412 25520
rect 531464 25508 531470 25560
rect 264974 24420 264980 24472
rect 265032 24460 265038 24472
rect 329926 24460 329932 24472
rect 265032 24432 329932 24460
rect 265032 24420 265038 24432
rect 329926 24420 329932 24432
rect 329984 24420 329990 24472
rect 384298 24420 384304 24472
rect 384356 24460 384362 24472
rect 487154 24460 487160 24472
rect 384356 24432 487160 24460
rect 384356 24420 384362 24432
rect 487154 24420 487160 24432
rect 487212 24420 487218 24472
rect 316126 24352 316132 24404
rect 316184 24392 316190 24404
rect 422386 24392 422392 24404
rect 316184 24364 422392 24392
rect 316184 24352 316190 24364
rect 422386 24352 422392 24364
rect 422444 24352 422450 24404
rect 187326 24284 187332 24336
rect 187384 24324 187390 24336
rect 407206 24324 407212 24336
rect 187384 24296 407212 24324
rect 187384 24284 187390 24296
rect 407206 24284 407212 24296
rect 407264 24284 407270 24336
rect 148318 24216 148324 24268
rect 148376 24256 148382 24268
rect 247678 24256 247684 24268
rect 148376 24228 247684 24256
rect 148376 24216 148382 24228
rect 247678 24216 247684 24228
rect 247736 24216 247742 24268
rect 269758 24216 269764 24268
rect 269816 24256 269822 24268
rect 523126 24256 523132 24268
rect 269816 24228 523132 24256
rect 269816 24216 269822 24228
rect 523126 24216 523132 24228
rect 523184 24216 523190 24268
rect 184934 24148 184940 24200
rect 184992 24188 184998 24200
rect 452746 24188 452752 24200
rect 184992 24160 452752 24188
rect 184992 24148 184998 24160
rect 452746 24148 452752 24160
rect 452804 24148 452810 24200
rect 70302 24080 70308 24132
rect 70360 24120 70366 24132
rect 92474 24120 92480 24132
rect 70360 24092 92480 24120
rect 70360 24080 70366 24092
rect 92474 24080 92480 24092
rect 92532 24080 92538 24132
rect 93670 24080 93676 24132
rect 93728 24120 93734 24132
rect 104894 24120 104900 24132
rect 93728 24092 104900 24120
rect 93728 24080 93734 24092
rect 104894 24080 104900 24092
rect 104952 24080 104958 24132
rect 161198 24080 161204 24132
rect 161256 24120 161262 24132
rect 521654 24120 521660 24132
rect 161256 24092 521660 24120
rect 161256 24080 161262 24092
rect 521654 24080 521660 24092
rect 521712 24080 521718 24132
rect 402238 23060 402244 23112
rect 402296 23100 402302 23112
rect 408494 23100 408500 23112
rect 402296 23072 408500 23100
rect 402296 23060 402302 23072
rect 408494 23060 408500 23072
rect 408552 23060 408558 23112
rect 200022 22992 200028 23044
rect 200080 23032 200086 23044
rect 354674 23032 354680 23044
rect 200080 23004 354680 23032
rect 200080 22992 200086 23004
rect 354674 22992 354680 23004
rect 354732 22992 354738 23044
rect 389818 22992 389824 23044
rect 389876 23032 389882 23044
rect 462314 23032 462320 23044
rect 389876 23004 462320 23032
rect 389876 22992 389882 23004
rect 462314 22992 462320 23004
rect 462372 22992 462378 23044
rect 267826 22924 267832 22976
rect 267884 22964 267890 22976
rect 434898 22964 434904 22976
rect 267884 22936 434904 22964
rect 267884 22924 267890 22936
rect 434898 22924 434904 22936
rect 434956 22924 434962 22976
rect 252462 22856 252468 22908
rect 252520 22896 252526 22908
rect 576118 22896 576124 22908
rect 252520 22868 576124 22896
rect 252520 22856 252526 22868
rect 576118 22856 576124 22868
rect 576176 22856 576182 22908
rect 125594 22788 125600 22840
rect 125652 22828 125658 22840
rect 467834 22828 467840 22840
rect 125652 22800 467840 22828
rect 125652 22788 125658 22800
rect 467834 22788 467840 22800
rect 467892 22788 467898 22840
rect 71590 22720 71596 22772
rect 71648 22760 71654 22772
rect 85574 22760 85580 22772
rect 71648 22732 85580 22760
rect 71648 22720 71654 22732
rect 85574 22720 85580 22732
rect 85632 22720 85638 22772
rect 156966 22720 156972 22772
rect 157024 22760 157030 22772
rect 535454 22760 535460 22772
rect 157024 22732 535460 22760
rect 157024 22720 157030 22732
rect 535454 22720 535460 22732
rect 535512 22720 535518 22772
rect 95142 22516 95148 22568
rect 95200 22556 95206 22568
rect 97994 22556 98000 22568
rect 95200 22528 98000 22556
rect 95200 22516 95206 22528
rect 97994 22516 98000 22528
rect 98052 22516 98058 22568
rect 316678 22108 316684 22160
rect 316736 22148 316742 22160
rect 324406 22148 324412 22160
rect 316736 22120 324412 22148
rect 316736 22108 316742 22120
rect 324406 22108 324412 22120
rect 324464 22108 324470 22160
rect 299566 21700 299572 21752
rect 299624 21740 299630 21752
rect 321646 21740 321652 21752
rect 299624 21712 321652 21740
rect 299624 21700 299630 21712
rect 321646 21700 321652 21712
rect 321704 21700 321710 21752
rect 287698 21632 287704 21684
rect 287756 21672 287762 21684
rect 448606 21672 448612 21684
rect 287756 21644 448612 21672
rect 287756 21632 287762 21644
rect 448606 21632 448612 21644
rect 448664 21632 448670 21684
rect 188706 21564 188712 21616
rect 188764 21604 188770 21616
rect 397454 21604 397460 21616
rect 188764 21576 397460 21604
rect 188764 21564 188770 21576
rect 397454 21564 397460 21576
rect 397512 21564 397518 21616
rect 182082 21496 182088 21548
rect 182140 21536 182146 21548
rect 429194 21536 429200 21548
rect 182140 21508 429200 21536
rect 182140 21496 182146 21508
rect 429194 21496 429200 21508
rect 429252 21496 429258 21548
rect 86954 21428 86960 21480
rect 87012 21468 87018 21480
rect 97442 21468 97448 21480
rect 87012 21440 97448 21468
rect 87012 21428 87018 21440
rect 97442 21428 97448 21440
rect 97500 21428 97506 21480
rect 180702 21428 180708 21480
rect 180760 21468 180766 21480
rect 436094 21468 436100 21480
rect 180760 21440 436100 21468
rect 180760 21428 180766 21440
rect 436094 21428 436100 21440
rect 436152 21428 436158 21480
rect 9674 21360 9680 21412
rect 9732 21400 9738 21412
rect 87782 21400 87788 21412
rect 9732 21372 87788 21400
rect 9732 21360 9738 21372
rect 87782 21360 87788 21372
rect 87840 21360 87846 21412
rect 179322 21360 179328 21412
rect 179380 21400 179386 21412
rect 442994 21400 443000 21412
rect 179380 21372 443000 21400
rect 179380 21360 179386 21372
rect 442994 21360 443000 21372
rect 443052 21360 443058 21412
rect 398926 20612 398932 20664
rect 398984 20652 398990 20664
rect 404446 20652 404452 20664
rect 398984 20624 404452 20652
rect 398984 20612 398990 20624
rect 404446 20612 404452 20624
rect 404504 20612 404510 20664
rect 296714 20272 296720 20324
rect 296772 20312 296778 20324
rect 323118 20312 323124 20324
rect 296772 20284 323124 20312
rect 296772 20272 296778 20284
rect 323118 20272 323124 20284
rect 323176 20272 323182 20324
rect 340966 20272 340972 20324
rect 341024 20312 341030 20324
rect 416774 20312 416780 20324
rect 341024 20284 416780 20312
rect 341024 20272 341030 20284
rect 416774 20272 416780 20284
rect 416832 20272 416838 20324
rect 201126 20204 201132 20256
rect 201184 20244 201190 20256
rect 347774 20244 347780 20256
rect 201184 20216 347780 20244
rect 201184 20204 201190 20216
rect 347774 20204 347780 20216
rect 347832 20204 347838 20256
rect 194502 20136 194508 20188
rect 194560 20176 194566 20188
rect 375374 20176 375380 20188
rect 194560 20148 375380 20176
rect 194560 20136 194566 20148
rect 375374 20136 375380 20148
rect 375432 20136 375438 20188
rect 388438 20136 388444 20188
rect 388496 20176 388502 20188
rect 469214 20176 469220 20188
rect 388496 20148 469220 20176
rect 388496 20136 388502 20148
rect 469214 20136 469220 20148
rect 469272 20136 469278 20188
rect 192846 20068 192852 20120
rect 192904 20108 192910 20120
rect 382366 20108 382372 20120
rect 192904 20080 382372 20108
rect 192904 20068 192910 20080
rect 382366 20068 382372 20080
rect 382424 20068 382430 20120
rect 385678 20068 385684 20120
rect 385736 20108 385742 20120
rect 480254 20108 480260 20120
rect 385736 20080 480260 20108
rect 385736 20068 385742 20080
rect 480254 20068 480260 20080
rect 480312 20068 480318 20120
rect 282178 20000 282184 20052
rect 282236 20040 282242 20052
rect 473446 20040 473452 20052
rect 282236 20012 473452 20040
rect 282236 20000 282242 20012
rect 473446 20000 473452 20012
rect 473504 20000 473510 20052
rect 44174 19932 44180 19984
rect 44232 19972 44238 19984
rect 134518 19972 134524 19984
rect 44232 19944 134524 19972
rect 44232 19932 44238 19944
rect 134518 19932 134524 19944
rect 134576 19932 134582 19984
rect 191742 19932 191748 19984
rect 191800 19972 191806 19984
rect 390554 19972 390560 19984
rect 191800 19944 390560 19972
rect 191800 19932 191806 19944
rect 390554 19932 390560 19944
rect 390612 19932 390618 19984
rect 398098 19932 398104 19984
rect 398156 19972 398162 19984
rect 426434 19972 426440 19984
rect 398156 19944 426440 19972
rect 398156 19932 398162 19944
rect 426434 19932 426440 19944
rect 426492 19932 426498 19984
rect 155862 18912 155868 18964
rect 155920 18952 155926 18964
rect 542354 18952 542360 18964
rect 155920 18924 542360 18952
rect 155920 18912 155926 18924
rect 542354 18912 542360 18924
rect 542412 18912 542418 18964
rect 153010 18844 153016 18896
rect 153068 18884 153074 18896
rect 553394 18884 553400 18896
rect 153068 18856 553400 18884
rect 153068 18844 153074 18856
rect 553394 18844 553400 18856
rect 553452 18844 553458 18896
rect 152826 18776 152832 18828
rect 152884 18816 152890 18828
rect 556154 18816 556160 18828
rect 152884 18788 556160 18816
rect 152884 18776 152890 18788
rect 556154 18776 556160 18788
rect 556212 18776 556218 18828
rect 151722 18708 151728 18760
rect 151780 18748 151786 18760
rect 560294 18748 560300 18760
rect 151780 18720 560300 18748
rect 151780 18708 151786 18720
rect 560294 18708 560300 18720
rect 560352 18708 560358 18760
rect 148870 18640 148876 18692
rect 148928 18680 148934 18692
rect 571334 18680 571340 18692
rect 148928 18652 571340 18680
rect 148928 18640 148934 18652
rect 571334 18640 571340 18652
rect 571392 18640 571398 18692
rect 60734 18572 60740 18624
rect 60792 18612 60798 18624
rect 76742 18612 76748 18624
rect 60792 18584 76748 18612
rect 60792 18572 60798 18584
rect 76742 18572 76748 18584
rect 76800 18572 76806 18624
rect 80054 18572 80060 18624
rect 80112 18612 80118 18624
rect 98822 18612 98828 18624
rect 80112 18584 98828 18612
rect 80112 18572 80118 18584
rect 98822 18572 98828 18584
rect 98880 18572 98886 18624
rect 103514 18572 103520 18624
rect 103572 18612 103578 18624
rect 119522 18612 119528 18624
rect 103572 18584 119528 18612
rect 103572 18572 103578 18584
rect 119522 18572 119528 18584
rect 119580 18572 119586 18624
rect 148686 18572 148692 18624
rect 148744 18612 148750 18624
rect 574094 18612 574100 18624
rect 148744 18584 574100 18612
rect 148744 18572 148750 18584
rect 574094 18572 574100 18584
rect 574152 18572 574158 18624
rect 280798 17756 280804 17808
rect 280856 17796 280862 17808
rect 477494 17796 477500 17808
rect 280856 17768 477500 17796
rect 280856 17756 280862 17768
rect 477494 17756 477500 17768
rect 477552 17756 477558 17808
rect 169386 17688 169392 17740
rect 169444 17728 169450 17740
rect 481726 17728 481732 17740
rect 169444 17700 481732 17728
rect 169444 17688 169450 17700
rect 481726 17688 481732 17700
rect 481784 17688 481790 17740
rect 169570 17620 169576 17672
rect 169628 17660 169634 17672
rect 485774 17660 485780 17672
rect 169628 17632 485780 17660
rect 169628 17620 169634 17632
rect 485774 17620 485780 17632
rect 485832 17620 485838 17672
rect 168282 17552 168288 17604
rect 168340 17592 168346 17604
rect 490006 17592 490012 17604
rect 168340 17564 490012 17592
rect 168340 17552 168346 17564
rect 490006 17552 490012 17564
rect 490064 17552 490070 17604
rect 166626 17484 166632 17536
rect 166684 17524 166690 17536
rect 492674 17524 492680 17536
rect 166684 17496 492680 17524
rect 166684 17484 166690 17496
rect 492674 17484 492680 17496
rect 492732 17484 492738 17536
rect 166810 17416 166816 17468
rect 166868 17456 166874 17468
rect 496814 17456 496820 17468
rect 166868 17428 496820 17456
rect 166868 17416 166874 17428
rect 496814 17416 496820 17428
rect 496872 17416 496878 17468
rect 165246 17348 165252 17400
rect 165304 17388 165310 17400
rect 499574 17388 499580 17400
rect 165304 17360 499580 17388
rect 165304 17348 165310 17360
rect 499574 17348 499580 17360
rect 499632 17348 499638 17400
rect 100754 17280 100760 17332
rect 100812 17320 100818 17332
rect 120718 17320 120724 17332
rect 100812 17292 120724 17320
rect 100812 17280 100818 17292
rect 120718 17280 120724 17292
rect 120776 17280 120782 17332
rect 165430 17280 165436 17332
rect 165488 17320 165494 17332
rect 503714 17320 503720 17332
rect 165488 17292 503720 17320
rect 165488 17280 165494 17292
rect 503714 17280 503720 17292
rect 503772 17280 503778 17332
rect 66254 17212 66260 17264
rect 66312 17252 66318 17264
rect 101582 17252 101588 17264
rect 66312 17224 101588 17252
rect 66312 17212 66318 17224
rect 101582 17212 101588 17224
rect 101640 17212 101646 17264
rect 164142 17212 164148 17264
rect 164200 17252 164206 17264
rect 506566 17252 506572 17264
rect 164200 17224 506572 17252
rect 164200 17212 164206 17224
rect 506566 17212 506572 17224
rect 506624 17212 506630 17264
rect 295978 16260 295984 16312
rect 296036 16300 296042 16312
rect 414290 16300 414296 16312
rect 296036 16272 414296 16300
rect 296036 16260 296042 16272
rect 414290 16260 414296 16272
rect 414348 16260 414354 16312
rect 294782 16192 294788 16244
rect 294840 16232 294846 16244
rect 417418 16232 417424 16244
rect 294840 16204 417424 16232
rect 294840 16192 294846 16204
rect 417418 16192 417424 16204
rect 417476 16192 417482 16244
rect 294598 16124 294604 16176
rect 294656 16164 294662 16176
rect 420914 16164 420920 16176
rect 294656 16136 420920 16164
rect 294656 16124 294662 16136
rect 420914 16124 420920 16136
rect 420972 16124 420978 16176
rect 220446 16056 220452 16108
rect 220504 16096 220510 16108
rect 266538 16096 266544 16108
rect 220504 16068 266544 16096
rect 220504 16056 220510 16068
rect 266538 16056 266544 16068
rect 266596 16056 266602 16108
rect 293218 16056 293224 16108
rect 293276 16096 293282 16108
rect 423766 16096 423772 16108
rect 293276 16068 423772 16096
rect 293276 16056 293282 16068
rect 423766 16056 423772 16068
rect 423824 16056 423830 16108
rect 188522 15988 188528 16040
rect 188580 16028 188586 16040
rect 238202 16028 238208 16040
rect 188580 16000 238208 16028
rect 188580 15988 188586 16000
rect 238202 15988 238208 16000
rect 238260 15988 238266 16040
rect 292022 15988 292028 16040
rect 292080 16028 292086 16040
rect 428458 16028 428464 16040
rect 292080 16000 428464 16028
rect 292080 15988 292086 16000
rect 428458 15988 428464 16000
rect 428516 15988 428522 16040
rect 73338 15920 73344 15972
rect 73396 15960 73402 15972
rect 100018 15960 100024 15972
rect 73396 15932 100024 15960
rect 73396 15920 73402 15932
rect 100018 15920 100024 15932
rect 100076 15920 100082 15972
rect 177574 15920 177580 15972
rect 177632 15960 177638 15972
rect 239398 15960 239404 15972
rect 177632 15932 239404 15960
rect 177632 15920 177638 15932
rect 239398 15920 239404 15932
rect 239456 15920 239462 15972
rect 291838 15920 291844 15972
rect 291896 15960 291902 15972
rect 432046 15960 432052 15972
rect 291896 15932 432052 15960
rect 291896 15920 291902 15932
rect 432046 15920 432052 15932
rect 432104 15920 432110 15972
rect 93946 15852 93952 15904
rect 94004 15892 94010 15904
rect 122282 15892 122288 15904
rect 94004 15864 122288 15892
rect 94004 15852 94010 15864
rect 122282 15852 122288 15864
rect 122340 15852 122346 15904
rect 135254 15852 135260 15904
rect 135312 15892 135318 15904
rect 250622 15892 250628 15904
rect 135312 15864 250628 15892
rect 135312 15852 135318 15864
rect 250622 15852 250628 15864
rect 250680 15852 250686 15904
rect 289078 15852 289084 15904
rect 289136 15892 289142 15904
rect 442626 15892 442632 15904
rect 289136 15864 442632 15892
rect 289136 15852 289142 15864
rect 442626 15852 442632 15864
rect 442684 15852 442690 15904
rect 268378 14968 268384 15020
rect 268436 15008 268442 15020
rect 534442 15008 534448 15020
rect 268436 14980 534448 15008
rect 268436 14968 268442 14980
rect 534442 14968 534448 14980
rect 534500 14968 534506 15020
rect 266998 14900 267004 14952
rect 267056 14940 267062 14952
rect 538214 14940 538220 14952
rect 267056 14912 538220 14940
rect 267056 14900 267062 14912
rect 538214 14900 538220 14912
rect 538272 14900 538278 14952
rect 265618 14832 265624 14884
rect 265676 14872 265682 14884
rect 541986 14872 541992 14884
rect 265676 14844 541992 14872
rect 265676 14832 265682 14844
rect 541986 14832 541992 14844
rect 542044 14832 542050 14884
rect 260742 14764 260748 14816
rect 260800 14804 260806 14816
rect 545482 14804 545488 14816
rect 260800 14776 545488 14804
rect 260800 14764 260806 14776
rect 545482 14764 545488 14776
rect 545540 14764 545546 14816
rect 259086 14696 259092 14748
rect 259144 14736 259150 14748
rect 548426 14736 548432 14748
rect 259144 14708 548432 14736
rect 259144 14696 259150 14708
rect 548426 14696 548432 14708
rect 548484 14696 548490 14748
rect 259270 14628 259276 14680
rect 259328 14668 259334 14680
rect 552658 14668 552664 14680
rect 259328 14640 552664 14668
rect 259328 14628 259334 14640
rect 552658 14628 552664 14640
rect 552716 14628 552722 14680
rect 185026 14560 185032 14612
rect 185084 14600 185090 14612
rect 238018 14600 238024 14612
rect 185084 14572 238024 14600
rect 185084 14560 185090 14572
rect 238018 14560 238024 14572
rect 238076 14560 238082 14612
rect 257982 14560 257988 14612
rect 258040 14600 258046 14612
rect 556246 14600 556252 14612
rect 258040 14572 556252 14600
rect 258040 14560 258046 14572
rect 556246 14560 556252 14572
rect 556304 14560 556310 14612
rect 53282 14492 53288 14544
rect 53340 14532 53346 14544
rect 79318 14532 79324 14544
rect 53340 14504 79324 14532
rect 53340 14492 53346 14504
rect 79318 14492 79324 14504
rect 79376 14492 79382 14544
rect 151078 14492 151084 14544
rect 151136 14532 151142 14544
rect 246482 14532 246488 14544
rect 151136 14504 246488 14532
rect 151136 14492 151142 14504
rect 246482 14492 246488 14504
rect 246540 14492 246546 14544
rect 256510 14492 256516 14544
rect 256568 14532 256574 14544
rect 559282 14532 559288 14544
rect 256568 14504 559288 14532
rect 256568 14492 256574 14504
rect 559282 14492 559288 14504
rect 559340 14492 559346 14544
rect 79226 14424 79232 14476
rect 79284 14464 79290 14476
rect 126422 14464 126428 14476
rect 79284 14436 126428 14464
rect 79284 14424 79290 14436
rect 126422 14424 126428 14436
rect 126480 14424 126486 14476
rect 127526 14424 127532 14476
rect 127584 14464 127590 14476
rect 251818 14464 251824 14476
rect 127584 14436 251824 14464
rect 127584 14424 127590 14436
rect 251818 14424 251824 14436
rect 251876 14424 251882 14476
rect 256326 14424 256332 14476
rect 256384 14464 256390 14476
rect 563054 14464 563060 14476
rect 256384 14436 563060 14464
rect 256384 14424 256390 14436
rect 563054 14424 563060 14436
rect 563112 14424 563118 14476
rect 307018 13608 307024 13660
rect 307076 13648 307082 13660
rect 367738 13648 367744 13660
rect 307076 13620 367744 13648
rect 307076 13608 307082 13620
rect 367738 13608 367744 13620
rect 367796 13608 367802 13660
rect 305638 13540 305644 13592
rect 305696 13580 305702 13592
rect 371234 13580 371240 13592
rect 305696 13552 371240 13580
rect 305696 13540 305702 13552
rect 371234 13540 371240 13552
rect 371292 13540 371298 13592
rect 304442 13472 304448 13524
rect 304500 13512 304506 13524
rect 374086 13512 374092 13524
rect 304500 13484 374092 13512
rect 304500 13472 304506 13484
rect 374086 13472 374092 13484
rect 374144 13472 374150 13524
rect 304258 13404 304264 13456
rect 304316 13444 304322 13456
rect 378410 13444 378416 13456
rect 304316 13416 378416 13444
rect 304316 13404 304322 13416
rect 378410 13404 378416 13416
rect 378468 13404 378474 13456
rect 401042 13404 401048 13456
rect 401100 13444 401106 13456
rect 415486 13444 415492 13456
rect 401100 13416 415492 13444
rect 401100 13404 401106 13416
rect 415486 13404 415492 13416
rect 415544 13404 415550 13456
rect 302878 13336 302884 13388
rect 302936 13376 302942 13388
rect 385954 13376 385960 13388
rect 302936 13348 385960 13376
rect 302936 13336 302942 13348
rect 385954 13336 385960 13348
rect 386012 13336 386018 13388
rect 387794 13336 387800 13388
rect 387852 13376 387858 13388
rect 405918 13376 405924 13388
rect 387852 13348 405924 13376
rect 387852 13336 387858 13348
rect 405918 13336 405924 13348
rect 405976 13336 405982 13388
rect 301498 13268 301504 13320
rect 301556 13308 301562 13320
rect 389450 13308 389456 13320
rect 301556 13280 389456 13308
rect 301556 13268 301562 13280
rect 389450 13268 389456 13280
rect 389508 13268 389514 13320
rect 390646 13268 390652 13320
rect 390704 13308 390710 13320
rect 406102 13308 406108 13320
rect 390704 13280 406108 13308
rect 390704 13268 390710 13280
rect 406102 13268 406108 13280
rect 406160 13268 406166 13320
rect 64322 13200 64328 13252
rect 64380 13240 64386 13252
rect 76558 13240 76564 13252
rect 64380 13212 76564 13240
rect 64380 13200 64386 13212
rect 76558 13200 76564 13212
rect 76616 13200 76622 13252
rect 216858 13200 216864 13252
rect 216916 13240 216922 13252
rect 231118 13240 231124 13252
rect 216916 13212 231124 13240
rect 216916 13200 216922 13212
rect 231118 13200 231124 13212
rect 231176 13200 231182 13252
rect 300118 13200 300124 13252
rect 300176 13240 300182 13252
rect 392486 13240 392492 13252
rect 300176 13212 392492 13240
rect 300176 13200 300182 13212
rect 392486 13200 392492 13212
rect 392544 13200 392550 13252
rect 399478 13200 399484 13252
rect 399536 13240 399542 13252
rect 420178 13240 420184 13252
rect 399536 13212 420184 13240
rect 399536 13200 399542 13212
rect 420178 13200 420184 13212
rect 420236 13200 420242 13252
rect 68646 13132 68652 13184
rect 68704 13172 68710 13184
rect 95786 13172 95792 13184
rect 68704 13144 95792 13172
rect 68704 13132 68710 13144
rect 95786 13132 95792 13144
rect 95844 13132 95850 13184
rect 151814 13132 151820 13184
rect 151872 13172 151878 13184
rect 356054 13172 356060 13184
rect 151872 13144 356060 13172
rect 151872 13132 151878 13144
rect 356054 13132 356060 13144
rect 356112 13132 356118 13184
rect 384298 13132 384304 13184
rect 384356 13172 384362 13184
rect 407298 13172 407304 13184
rect 384356 13144 407304 13172
rect 384356 13132 384362 13144
rect 407298 13132 407304 13144
rect 407356 13132 407362 13184
rect 75914 13064 75920 13116
rect 75972 13104 75978 13116
rect 126238 13104 126244 13116
rect 75972 13076 126244 13104
rect 75972 13064 75978 13076
rect 126238 13064 126244 13076
rect 126296 13064 126302 13116
rect 147858 13064 147864 13116
rect 147916 13104 147922 13116
rect 357802 13104 357808 13116
rect 147916 13076 357808 13104
rect 147916 13064 147922 13076
rect 357802 13064 357808 13076
rect 357860 13064 357866 13116
rect 393958 13064 393964 13116
rect 394016 13104 394022 13116
rect 445018 13104 445024 13116
rect 394016 13076 445024 13104
rect 394016 13064 394022 13076
rect 445018 13064 445024 13076
rect 445076 13064 445082 13116
rect 312538 12180 312544 12232
rect 312596 12220 312602 12232
rect 339494 12220 339500 12232
rect 312596 12192 339500 12220
rect 312596 12180 312602 12192
rect 339494 12180 339500 12192
rect 339552 12180 339558 12232
rect 312722 12112 312728 12164
rect 312780 12152 312786 12164
rect 342254 12152 342260 12164
rect 312780 12124 342260 12152
rect 312780 12112 312786 12124
rect 342254 12112 342260 12124
rect 342312 12112 342318 12164
rect 311342 12044 311348 12096
rect 311400 12084 311406 12096
rect 346946 12084 346952 12096
rect 311400 12056 346952 12084
rect 311400 12044 311406 12056
rect 346946 12044 346952 12056
rect 347004 12044 347010 12096
rect 400858 12044 400864 12096
rect 400916 12084 400922 12096
rect 412634 12084 412640 12096
rect 400916 12056 412640 12084
rect 400916 12044 400922 12056
rect 412634 12044 412640 12056
rect 412692 12044 412698 12096
rect 211062 11976 211068 12028
rect 211120 12016 211126 12028
rect 305546 12016 305552 12028
rect 211120 11988 305552 12016
rect 211120 11976 211126 11988
rect 305546 11976 305552 11988
rect 305604 11976 305610 12028
rect 311158 11976 311164 12028
rect 311216 12016 311222 12028
rect 349246 12016 349252 12028
rect 311216 11988 349252 12016
rect 311216 11976 311222 11988
rect 349246 11976 349252 11988
rect 349304 11976 349310 12028
rect 396718 11976 396724 12028
rect 396776 12016 396782 12028
rect 430850 12016 430856 12028
rect 396776 11988 430856 12016
rect 396776 11976 396782 11988
rect 430850 11976 430856 11988
rect 430908 11976 430914 12028
rect 153010 11908 153016 11960
rect 153068 11948 153074 11960
rect 246298 11948 246304 11960
rect 153068 11920 246304 11948
rect 153068 11908 153074 11920
rect 246298 11908 246304 11920
rect 246356 11908 246362 11960
rect 309778 11908 309784 11960
rect 309836 11948 309842 11960
rect 353570 11948 353576 11960
rect 309836 11920 353576 11948
rect 309836 11908 309842 11920
rect 353570 11908 353576 11920
rect 353628 11908 353634 11960
rect 365806 11908 365812 11960
rect 365864 11948 365870 11960
rect 411346 11948 411352 11960
rect 365864 11920 411352 11948
rect 365864 11908 365870 11920
rect 411346 11908 411352 11920
rect 411404 11908 411410 11960
rect 209406 11840 209412 11892
rect 209464 11880 209470 11892
rect 312170 11880 312176 11892
rect 209464 11852 312176 11880
rect 209464 11840 209470 11852
rect 312170 11840 312176 11852
rect 312228 11840 312234 11892
rect 313918 11840 313924 11892
rect 313976 11880 313982 11892
rect 335446 11880 335452 11892
rect 313976 11852 335452 11880
rect 313976 11840 313982 11852
rect 335446 11840 335452 11852
rect 335504 11840 335510 11892
rect 338666 11840 338672 11892
rect 338724 11880 338730 11892
rect 418246 11880 418252 11892
rect 338724 11852 418252 11880
rect 338724 11840 338730 11852
rect 418246 11840 418252 11852
rect 418304 11840 418310 11892
rect 144454 11772 144460 11824
rect 144512 11812 144518 11824
rect 357618 11812 357624 11824
rect 144512 11784 357624 11812
rect 144512 11772 144518 11784
rect 357618 11772 357624 11784
rect 357676 11772 357682 11824
rect 392578 11772 392584 11824
rect 392636 11812 392642 11824
rect 451642 11812 451648 11824
rect 392636 11784 451648 11812
rect 392636 11772 392642 11784
rect 451642 11772 451648 11784
rect 451700 11772 451706 11824
rect 65058 11704 65064 11756
rect 65116 11744 65122 11756
rect 128998 11744 129004 11756
rect 65116 11716 129004 11744
rect 65116 11704 65122 11716
rect 128998 11704 129004 11716
rect 129056 11704 129062 11756
rect 168374 11704 168380 11756
rect 168432 11744 168438 11756
rect 169570 11744 169576 11756
rect 168432 11716 169576 11744
rect 168432 11704 168438 11716
rect 169570 11704 169576 11716
rect 169628 11704 169634 11756
rect 184934 11704 184940 11756
rect 184992 11744 184998 11756
rect 186130 11744 186136 11756
rect 184992 11716 186136 11744
rect 184992 11704 184998 11716
rect 186130 11704 186136 11716
rect 186188 11704 186194 11756
rect 425698 11744 425704 11756
rect 190426 11716 425704 11744
rect 183186 11636 183192 11688
rect 183244 11676 183250 11688
rect 190426 11676 190454 11716
rect 425698 11704 425704 11716
rect 425756 11704 425762 11756
rect 183244 11648 190454 11676
rect 183244 11636 183250 11648
rect 259454 11636 259460 11688
rect 259512 11676 259518 11688
rect 260650 11676 260656 11688
rect 259512 11648 260656 11676
rect 259512 11636 259518 11648
rect 260650 11636 260656 11648
rect 260708 11636 260714 11688
rect 91554 11024 91560 11076
rect 91612 11064 91618 11076
rect 95878 11064 95884 11076
rect 91612 11036 95884 11064
rect 91612 11024 91618 11036
rect 95878 11024 95884 11036
rect 95936 11024 95942 11076
rect 217686 10684 217692 10736
rect 217744 10724 217750 10736
rect 276658 10724 276664 10736
rect 217744 10696 276664 10724
rect 217744 10684 217750 10696
rect 276658 10684 276664 10696
rect 276716 10684 276722 10736
rect 216306 10616 216312 10668
rect 216364 10656 216370 10668
rect 280706 10656 280712 10668
rect 216364 10628 280712 10656
rect 216364 10616 216370 10628
rect 280706 10616 280712 10628
rect 280764 10616 280770 10668
rect 286594 10616 286600 10668
rect 286652 10656 286658 10668
rect 324774 10656 324780 10668
rect 286652 10628 324780 10656
rect 286652 10616 286658 10628
rect 324774 10616 324780 10628
rect 324832 10616 324838 10668
rect 370130 10616 370136 10668
rect 370188 10656 370194 10668
rect 409966 10656 409972 10668
rect 370188 10628 409972 10656
rect 370188 10616 370194 10628
rect 409966 10616 409972 10628
rect 410024 10616 410030 10668
rect 215202 10548 215208 10600
rect 215260 10588 215266 10600
rect 287330 10588 287336 10600
rect 215260 10560 287336 10588
rect 215260 10548 215266 10560
rect 287330 10548 287336 10560
rect 287388 10548 287394 10600
rect 289814 10548 289820 10600
rect 289872 10588 289878 10600
rect 324590 10588 324596 10600
rect 289872 10560 324596 10588
rect 289872 10548 289878 10560
rect 324590 10548 324596 10560
rect 324648 10548 324654 10600
rect 363506 10548 363512 10600
rect 363564 10588 363570 10600
rect 412910 10588 412916 10600
rect 363564 10560 412916 10588
rect 363564 10548 363570 10560
rect 412910 10548 412916 10560
rect 412968 10548 412974 10600
rect 213546 10480 213552 10532
rect 213604 10520 213610 10532
rect 291378 10520 291384 10532
rect 213604 10492 291384 10520
rect 213604 10480 213610 10492
rect 291378 10480 291384 10492
rect 291436 10480 291442 10532
rect 293218 10480 293224 10532
rect 293276 10520 293282 10532
rect 323302 10520 323308 10532
rect 293276 10492 323308 10520
rect 293276 10480 293282 10492
rect 323302 10480 323308 10492
rect 323360 10480 323366 10532
rect 359458 10480 359464 10532
rect 359516 10520 359522 10532
rect 412726 10520 412732 10532
rect 359516 10492 412732 10520
rect 359516 10480 359522 10492
rect 412726 10480 412732 10492
rect 412784 10480 412790 10532
rect 213730 10412 213736 10464
rect 213788 10452 213794 10464
rect 294874 10452 294880 10464
rect 213788 10424 294880 10452
rect 213788 10412 213794 10424
rect 294874 10412 294880 10424
rect 294932 10412 294938 10464
rect 314654 10412 314660 10464
rect 314712 10452 314718 10464
rect 318886 10452 318892 10464
rect 314712 10424 318892 10452
rect 314712 10412 314718 10424
rect 318886 10412 318892 10424
rect 318944 10412 318950 10464
rect 356330 10412 356336 10464
rect 356388 10452 356394 10464
rect 414014 10452 414020 10464
rect 356388 10424 414020 10452
rect 356388 10412 356394 10424
rect 414014 10412 414020 10424
rect 414072 10412 414078 10464
rect 72970 10344 72976 10396
rect 73028 10384 73034 10396
rect 81618 10384 81624 10396
rect 73028 10356 81624 10384
rect 73028 10344 73034 10356
rect 81618 10344 81624 10356
rect 81676 10344 81682 10396
rect 84194 10344 84200 10396
rect 84252 10384 84258 10396
rect 97258 10384 97264 10396
rect 84252 10356 97264 10384
rect 84252 10344 84258 10356
rect 97258 10344 97264 10356
rect 97316 10344 97322 10396
rect 212166 10344 212172 10396
rect 212224 10384 212230 10396
rect 298094 10384 298100 10396
rect 212224 10356 298100 10384
rect 212224 10344 212230 10356
rect 298094 10344 298100 10356
rect 298152 10344 298158 10396
rect 307938 10344 307944 10396
rect 307996 10384 308002 10396
rect 320542 10384 320548 10396
rect 307996 10356 320548 10384
rect 307996 10344 308002 10356
rect 320542 10344 320548 10356
rect 320600 10344 320606 10396
rect 352834 10344 352840 10396
rect 352892 10384 352898 10396
rect 414106 10384 414112 10396
rect 352892 10356 414112 10384
rect 352892 10344 352898 10356
rect 414106 10344 414112 10356
rect 414164 10344 414170 10396
rect 47394 10276 47400 10328
rect 47452 10316 47458 10328
rect 133138 10316 133144 10328
rect 47452 10288 133144 10316
rect 47452 10276 47458 10288
rect 133138 10276 133144 10288
rect 133196 10276 133202 10328
rect 212350 10276 212356 10328
rect 212408 10316 212414 10328
rect 301498 10316 301504 10328
rect 212408 10288 301504 10316
rect 212408 10276 212414 10288
rect 301498 10276 301504 10288
rect 301556 10276 301562 10328
rect 303890 10276 303896 10328
rect 303948 10316 303954 10328
rect 320358 10316 320364 10328
rect 303948 10288 320364 10316
rect 303948 10276 303954 10288
rect 320358 10276 320364 10288
rect 320416 10276 320422 10328
rect 345014 10276 345020 10328
rect 345072 10316 345078 10328
rect 416958 10316 416964 10328
rect 345072 10288 416964 10316
rect 345072 10276 345078 10288
rect 416958 10276 416964 10288
rect 417016 10276 417022 10328
rect 310238 9324 310244 9376
rect 310296 9364 310302 9376
rect 425146 9364 425152 9376
rect 310296 9336 425152 9364
rect 310296 9324 310302 9336
rect 425146 9324 425152 9336
rect 425204 9324 425210 9376
rect 306742 9256 306748 9308
rect 306800 9296 306806 9308
rect 425330 9296 425336 9308
rect 306800 9268 425336 9296
rect 306800 9256 306806 9268
rect 425330 9256 425336 9268
rect 425388 9256 425394 9308
rect 227622 9188 227628 9240
rect 227680 9228 227686 9240
rect 234614 9228 234620 9240
rect 227680 9200 234620 9228
rect 227680 9188 227686 9200
rect 234614 9188 234620 9200
rect 234672 9188 234678 9240
rect 296070 9188 296076 9240
rect 296128 9228 296134 9240
rect 427906 9228 427912 9240
rect 296128 9200 427912 9228
rect 296128 9188 296134 9200
rect 427906 9188 427912 9200
rect 427964 9188 427970 9240
rect 224770 9120 224776 9172
rect 224828 9160 224834 9172
rect 245194 9160 245200 9172
rect 224828 9132 245200 9160
rect 224828 9120 224834 9132
rect 245194 9120 245200 9132
rect 245252 9120 245258 9172
rect 292574 9120 292580 9172
rect 292632 9160 292638 9172
rect 429562 9160 429568 9172
rect 292632 9132 429568 9160
rect 292632 9120 292638 9132
rect 429562 9120 429568 9132
rect 429620 9120 429626 9172
rect 77386 9052 77392 9104
rect 77444 9092 77450 9104
rect 77444 9064 84194 9092
rect 77444 9052 77450 9064
rect 72786 8984 72792 9036
rect 72844 9024 72850 9036
rect 78582 9024 78588 9036
rect 72844 8996 78588 9024
rect 72844 8984 72850 8996
rect 78582 8984 78588 8996
rect 78640 8984 78646 9036
rect 84166 9024 84194 9064
rect 93762 9052 93768 9104
rect 93820 9092 93826 9104
rect 102226 9092 102232 9104
rect 93820 9064 102232 9092
rect 93820 9052 93826 9064
rect 102226 9052 102232 9064
rect 102284 9052 102290 9104
rect 224862 9052 224868 9104
rect 224920 9092 224926 9104
rect 248782 9092 248788 9104
rect 224920 9064 248788 9092
rect 224920 9052 224926 9064
rect 248782 9052 248788 9064
rect 248840 9052 248846 9104
rect 288986 9052 288992 9104
rect 289044 9092 289050 9104
rect 429378 9092 429384 9104
rect 289044 9064 429384 9092
rect 289044 9052 289050 9064
rect 429378 9052 429384 9064
rect 429436 9052 429442 9104
rect 98638 9024 98644 9036
rect 84166 8996 98644 9024
rect 98638 8984 98644 8996
rect 98696 8984 98702 9036
rect 223482 8984 223488 9036
rect 223540 9024 223546 9036
rect 252370 9024 252376 9036
rect 223540 8996 252376 9024
rect 223540 8984 223546 8996
rect 252370 8984 252376 8996
rect 252428 8984 252434 9036
rect 285398 8984 285404 9036
rect 285456 9024 285462 9036
rect 430666 9024 430672 9036
rect 285456 8996 430672 9024
rect 285456 8984 285462 8996
rect 430666 8984 430672 8996
rect 430724 8984 430730 9036
rect 62022 8916 62028 8968
rect 62080 8956 62086 8968
rect 130378 8956 130384 8968
rect 62080 8928 130384 8956
rect 62080 8916 62086 8928
rect 130378 8916 130384 8928
rect 130436 8916 130442 8968
rect 131758 8916 131764 8968
rect 131816 8956 131822 8968
rect 250438 8956 250444 8968
rect 131816 8928 250444 8956
rect 131816 8916 131822 8928
rect 250438 8916 250444 8928
rect 250496 8916 250502 8968
rect 281902 8916 281908 8968
rect 281960 8956 281966 8968
rect 430574 8956 430580 8968
rect 281960 8928 430580 8956
rect 281960 8916 281966 8928
rect 430574 8916 430580 8928
rect 430632 8916 430638 8968
rect 223942 8372 223948 8424
rect 224000 8412 224006 8424
rect 229922 8412 229928 8424
rect 224000 8384 229928 8412
rect 224000 8372 224006 8384
rect 229922 8372 229928 8384
rect 229980 8372 229986 8424
rect 229002 8304 229008 8356
rect 229060 8344 229066 8356
rect 231026 8344 231032 8356
rect 229060 8316 231032 8344
rect 229060 8304 229066 8316
rect 231026 8304 231032 8316
rect 231084 8304 231090 8356
rect 227530 8168 227536 8220
rect 227588 8208 227594 8220
rect 228358 8208 228364 8220
rect 227588 8180 228364 8208
rect 227588 8168 227594 8180
rect 228358 8168 228364 8180
rect 228416 8168 228422 8220
rect 92382 7964 92388 8016
rect 92440 8004 92446 8016
rect 109310 8004 109316 8016
rect 92440 7976 109316 8004
rect 92440 7964 92446 7976
rect 109310 7964 109316 7976
rect 109368 7964 109374 8016
rect 249978 7964 249984 8016
rect 250036 8004 250042 8016
rect 439222 8004 439228 8016
rect 250036 7976 439228 8004
rect 250036 7964 250042 7976
rect 439222 7964 439228 7976
rect 439280 7964 439286 8016
rect 90726 7896 90732 7948
rect 90784 7936 90790 7948
rect 116394 7936 116400 7948
rect 90784 7908 116400 7936
rect 90784 7896 90790 7908
rect 116394 7896 116400 7908
rect 116452 7896 116458 7948
rect 170766 7896 170772 7948
rect 170824 7936 170830 7948
rect 242342 7936 242348 7948
rect 170824 7908 242348 7936
rect 170824 7896 170830 7908
rect 242342 7896 242348 7908
rect 242400 7896 242406 7948
rect 246390 7896 246396 7948
rect 246448 7936 246454 7948
rect 439038 7936 439044 7948
rect 246448 7908 439044 7936
rect 246448 7896 246454 7908
rect 439038 7896 439044 7908
rect 439096 7896 439102 7948
rect 89530 7828 89536 7880
rect 89588 7868 89594 7880
rect 119890 7868 119896 7880
rect 89588 7840 119896 7868
rect 89588 7828 89594 7840
rect 119890 7828 119896 7840
rect 119948 7828 119954 7880
rect 195606 7828 195612 7880
rect 195664 7868 195670 7880
rect 235258 7868 235264 7880
rect 195664 7840 235264 7868
rect 195664 7828 195670 7840
rect 235258 7828 235264 7840
rect 235316 7828 235322 7880
rect 239306 7828 239312 7880
rect 239364 7868 239370 7880
rect 440418 7868 440424 7880
rect 239364 7840 440424 7868
rect 239364 7828 239370 7840
rect 440418 7828 440424 7840
rect 440476 7828 440482 7880
rect 45462 7760 45468 7812
rect 45520 7800 45526 7812
rect 106918 7800 106924 7812
rect 45520 7772 106924 7800
rect 45520 7760 45526 7772
rect 106918 7760 106924 7772
rect 106976 7760 106982 7812
rect 209866 7760 209872 7812
rect 209924 7800 209930 7812
rect 232498 7800 232504 7812
rect 209924 7772 232504 7800
rect 209924 7760 209930 7772
rect 232498 7760 232504 7772
rect 232556 7760 232562 7812
rect 235810 7760 235816 7812
rect 235868 7800 235874 7812
rect 441706 7800 441712 7812
rect 235868 7772 441712 7800
rect 235868 7760 235874 7772
rect 441706 7760 441712 7772
rect 441764 7760 441770 7812
rect 38378 7692 38384 7744
rect 38436 7732 38442 7744
rect 108298 7732 108304 7744
rect 38436 7704 108304 7732
rect 38436 7692 38442 7704
rect 108298 7692 108304 7704
rect 108356 7692 108362 7744
rect 232222 7692 232228 7744
rect 232280 7732 232286 7744
rect 443178 7732 443184 7744
rect 232280 7704 443184 7732
rect 232280 7692 232286 7704
rect 443178 7692 443184 7704
rect 443236 7692 443242 7744
rect 31294 7624 31300 7676
rect 31352 7664 31358 7676
rect 109678 7664 109684 7676
rect 31352 7636 109684 7664
rect 31352 7624 31358 7636
rect 109678 7624 109684 7636
rect 109736 7624 109742 7676
rect 228726 7624 228732 7676
rect 228784 7664 228790 7676
rect 443362 7664 443368 7676
rect 228784 7636 443368 7664
rect 228784 7624 228790 7636
rect 443362 7624 443368 7636
rect 443420 7624 443426 7676
rect 23014 7556 23020 7608
rect 23072 7596 23078 7608
rect 111058 7596 111064 7608
rect 23072 7568 111064 7596
rect 23072 7556 23078 7568
rect 111058 7556 111064 7568
rect 111116 7556 111122 7608
rect 132954 7556 132960 7608
rect 133012 7596 133018 7608
rect 465350 7596 465356 7608
rect 133012 7568 465356 7596
rect 133012 7556 133018 7568
rect 465350 7556 465356 7568
rect 465408 7556 465414 7608
rect 93854 7488 93860 7540
rect 93912 7528 93918 7540
rect 94774 7528 94780 7540
rect 93912 7500 94780 7528
rect 93912 7488 93918 7500
rect 94774 7488 94780 7500
rect 94832 7488 94838 7540
rect 220446 6740 220452 6792
rect 220504 6780 220510 6792
rect 229738 6780 229744 6792
rect 220504 6752 229744 6780
rect 220504 6740 220510 6752
rect 229738 6740 229744 6752
rect 229796 6740 229802 6792
rect 202690 6672 202696 6724
rect 202748 6712 202754 6724
rect 233878 6712 233884 6724
rect 202748 6684 233884 6712
rect 202748 6672 202754 6684
rect 233878 6672 233884 6684
rect 233936 6672 233942 6724
rect 174262 6604 174268 6656
rect 174320 6644 174326 6656
rect 240778 6644 240784 6656
rect 174320 6616 240784 6644
rect 174320 6604 174326 6616
rect 240778 6604 240784 6616
rect 240836 6604 240842 6656
rect 167178 6536 167184 6588
rect 167236 6576 167242 6588
rect 242158 6576 242164 6588
rect 167236 6548 242164 6576
rect 167236 6536 167242 6548
rect 242158 6536 242164 6548
rect 242216 6536 242222 6588
rect 247586 6536 247592 6588
rect 247644 6576 247650 6588
rect 334066 6576 334072 6588
rect 247644 6548 334072 6576
rect 247644 6536 247650 6548
rect 334066 6536 334072 6548
rect 334124 6536 334130 6588
rect 70302 6468 70308 6520
rect 70360 6508 70366 6520
rect 101398 6508 101404 6520
rect 70360 6480 101404 6508
rect 70360 6468 70366 6480
rect 101398 6468 101404 6480
rect 101456 6468 101462 6520
rect 192018 6468 192024 6520
rect 192076 6508 192082 6520
rect 236638 6508 236644 6520
rect 192076 6480 236644 6508
rect 192076 6468 192082 6480
rect 236638 6468 236644 6480
rect 236696 6468 236702 6520
rect 240502 6468 240508 6520
rect 240560 6508 240566 6520
rect 335538 6508 335544 6520
rect 240560 6480 335544 6508
rect 240560 6468 240566 6480
rect 335538 6468 335544 6480
rect 335596 6468 335602 6520
rect 63218 6400 63224 6452
rect 63276 6440 63282 6452
rect 102962 6440 102968 6452
rect 63276 6412 102968 6440
rect 63276 6400 63282 6412
rect 102962 6400 102968 6412
rect 103020 6400 103026 6452
rect 229830 6400 229836 6452
rect 229888 6440 229894 6452
rect 338206 6440 338212 6452
rect 229888 6412 338212 6440
rect 229888 6400 229894 6412
rect 338206 6400 338212 6412
rect 338264 6400 338270 6452
rect 59630 6332 59636 6384
rect 59688 6372 59694 6384
rect 102778 6372 102784 6384
rect 59688 6344 102784 6372
rect 59688 6332 59694 6344
rect 102778 6332 102784 6344
rect 102836 6332 102842 6384
rect 226334 6332 226340 6384
rect 226392 6372 226398 6384
rect 338114 6372 338120 6384
rect 226392 6344 338120 6372
rect 226392 6332 226398 6344
rect 338114 6332 338120 6344
rect 338172 6332 338178 6384
rect 56042 6264 56048 6316
rect 56100 6304 56106 6316
rect 104158 6304 104164 6316
rect 56100 6276 104164 6304
rect 56100 6264 56106 6276
rect 104158 6264 104164 6276
rect 104216 6264 104222 6316
rect 222746 6264 222752 6316
rect 222804 6304 222810 6316
rect 339586 6304 339592 6316
rect 222804 6276 339592 6304
rect 222804 6264 222810 6276
rect 339586 6264 339592 6276
rect 339644 6264 339650 6316
rect 364978 6264 364984 6316
rect 365036 6304 365042 6316
rect 569126 6304 569132 6316
rect 365036 6276 569132 6304
rect 365036 6264 365042 6276
rect 569126 6264 569132 6276
rect 569184 6264 569190 6316
rect 52546 6196 52552 6248
rect 52604 6236 52610 6248
rect 105814 6236 105820 6248
rect 52604 6208 105820 6236
rect 52604 6196 52610 6208
rect 105814 6196 105820 6208
rect 105872 6196 105878 6248
rect 219250 6196 219256 6248
rect 219308 6236 219314 6248
rect 341150 6236 341156 6248
rect 219308 6208 341156 6236
rect 219308 6196 219314 6208
rect 341150 6196 341156 6208
rect 341208 6196 341214 6248
rect 363782 6196 363788 6248
rect 363840 6236 363846 6248
rect 572714 6236 572720 6248
rect 363840 6208 572720 6236
rect 363840 6196 363846 6208
rect 572714 6196 572720 6208
rect 572772 6196 572778 6248
rect 48958 6128 48964 6180
rect 49016 6168 49022 6180
rect 105538 6168 105544 6180
rect 49016 6140 105544 6168
rect 49016 6128 49022 6140
rect 105538 6128 105544 6140
rect 105596 6128 105602 6180
rect 108114 6128 108120 6180
rect 108172 6168 108178 6180
rect 119338 6168 119344 6180
rect 108172 6140 119344 6168
rect 108172 6128 108178 6140
rect 119338 6128 119344 6140
rect 119396 6128 119402 6180
rect 134150 6128 134156 6180
rect 134208 6168 134214 6180
rect 360286 6168 360292 6180
rect 134208 6140 360292 6168
rect 134208 6128 134214 6140
rect 360286 6128 360292 6140
rect 360344 6128 360350 6180
rect 363598 6128 363604 6180
rect 363656 6168 363662 6180
rect 576302 6168 576308 6180
rect 363656 6140 576308 6168
rect 363656 6128 363662 6140
rect 576302 6128 576308 6140
rect 576360 6128 576366 6180
rect 403066 5856 403072 5908
rect 403124 5856 403130 5908
rect 402974 5652 402980 5704
rect 403032 5692 403038 5704
rect 403084 5692 403112 5856
rect 403032 5664 403112 5692
rect 403032 5652 403038 5664
rect 340138 5312 340144 5364
rect 340196 5352 340202 5364
rect 346394 5352 346400 5364
rect 340196 5324 346400 5352
rect 340196 5312 340202 5324
rect 346394 5312 346400 5324
rect 346452 5312 346458 5364
rect 212166 5244 212172 5296
rect 212224 5284 212230 5296
rect 342346 5284 342352 5296
rect 212224 5256 342352 5284
rect 212224 5244 212230 5256
rect 342346 5244 342352 5256
rect 342404 5244 342410 5296
rect 71406 5176 71412 5228
rect 71464 5216 71470 5228
rect 89162 5216 89168 5228
rect 71464 5188 89168 5216
rect 71464 5176 71470 5188
rect 89162 5176 89168 5188
rect 89220 5176 89226 5228
rect 97442 5176 97448 5228
rect 97500 5216 97506 5228
rect 122098 5216 122104 5228
rect 97500 5188 122104 5216
rect 97500 5176 97506 5188
rect 122098 5176 122104 5188
rect 122156 5176 122162 5228
rect 208578 5176 208584 5228
rect 208636 5216 208642 5228
rect 342530 5216 342536 5228
rect 208636 5188 342536 5216
rect 208636 5176 208642 5188
rect 342530 5176 342536 5188
rect 342588 5176 342594 5228
rect 72602 5108 72608 5160
rect 72660 5148 72666 5160
rect 72660 5120 79456 5148
rect 72660 5108 72666 5120
rect 69106 5040 69112 5092
rect 69164 5080 69170 5092
rect 69164 5052 79180 5080
rect 69164 5040 69170 5052
rect 71498 4904 71504 4956
rect 71556 4944 71562 4956
rect 75178 4944 75184 4956
rect 71556 4916 75184 4944
rect 71556 4904 71562 4916
rect 75178 4904 75184 4916
rect 75236 4904 75242 4956
rect 79152 4944 79180 5052
rect 79428 5012 79456 5120
rect 86862 5108 86868 5160
rect 86920 5148 86926 5160
rect 123478 5148 123484 5160
rect 86920 5120 123484 5148
rect 86920 5108 86926 5120
rect 123478 5108 123484 5120
rect 123536 5108 123542 5160
rect 201494 5108 201500 5160
rect 201552 5148 201558 5160
rect 345106 5148 345112 5160
rect 201552 5120 345112 5148
rect 201552 5108 201558 5120
rect 345106 5108 345112 5120
rect 345164 5108 345170 5160
rect 83274 5040 83280 5092
rect 83332 5080 83338 5092
rect 124858 5080 124864 5092
rect 83332 5052 124864 5080
rect 83332 5040 83338 5052
rect 124858 5040 124864 5052
rect 124916 5040 124922 5092
rect 197906 5040 197912 5092
rect 197964 5080 197970 5092
rect 345382 5080 345388 5092
rect 197964 5052 345388 5080
rect 197964 5040 197970 5052
rect 345382 5040 345388 5052
rect 345440 5040 345446 5092
rect 378778 5040 378784 5092
rect 378836 5080 378842 5092
rect 508866 5080 508872 5092
rect 378836 5052 508872 5080
rect 378836 5040 378842 5052
rect 508866 5040 508872 5052
rect 508924 5040 508930 5092
rect 127802 5012 127808 5024
rect 79428 4984 127808 5012
rect 127802 4972 127808 4984
rect 127860 4972 127866 5024
rect 194410 4972 194416 5024
rect 194468 5012 194474 5024
rect 346486 5012 346492 5024
rect 194468 4984 346492 5012
rect 194468 4972 194474 4984
rect 346486 4972 346492 4984
rect 346544 4972 346550 5024
rect 378962 4972 378968 5024
rect 379020 5012 379026 5024
rect 512454 5012 512460 5024
rect 379020 4984 512460 5012
rect 379020 4972 379026 4984
rect 512454 4972 512460 4984
rect 512512 4972 512518 5024
rect 127618 4944 127624 4956
rect 79152 4916 127624 4944
rect 127618 4904 127624 4916
rect 127676 4904 127682 4956
rect 190822 4904 190828 4956
rect 190880 4944 190886 4956
rect 340138 4944 340144 4956
rect 190880 4916 340144 4944
rect 190880 4904 190886 4916
rect 340138 4904 340144 4916
rect 340196 4904 340202 4956
rect 377398 4904 377404 4956
rect 377456 4944 377462 4956
rect 515950 4944 515956 4956
rect 377456 4916 515956 4944
rect 377456 4904 377462 4916
rect 515950 4904 515956 4916
rect 516008 4904 516014 4956
rect 14734 4836 14740 4888
rect 14792 4876 14798 4888
rect 87598 4876 87604 4888
rect 14792 4848 87604 4876
rect 14792 4836 14798 4848
rect 87598 4836 87604 4848
rect 87656 4836 87662 4888
rect 90358 4836 90364 4888
rect 90416 4876 90422 4888
rect 123662 4876 123668 4888
rect 90416 4848 123668 4876
rect 90416 4836 90422 4848
rect 123662 4836 123668 4848
rect 123720 4836 123726 4888
rect 187326 4836 187332 4888
rect 187384 4876 187390 4888
rect 347866 4876 347872 4888
rect 187384 4848 347872 4876
rect 187384 4836 187390 4848
rect 347866 4836 347872 4848
rect 347924 4836 347930 4888
rect 376110 4836 376116 4888
rect 376168 4876 376174 4888
rect 519538 4876 519544 4888
rect 376168 4848 519544 4876
rect 376168 4836 376174 4848
rect 519538 4836 519544 4848
rect 519596 4836 519602 4888
rect 12342 4768 12348 4820
rect 12400 4808 12406 4820
rect 140038 4808 140044 4820
rect 12400 4780 140044 4808
rect 12400 4768 12406 4780
rect 140038 4768 140044 4780
rect 140096 4768 140102 4820
rect 183738 4768 183744 4820
rect 183796 4808 183802 4820
rect 349430 4808 349436 4820
rect 183796 4780 349436 4808
rect 183796 4768 183802 4780
rect 349430 4768 349436 4780
rect 349488 4768 349494 4820
rect 371878 4768 371884 4820
rect 371936 4808 371942 4820
rect 537202 4808 537208 4820
rect 371936 4780 537208 4808
rect 371936 4768 371942 4780
rect 537202 4768 537208 4780
rect 537260 4768 537266 4820
rect 74442 4632 74448 4684
rect 74500 4672 74506 4684
rect 74994 4672 75000 4684
rect 74500 4644 75000 4672
rect 74500 4632 74506 4644
rect 74994 4632 75000 4644
rect 75052 4632 75058 4684
rect 67910 4428 67916 4480
rect 67968 4468 67974 4480
rect 75362 4468 75368 4480
rect 67968 4440 75368 4468
rect 67968 4428 67974 4440
rect 75362 4428 75368 4440
rect 75420 4428 75426 4480
rect 209774 4156 209780 4208
rect 209832 4196 209838 4208
rect 210970 4196 210976 4208
rect 209832 4168 210976 4196
rect 209832 4156 209838 4168
rect 210970 4156 210976 4168
rect 211028 4156 211034 4208
rect 267734 4156 267740 4208
rect 267792 4196 267798 4208
rect 268470 4196 268476 4208
rect 267792 4168 268476 4196
rect 267792 4156 267798 4168
rect 268470 4156 268476 4168
rect 268528 4156 268534 4208
rect 299566 4156 299572 4208
rect 299624 4196 299630 4208
rect 300762 4196 300768 4208
rect 299624 4168 300768 4196
rect 299624 4156 299630 4168
rect 300762 4156 300768 4168
rect 300820 4156 300826 4208
rect 316126 4156 316132 4208
rect 316184 4196 316190 4208
rect 317322 4196 317328 4208
rect 316184 4168 317328 4196
rect 316184 4156 316190 4168
rect 317322 4156 317328 4168
rect 317380 4156 317386 4208
rect 2866 4088 2872 4140
rect 2924 4128 2930 4140
rect 7558 4128 7564 4140
rect 2924 4100 7564 4128
rect 2924 4088 2930 4100
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 67266 4088 67272 4140
rect 67324 4128 67330 4140
rect 106918 4128 106924 4140
rect 67324 4100 106924 4128
rect 67324 4088 67330 4100
rect 106918 4088 106924 4100
rect 106976 4088 106982 4140
rect 141234 4088 141240 4140
rect 141292 4128 141298 4140
rect 142798 4128 142804 4140
rect 141292 4100 142804 4128
rect 141292 4088 141298 4100
rect 142798 4088 142804 4100
rect 142856 4088 142862 4140
rect 177666 4088 177672 4140
rect 177724 4128 177730 4140
rect 450906 4128 450912 4140
rect 177724 4100 450912 4128
rect 177724 4088 177730 4100
rect 450906 4088 450912 4100
rect 450964 4088 450970 4140
rect 566458 4088 566464 4140
rect 566516 4128 566522 4140
rect 568022 4128 568028 4140
rect 566516 4100 568028 4128
rect 566516 4088 566522 4100
rect 568022 4088 568028 4100
rect 568080 4088 568086 4140
rect 576118 4088 576124 4140
rect 576176 4128 576182 4140
rect 577406 4128 577412 4140
rect 576176 4100 577412 4128
rect 576176 4088 576182 4100
rect 577406 4088 577412 4100
rect 577464 4088 577470 4140
rect 39574 4020 39580 4072
rect 39632 4060 39638 4072
rect 82078 4060 82084 4072
rect 39632 4032 82084 4060
rect 39632 4020 39638 4032
rect 82078 4020 82084 4032
rect 82136 4020 82142 4072
rect 176562 4020 176568 4072
rect 176620 4060 176626 4072
rect 454494 4060 454500 4072
rect 176620 4032 454500 4060
rect 176620 4020 176626 4032
rect 454494 4020 454500 4032
rect 454552 4020 454558 4072
rect 66162 3952 66168 4004
rect 66220 3992 66226 4004
rect 110506 3992 110512 4004
rect 66220 3964 110512 3992
rect 66220 3952 66226 3964
rect 110506 3952 110512 3964
rect 110564 3952 110570 4004
rect 174906 3952 174912 4004
rect 174964 3992 174970 4004
rect 458082 3992 458088 4004
rect 174964 3964 458088 3992
rect 174964 3952 174970 3964
rect 458082 3952 458088 3964
rect 458140 3952 458146 4004
rect 35986 3884 35992 3936
rect 36044 3924 36050 3936
rect 83458 3924 83464 3936
rect 36044 3896 83464 3924
rect 36044 3884 36050 3896
rect 83458 3884 83464 3896
rect 83516 3884 83522 3936
rect 175090 3884 175096 3936
rect 175148 3924 175154 3936
rect 461578 3924 461584 3936
rect 175148 3896 461584 3924
rect 175148 3884 175154 3896
rect 461578 3884 461584 3896
rect 461636 3884 461642 3936
rect 64690 3816 64696 3868
rect 64748 3856 64754 3868
rect 114002 3856 114008 3868
rect 64748 3828 114008 3856
rect 64748 3816 64754 3828
rect 114002 3816 114008 3828
rect 114060 3816 114066 3868
rect 173710 3816 173716 3868
rect 173768 3856 173774 3868
rect 465166 3856 465172 3868
rect 173768 3828 465172 3856
rect 173768 3816 173774 3828
rect 465166 3816 465172 3828
rect 465224 3816 465230 3868
rect 32398 3748 32404 3800
rect 32456 3788 32462 3800
rect 83642 3788 83648 3800
rect 32456 3760 83648 3788
rect 32456 3748 32462 3760
rect 83642 3748 83648 3760
rect 83700 3748 83706 3800
rect 173526 3748 173532 3800
rect 173584 3788 173590 3800
rect 468662 3788 468668 3800
rect 173584 3760 468668 3788
rect 173584 3748 173590 3760
rect 468662 3748 468668 3760
rect 468720 3748 468726 3800
rect 64506 3680 64512 3732
rect 64564 3720 64570 3732
rect 117590 3720 117596 3732
rect 64564 3692 117596 3720
rect 64564 3680 64570 3692
rect 117590 3680 117596 3692
rect 117648 3680 117654 3732
rect 172422 3680 172428 3732
rect 172480 3720 172486 3732
rect 472250 3720 472256 3732
rect 172480 3692 472256 3720
rect 172480 3680 172486 3692
rect 472250 3680 472256 3692
rect 472308 3680 472314 3732
rect 63402 3612 63408 3664
rect 63460 3652 63466 3664
rect 121086 3652 121092 3664
rect 63460 3624 121092 3652
rect 63460 3612 63466 3624
rect 121086 3612 121092 3624
rect 121144 3612 121150 3664
rect 142430 3612 142436 3664
rect 142488 3652 142494 3664
rect 146938 3652 146944 3664
rect 142488 3624 146944 3652
rect 142488 3612 142494 3624
rect 146938 3612 146944 3624
rect 146996 3612 147002 3664
rect 170950 3612 170956 3664
rect 171008 3652 171014 3664
rect 475746 3652 475752 3664
rect 171008 3624 475752 3652
rect 171008 3612 171014 3624
rect 475746 3612 475752 3624
rect 475804 3612 475810 3664
rect 28902 3544 28908 3596
rect 28960 3584 28966 3596
rect 84838 3584 84844 3596
rect 28960 3556 84844 3584
rect 28960 3544 28966 3556
rect 84838 3544 84844 3556
rect 84896 3544 84902 3596
rect 115198 3544 115204 3596
rect 115256 3584 115262 3596
rect 117958 3584 117964 3596
rect 115256 3556 117964 3584
rect 115256 3544 115262 3556
rect 117958 3544 117964 3556
rect 118016 3544 118022 3596
rect 144546 3544 144552 3596
rect 144604 3584 144610 3596
rect 144604 3556 144684 3584
rect 144604 3544 144610 3556
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 3418 3516 3424 3528
rect 624 3488 3424 3516
rect 624 3476 630 3488
rect 3418 3476 3424 3488
rect 3476 3476 3482 3528
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 10318 3516 10324 3528
rect 7708 3488 10324 3516
rect 7708 3476 7714 3488
rect 10318 3476 10324 3488
rect 10376 3476 10382 3528
rect 11146 3476 11152 3528
rect 11204 3516 11210 3528
rect 61378 3516 61384 3528
rect 11204 3488 61384 3516
rect 11204 3476 11210 3488
rect 61378 3476 61384 3488
rect 61436 3476 61442 3528
rect 63310 3476 63316 3528
rect 63368 3516 63374 3528
rect 124674 3516 124680 3528
rect 63368 3488 124680 3516
rect 63368 3476 63374 3488
rect 124674 3476 124680 3488
rect 124732 3476 124738 3528
rect 4062 3408 4068 3460
rect 4120 3448 4126 3460
rect 11698 3448 11704 3460
rect 4120 3420 11704 3448
rect 4120 3408 4126 3420
rect 11698 3408 11704 3420
rect 11756 3408 11762 3460
rect 24210 3408 24216 3460
rect 24268 3448 24274 3460
rect 85022 3448 85028 3460
rect 24268 3420 85028 3448
rect 24268 3408 24274 3420
rect 85022 3408 85028 3420
rect 85080 3408 85086 3460
rect 89622 3408 89628 3460
rect 89680 3448 89686 3460
rect 123478 3448 123484 3460
rect 89680 3420 123484 3448
rect 89680 3408 89686 3420
rect 123478 3408 123484 3420
rect 123536 3408 123542 3460
rect 144656 3448 144684 3556
rect 146202 3544 146208 3596
rect 146260 3584 146266 3596
rect 580994 3584 581000 3596
rect 146260 3556 581000 3584
rect 146260 3544 146266 3556
rect 580994 3544 581000 3556
rect 581052 3544 581058 3596
rect 145926 3476 145932 3528
rect 145984 3516 145990 3528
rect 148318 3516 148324 3528
rect 145984 3488 148324 3516
rect 145984 3476 145990 3488
rect 148318 3476 148324 3488
rect 148376 3476 148382 3528
rect 149514 3476 149520 3528
rect 149572 3516 149578 3528
rect 151078 3516 151084 3528
rect 149572 3488 151084 3516
rect 149572 3476 149578 3488
rect 151078 3476 151084 3488
rect 151136 3476 151142 3528
rect 160094 3476 160100 3528
rect 160152 3516 160158 3528
rect 161290 3516 161296 3528
rect 160152 3488 161296 3516
rect 160152 3476 160158 3488
rect 161290 3476 161296 3488
rect 161348 3476 161354 3528
rect 170858 3476 170864 3528
rect 170916 3516 170922 3528
rect 479334 3516 479340 3528
rect 170916 3488 479340 3516
rect 170916 3476 170922 3488
rect 479334 3476 479340 3488
rect 479392 3476 479398 3528
rect 489914 3476 489920 3528
rect 489972 3516 489978 3528
rect 490742 3516 490748 3528
rect 489972 3488 490748 3516
rect 489972 3476 489978 3488
rect 490742 3476 490748 3488
rect 490800 3476 490806 3528
rect 498194 3476 498200 3528
rect 498252 3516 498258 3528
rect 499022 3516 499028 3528
rect 498252 3488 499028 3516
rect 498252 3476 498258 3488
rect 499022 3476 499028 3488
rect 499080 3476 499086 3528
rect 539594 3476 539600 3528
rect 539652 3516 539658 3528
rect 540422 3516 540428 3528
rect 539652 3488 540428 3516
rect 539652 3476 539658 3488
rect 540422 3476 540428 3488
rect 540480 3476 540486 3528
rect 548518 3476 548524 3528
rect 548576 3516 548582 3528
rect 550266 3516 550272 3528
rect 548576 3488 550272 3516
rect 548576 3476 548582 3488
rect 550266 3476 550272 3488
rect 550324 3476 550330 3528
rect 556154 3476 556160 3528
rect 556212 3516 556218 3528
rect 556982 3516 556988 3528
rect 556212 3488 556988 3516
rect 556212 3476 556218 3488
rect 556982 3476 556988 3488
rect 557040 3476 557046 3528
rect 564434 3476 564440 3528
rect 564492 3516 564498 3528
rect 565262 3516 565268 3528
rect 564492 3488 565268 3516
rect 564492 3476 564498 3488
rect 565262 3476 565268 3488
rect 565320 3476 565326 3528
rect 582190 3448 582196 3460
rect 144656 3420 582196 3448
rect 582190 3408 582196 3420
rect 582248 3408 582254 3460
rect 41874 3340 41880 3392
rect 41932 3380 41938 3392
rect 43438 3380 43444 3392
rect 41932 3352 43444 3380
rect 41932 3340 41938 3352
rect 43438 3340 43444 3352
rect 43496 3340 43502 3392
rect 80974 3380 80980 3392
rect 45526 3352 80980 3380
rect 13538 3272 13544 3324
rect 13596 3312 13602 3324
rect 18598 3312 18604 3324
rect 13596 3284 18604 3312
rect 13596 3272 13602 3284
rect 18598 3272 18604 3284
rect 18656 3272 18662 3324
rect 43070 3272 43076 3324
rect 43128 3312 43134 3324
rect 45526 3312 45554 3352
rect 80974 3340 80980 3352
rect 81032 3340 81038 3392
rect 117222 3340 117228 3392
rect 117280 3380 117286 3392
rect 118786 3380 118792 3392
rect 117280 3352 118792 3380
rect 117280 3340 117286 3352
rect 118786 3340 118792 3352
rect 118844 3340 118850 3392
rect 177942 3340 177948 3392
rect 178000 3380 178006 3392
rect 447410 3380 447416 3392
rect 178000 3352 447416 3380
rect 178000 3340 178006 3352
rect 447410 3340 447416 3352
rect 447468 3340 447474 3392
rect 448606 3340 448612 3392
rect 448664 3380 448670 3392
rect 449802 3380 449808 3392
rect 448664 3352 449808 3380
rect 448664 3340 448670 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 43128 3284 45554 3312
rect 43128 3272 43134 3284
rect 46658 3272 46664 3324
rect 46716 3312 46722 3324
rect 80698 3312 80704 3324
rect 46716 3284 80704 3312
rect 46716 3272 46722 3284
rect 80698 3272 80704 3284
rect 80756 3272 80762 3324
rect 115842 3272 115848 3324
rect 115900 3312 115906 3324
rect 122282 3312 122288 3324
rect 115900 3284 122288 3312
rect 115900 3272 115906 3284
rect 122282 3272 122288 3284
rect 122340 3272 122346 3324
rect 156598 3272 156604 3324
rect 156656 3312 156662 3324
rect 244918 3312 244924 3324
rect 156656 3284 244924 3312
rect 156656 3272 156662 3284
rect 244918 3272 244924 3284
rect 244976 3272 244982 3324
rect 307754 3272 307760 3324
rect 307812 3312 307818 3324
rect 309042 3312 309048 3324
rect 307812 3284 309048 3312
rect 307812 3272 307818 3284
rect 309042 3272 309048 3284
rect 309100 3272 309106 3324
rect 324406 3272 324412 3324
rect 324464 3312 324470 3324
rect 325602 3312 325608 3324
rect 324464 3284 325608 3312
rect 324464 3272 324470 3284
rect 325602 3272 325608 3284
rect 325660 3272 325666 3324
rect 332594 3272 332600 3324
rect 332652 3312 332658 3324
rect 333882 3312 333888 3324
rect 332652 3284 333888 3312
rect 332652 3272 332658 3284
rect 333882 3272 333888 3284
rect 333940 3272 333946 3324
rect 340966 3272 340972 3324
rect 341024 3312 341030 3324
rect 342162 3312 342168 3324
rect 341024 3284 342168 3312
rect 341024 3272 341030 3284
rect 342162 3272 342168 3284
rect 342220 3272 342226 3324
rect 349246 3272 349252 3324
rect 349304 3312 349310 3324
rect 350442 3312 350448 3324
rect 349304 3284 350448 3312
rect 349304 3272 349310 3284
rect 350442 3272 350448 3284
rect 350500 3272 350506 3324
rect 357526 3272 357532 3324
rect 357584 3312 357590 3324
rect 358722 3312 358728 3324
rect 357584 3284 358728 3312
rect 357584 3272 357590 3284
rect 358722 3272 358728 3284
rect 358780 3272 358786 3324
rect 365806 3272 365812 3324
rect 365864 3312 365870 3324
rect 367002 3312 367008 3324
rect 365864 3284 367008 3312
rect 365864 3272 365870 3284
rect 367002 3272 367008 3284
rect 367060 3272 367066 3324
rect 374086 3272 374092 3324
rect 374144 3312 374150 3324
rect 375282 3312 375288 3324
rect 374144 3284 375288 3312
rect 374144 3272 374150 3284
rect 375282 3272 375288 3284
rect 375340 3272 375346 3324
rect 382366 3272 382372 3324
rect 382424 3312 382430 3324
rect 383562 3312 383568 3324
rect 382424 3284 383568 3312
rect 382424 3272 382430 3284
rect 383562 3272 383568 3284
rect 383620 3272 383626 3324
rect 390646 3272 390652 3324
rect 390704 3312 390710 3324
rect 391842 3312 391848 3324
rect 390704 3284 391848 3312
rect 390704 3272 390710 3284
rect 391842 3272 391848 3284
rect 391900 3272 391906 3324
rect 398834 3272 398840 3324
rect 398892 3312 398898 3324
rect 400122 3312 400128 3324
rect 398892 3284 400128 3312
rect 398892 3272 398898 3284
rect 400122 3272 400128 3284
rect 400180 3272 400186 3324
rect 407206 3272 407212 3324
rect 407264 3312 407270 3324
rect 408402 3312 408408 3324
rect 407264 3284 408408 3312
rect 407264 3272 407270 3284
rect 408402 3272 408408 3284
rect 408460 3272 408466 3324
rect 415486 3272 415492 3324
rect 415544 3312 415550 3324
rect 416682 3312 416688 3324
rect 415544 3284 416688 3312
rect 415544 3272 415550 3284
rect 416682 3272 416688 3284
rect 416740 3272 416746 3324
rect 423766 3272 423772 3324
rect 423824 3312 423830 3324
rect 424962 3312 424968 3324
rect 423824 3284 424968 3312
rect 423824 3272 423830 3284
rect 424962 3272 424968 3284
rect 425020 3272 425026 3324
rect 431954 3272 431960 3324
rect 432012 3312 432018 3324
rect 433242 3312 433248 3324
rect 432012 3284 433248 3312
rect 432012 3272 432018 3284
rect 433242 3272 433248 3284
rect 433300 3272 433306 3324
rect 440234 3272 440240 3324
rect 440292 3312 440298 3324
rect 441522 3312 441528 3324
rect 440292 3284 441528 3312
rect 440292 3272 440298 3284
rect 441522 3272 441528 3284
rect 441580 3272 441586 3324
rect 67450 3204 67456 3256
rect 67508 3244 67514 3256
rect 103330 3244 103336 3256
rect 67508 3216 103336 3244
rect 67508 3204 67514 3216
rect 103330 3204 103336 3216
rect 103388 3204 103394 3256
rect 160094 3204 160100 3256
rect 160152 3244 160158 3256
rect 243538 3244 243544 3256
rect 160152 3216 243544 3244
rect 160152 3204 160158 3216
rect 243538 3204 243544 3216
rect 243596 3204 243602 3256
rect 136450 3136 136456 3188
rect 136508 3176 136514 3188
rect 137278 3176 137284 3188
rect 136508 3148 137284 3176
rect 136508 3136 136514 3148
rect 137278 3136 137284 3148
rect 137336 3136 137342 3188
rect 138842 3136 138848 3188
rect 138900 3176 138906 3188
rect 141418 3176 141424 3188
rect 138900 3148 141424 3176
rect 138900 3136 138906 3148
rect 141418 3136 141424 3148
rect 141476 3136 141482 3188
rect 8754 3000 8760 3052
rect 8812 3040 8818 3052
rect 14458 3040 14464 3052
rect 8812 3012 14464 3040
rect 8812 3000 8818 3012
rect 14458 3000 14464 3012
rect 14516 3000 14522 3052
<< via1 >>
rect 1400 444388 1452 444440
rect 57612 444388 57664 444440
rect 63316 59712 63368 59764
rect 64328 59712 64380 59764
rect 72792 59712 72844 59764
rect 75092 59712 75144 59764
rect 78588 59712 78640 59764
rect 79968 59712 80020 59764
rect 92388 59712 92440 59764
rect 93860 59712 93912 59764
rect 98644 59712 98696 59764
rect 101404 59712 101456 59764
rect 102784 59712 102836 59764
rect 105636 59780 105688 59832
rect 110328 59780 110380 59832
rect 111340 59780 111392 59832
rect 229468 59780 229520 59832
rect 230664 59780 230716 59832
rect 105544 59712 105596 59764
rect 108028 59712 108080 59764
rect 111064 59712 111116 59764
rect 113732 59712 113784 59764
rect 114008 59712 114060 59764
rect 116216 59712 116268 59764
rect 119528 59712 119580 59764
rect 122012 59712 122064 59764
rect 124864 59712 124916 59764
rect 126428 59712 126480 59764
rect 127624 59712 127676 59764
rect 130200 59712 130252 59764
rect 140688 59712 140740 59764
rect 141700 59712 141752 59764
rect 150072 59712 150124 59764
rect 151912 59712 151964 59764
rect 157156 59712 157208 59764
rect 158168 59712 158220 59764
rect 172428 59712 172480 59764
rect 173348 59712 173400 59764
rect 182088 59712 182140 59764
rect 183744 59712 183796 59764
rect 192852 59712 192904 59764
rect 194416 59712 194468 59764
rect 199844 59712 199896 59764
rect 200212 59712 200264 59764
rect 201316 59712 201368 59764
rect 202788 59712 202840 59764
rect 208216 59712 208268 59764
rect 209412 59712 209464 59764
rect 213552 59712 213604 59764
rect 215852 59712 215904 59764
rect 232504 59712 232556 59764
rect 234804 59712 234856 59764
rect 238024 59712 238076 59764
rect 240508 59780 240560 59832
rect 296996 59780 297048 59832
rect 298928 59780 298980 59832
rect 380072 59780 380124 59832
rect 382924 59780 382976 59832
rect 239404 59712 239456 59764
rect 242164 59712 242216 59764
rect 244188 59712 244240 59764
rect 245476 59712 245528 59764
rect 249064 59712 249116 59764
rect 251272 59712 251324 59764
rect 267464 59712 267516 59764
rect 269948 59712 270000 59764
rect 270684 59712 270736 59764
rect 271880 59712 271932 59764
rect 277216 59712 277268 59764
rect 277860 59712 277912 59764
rect 283012 59712 283064 59764
rect 284300 59712 284352 59764
rect 287888 59712 287940 59764
rect 290648 59712 290700 59764
rect 293684 59712 293736 59764
rect 295984 59712 296036 59764
rect 296536 59712 296588 59764
rect 298744 59712 298796 59764
rect 301964 59712 302016 59764
rect 304264 59712 304316 59764
rect 314292 59712 314344 59764
rect 316684 59712 316736 59764
rect 320824 59712 320876 59764
rect 323124 59712 323176 59764
rect 324964 59712 325016 59764
rect 327356 59712 327408 59764
rect 334900 59712 334952 59764
rect 336924 59712 336976 59764
rect 339040 59712 339092 59764
rect 341156 59712 341208 59764
rect 341524 59712 341576 59764
rect 342536 59712 342588 59764
rect 343088 59712 343140 59764
rect 345112 59712 345164 59764
rect 359556 59712 359608 59764
rect 361764 59712 361816 59764
rect 363696 59712 363748 59764
rect 366364 59712 366416 59764
rect 367008 59712 367060 59764
rect 369124 59712 369176 59764
rect 369400 59712 369452 59764
rect 24860 59644 24912 59696
rect 61016 59644 61068 59696
rect 95884 59644 95936 59696
rect 97356 59644 97408 59696
rect 236644 59644 236696 59696
rect 238852 59644 238904 59696
rect 269856 59644 269908 59696
rect 272524 59644 272576 59696
rect 286324 59644 286376 59696
rect 288440 59644 288492 59696
rect 300308 59644 300360 59696
rect 302884 59644 302936 59696
rect 312544 59644 312596 59696
rect 313924 59644 313976 59696
rect 365168 59644 365220 59696
rect 366548 59644 366600 59696
rect 371056 59712 371108 59764
rect 372620 59712 372672 59764
rect 376024 59712 376076 59764
rect 378968 59712 379020 59764
rect 379428 59712 379480 59764
rect 380164 59712 380216 59764
rect 380992 59712 381044 59764
rect 382280 59712 382332 59764
rect 387524 59712 387576 59764
rect 389824 59712 389876 59764
rect 391664 59712 391716 59764
rect 393964 59712 394016 59764
rect 397460 59712 397512 59764
rect 399484 59712 399536 59764
rect 402336 59712 402388 59764
rect 404452 59712 404504 59764
rect 406476 59712 406528 59764
rect 408500 59712 408552 59764
rect 410616 59712 410668 59764
rect 412824 59712 412876 59764
rect 425520 59712 425572 59764
rect 426532 59712 426584 59764
rect 427084 59712 427136 59764
rect 429568 59712 429620 59764
rect 431224 59712 431276 59764
rect 433616 59712 433668 59764
rect 436928 59712 436980 59764
rect 439228 59712 439280 59764
rect 441896 59712 441948 59764
rect 443184 59712 443236 59764
rect 446864 59712 446916 59764
rect 448796 59712 448848 59764
rect 457536 59712 457588 59764
rect 459928 59712 459980 59764
rect 464160 59712 464212 59764
rect 465356 59712 465408 59764
rect 371332 59644 371384 59696
rect 390008 59644 390060 59696
rect 392584 59644 392636 59696
rect 19340 59576 19392 59628
rect 60464 59576 60516 59628
rect 67456 59576 67508 59628
rect 69296 59576 69348 59628
rect 75368 59576 75420 59628
rect 77484 59576 77536 59628
rect 87604 59576 87656 59628
rect 89076 59576 89128 59628
rect 118148 59576 118200 59628
rect 120356 59576 120408 59628
rect 130568 59576 130620 59628
rect 131948 59576 132000 59628
rect 140044 59576 140096 59628
rect 141700 59576 141752 59628
rect 150256 59576 150308 59628
rect 151636 59576 151688 59628
rect 165436 59576 165488 59628
rect 166448 59576 166500 59628
rect 174912 59576 174964 59628
rect 177120 59576 177172 59628
rect 217692 59576 217744 59628
rect 219164 59576 219216 59628
rect 227628 59576 227680 59628
rect 229008 59576 229060 59628
rect 246488 59576 246540 59628
rect 248880 59576 248932 59628
rect 256332 59576 256384 59628
rect 257804 59576 257856 59628
rect 259092 59576 259144 59628
rect 261116 59576 261168 59628
rect 280344 59576 280396 59628
rect 282184 59576 282236 59628
rect 306012 59576 306064 59628
rect 307208 59576 307260 59628
rect 310152 59576 310204 59628
rect 312728 59576 312780 59628
rect 376024 59576 376076 59628
rect 377404 59576 377456 59628
rect 393320 59576 393372 59628
rect 395344 59576 395396 59628
rect 413100 59576 413152 59628
rect 414112 59576 414164 59628
rect 416412 59576 416464 59628
rect 418252 59576 418304 59628
rect 449256 59576 449308 59628
rect 449900 59576 449952 59628
rect 453396 59576 453448 59628
rect 455696 59576 455748 59628
rect 15200 59508 15252 59560
rect 59360 59508 59412 59560
rect 247868 59508 247920 59560
rect 250536 59508 250588 59560
rect 5540 59440 5592 59492
rect 57612 59440 57664 59492
rect 85028 59440 85080 59492
rect 87420 59440 87472 59492
rect 89536 59440 89588 59492
rect 91560 59440 91612 59492
rect 166632 59440 166684 59492
rect 168932 59440 168984 59492
rect 169392 59440 169444 59492
rect 171416 59440 171468 59492
rect 179328 59440 179380 59492
rect 180432 59440 180484 59492
rect 188896 59440 188948 59492
rect 190276 59440 190328 59492
rect 4160 59372 4212 59424
rect 57980 59372 58032 59424
rect 138112 59372 138164 59424
rect 139308 59372 139360 59424
rect 188712 59372 188764 59424
rect 190552 59440 190604 59492
rect 205272 59440 205324 59492
rect 207572 59440 207624 59492
rect 246304 59440 246356 59492
rect 247960 59440 248012 59492
rect 272248 59440 272300 59492
rect 273260 59440 273312 59492
rect 273904 59440 273956 59492
rect 276664 59440 276716 59492
rect 308496 59440 308548 59492
rect 311164 59440 311216 59492
rect 329104 59440 329156 59492
rect 331312 59440 331364 59492
rect 344744 59440 344796 59492
rect 346492 59440 346544 59492
rect 351368 59440 351420 59492
rect 353576 59440 353628 59492
rect 372712 59440 372764 59492
rect 374000 59440 374052 59492
rect 398104 59440 398156 59492
rect 401048 59440 401100 59492
rect 408132 59440 408184 59492
rect 409880 59440 409932 59492
rect 428740 59440 428792 59492
rect 430672 59440 430724 59492
rect 432052 59440 432104 59492
rect 433432 59440 433484 59492
rect 455052 59440 455104 59492
rect 456984 59440 457036 59492
rect 459192 59440 459244 59492
rect 461216 59440 461268 59492
rect 306840 59304 306892 59356
rect 308404 59304 308456 59356
rect 310520 59304 310572 59356
rect 316960 59304 317012 59356
rect 325792 59304 325844 59356
rect 327172 59304 327224 59356
rect 384120 59304 384172 59356
rect 385684 59304 385736 59356
rect 123484 59236 123536 59288
rect 126152 59236 126204 59288
rect 82084 58964 82136 59016
rect 84200 58964 84252 59016
rect 401600 58964 401652 59016
rect 405740 58964 405792 59016
rect 147588 58896 147640 58948
rect 148692 58896 148744 58948
rect 251180 58896 251232 58948
rect 330300 58896 330352 58948
rect 383660 58896 383712 58948
rect 483020 58896 483072 58948
rect 320180 58828 320232 58880
rect 419540 58828 419592 58880
rect 162860 58760 162912 58812
rect 244188 58760 244240 58812
rect 271880 58760 271932 58812
rect 513380 58760 513432 58812
rect 56600 58692 56652 58744
rect 78588 58692 78640 58744
rect 193220 58692 193272 58744
rect 449716 58692 449768 58744
rect 7564 58624 7616 58676
rect 142068 58624 142120 58676
rect 157248 58624 157300 58676
rect 546500 58624 546552 58676
rect 80888 58488 80940 58540
rect 83280 58488 83332 58540
rect 291752 58488 291804 58540
rect 293224 58488 293276 58540
rect 293408 58488 293460 58540
rect 294788 58488 294840 58540
rect 148692 58352 148744 58404
rect 149980 58352 150032 58404
rect 314660 57536 314712 57588
rect 328460 57536 328512 57588
rect 331220 57536 331272 57588
rect 416872 57536 416924 57588
rect 233240 57468 233292 57520
rect 335360 57468 335412 57520
rect 382280 57468 382332 57520
rect 489920 57468 489972 57520
rect 190368 57400 190420 57452
rect 393320 57400 393372 57452
rect 273260 57332 273312 57384
rect 506480 57332 506532 57384
rect 34520 57264 34572 57316
rect 110328 57264 110380 57316
rect 195980 57264 196032 57316
rect 451280 57264 451332 57316
rect 51080 57196 51132 57248
rect 131120 57196 131172 57248
rect 164056 57196 164108 57248
rect 517520 57196 517572 57248
rect 349160 56176 349212 56228
rect 412916 56176 412968 56228
rect 172520 56108 172572 56160
rect 348424 56108 348476 56160
rect 380808 56108 380860 56160
rect 500960 56108 501012 56160
rect 194416 56040 194468 56092
rect 386420 56040 386472 56092
rect 274640 55972 274692 56024
rect 502340 55972 502392 56024
rect 209780 55904 209832 55956
rect 447140 55904 447192 55956
rect 53840 55836 53892 55888
rect 132040 55836 132092 55888
rect 162768 55836 162820 55888
rect 524420 55836 524472 55888
rect 205456 54748 205508 54800
rect 329840 54748 329892 54800
rect 376760 54748 376812 54800
rect 408684 54748 408736 54800
rect 284300 54680 284352 54732
rect 459560 54680 459612 54732
rect 226156 54612 226208 54664
rect 241520 54612 241572 54664
rect 252560 54612 252612 54664
rect 437480 54612 437532 54664
rect 110512 54544 110564 54596
rect 118148 54544 118200 54596
rect 126980 54544 127032 54596
rect 361580 54544 361632 54596
rect 374000 54544 374052 54596
rect 525800 54544 525852 54596
rect 33140 54476 33192 54528
rect 136088 54476 136140 54528
rect 180800 54476 180852 54528
rect 239588 54476 239640 54528
rect 253848 54476 253900 54528
rect 572720 54476 572772 54528
rect 308588 53388 308640 53440
rect 360200 53388 360252 53440
rect 225972 53320 226024 53372
rect 237380 53320 237432 53372
rect 258080 53320 258132 53372
rect 331496 53320 331548 53372
rect 205640 53252 205692 53304
rect 234068 53252 234120 53304
rect 288440 53252 288492 53304
rect 445760 53252 445812 53304
rect 197084 53184 197136 53236
rect 365720 53184 365772 53236
rect 372620 53184 372672 53236
rect 532700 53184 532752 53236
rect 222016 53116 222068 53168
rect 255320 53116 255372 53168
rect 259460 53116 259512 53168
rect 436192 53116 436244 53168
rect 57980 53048 58032 53100
rect 130568 53048 130620 53100
rect 146300 53048 146352 53100
rect 462320 53048 462372 53100
rect 298928 52028 298980 52080
rect 398840 52028 398892 52080
rect 236000 51960 236052 52012
rect 336924 51960 336976 52012
rect 371332 51960 371384 52012
rect 539600 51960 539652 52012
rect 263600 51892 263652 51944
rect 434720 51892 434772 51944
rect 183376 51824 183428 51876
rect 422300 51824 422352 51876
rect 143540 51756 143592 51808
rect 463792 51756 463844 51808
rect 16580 51688 16632 51740
rect 140688 51688 140740 51740
rect 158628 51688 158680 51740
rect 528560 51688 528612 51740
rect 203984 50600 204036 50652
rect 332600 50600 332652 50652
rect 380900 50600 380952 50652
rect 408500 50600 408552 50652
rect 286508 50532 286560 50584
rect 457076 50532 457128 50584
rect 204260 50464 204312 50516
rect 343640 50464 343692 50516
rect 370688 50464 370740 50516
rect 543740 50464 543792 50516
rect 20720 50396 20772 50448
rect 138848 50396 138900 50448
rect 146944 50396 146996 50448
rect 247868 50396 247920 50448
rect 278136 50396 278188 50448
rect 488540 50396 488592 50448
rect 137284 50328 137336 50380
rect 465080 50328 465132 50380
rect 208216 49308 208268 49360
rect 316040 49308 316092 49360
rect 394700 49308 394752 49360
rect 404360 49308 404412 49360
rect 290648 49240 290700 49292
rect 438860 49240 438912 49292
rect 256700 49172 256752 49224
rect 436376 49172 436428 49224
rect 136640 49104 136692 49156
rect 358912 49104 358964 49156
rect 369124 49104 369176 49156
rect 550640 49104 550692 49156
rect 186136 49036 186188 49088
rect 411260 49036 411312 49088
rect 29000 48968 29052 49020
rect 137376 48968 137428 49020
rect 150440 48968 150492 49020
rect 461032 48968 461084 49020
rect 204168 47880 204220 47932
rect 336740 47880 336792 47932
rect 168380 47812 168432 47864
rect 351920 47812 351972 47864
rect 398288 47812 398340 47864
rect 423680 47812 423732 47864
rect 242900 47744 242952 47796
rect 440240 47744 440292 47796
rect 154580 47676 154632 47728
rect 354864 47676 354916 47728
rect 367928 47676 367980 47728
rect 554780 47676 554832 47728
rect 279424 47608 279476 47660
rect 484400 47608 484452 47660
rect 26240 47540 26292 47592
rect 138664 47540 138716 47592
rect 185952 47540 186004 47592
rect 415400 47540 415452 47592
rect 308404 46520 308456 46572
rect 357440 46520 357492 46572
rect 276020 46452 276072 46504
rect 327172 46452 327224 46504
rect 387248 46452 387300 46504
rect 473360 46452 473412 46504
rect 296996 46384 297048 46436
rect 407120 46384 407172 46436
rect 161480 46316 161532 46368
rect 353392 46316 353444 46368
rect 366548 46316 366600 46368
rect 561680 46316 561732 46368
rect 224960 46248 225012 46300
rect 444472 46248 444524 46300
rect 35900 46180 35952 46232
rect 135904 46180 135956 46232
rect 154304 46180 154356 46232
rect 548524 46180 548576 46232
rect 271880 45160 271932 45212
rect 328644 45160 328696 45212
rect 307208 45092 307260 45144
rect 364340 45092 364392 45144
rect 217876 45024 217928 45076
rect 273260 45024 273312 45076
rect 290464 45024 290516 45076
rect 434720 45024 434772 45076
rect 197268 44956 197320 45008
rect 361580 44956 361632 45008
rect 388628 44956 388680 45008
rect 465264 44956 465316 45008
rect 165620 44888 165672 44940
rect 353576 44888 353628 44940
rect 366364 44888 366416 44940
rect 564440 44888 564492 44940
rect 40040 44820 40092 44872
rect 134708 44820 134760 44872
rect 220820 44820 220872 44872
rect 444380 44820 444432 44872
rect 201316 43732 201368 43784
rect 343640 43732 343692 43784
rect 270500 43664 270552 43716
rect 433432 43664 433484 43716
rect 158720 43596 158772 43648
rect 354956 43596 355008 43648
rect 390008 43596 390060 43648
rect 458180 43596 458232 43648
rect 181996 43528 182048 43580
rect 431960 43528 432012 43580
rect 175280 43460 175332 43512
rect 455512 43460 455564 43512
rect 11704 43392 11756 43444
rect 115204 43392 115256 43444
rect 255136 43392 255188 43444
rect 569960 43392 570012 43444
rect 209596 42372 209648 42424
rect 307760 42372 307812 42424
rect 299480 42304 299532 42356
rect 426532 42304 426584 42356
rect 195796 42236 195848 42288
rect 372620 42236 372672 42288
rect 142804 42168 142856 42220
rect 358820 42168 358872 42220
rect 392768 42168 392820 42220
rect 448520 42168 448572 42220
rect 272524 42100 272576 42152
rect 516140 42100 516192 42152
rect 3424 42032 3476 42084
rect 142896 42032 142948 42084
rect 182180 42032 182232 42084
rect 454040 42032 454092 42084
rect 253940 41012 253992 41064
rect 332692 41012 332744 41064
rect 303068 40944 303120 40996
rect 382280 40944 382332 40996
rect 193036 40876 193088 40928
rect 379520 40876 379572 40928
rect 387064 40876 387116 40928
rect 476120 40876 476172 40928
rect 282368 40808 282420 40860
rect 470600 40808 470652 40860
rect 178040 40740 178092 40792
rect 455696 40740 455748 40792
rect 14464 40672 14516 40724
rect 114008 40672 114060 40724
rect 139400 40672 139452 40724
rect 463976 40672 464028 40724
rect 278780 39652 278832 39704
rect 327356 39652 327408 39704
rect 216496 39584 216548 39636
rect 284300 39584 284352 39636
rect 313280 39584 313332 39636
rect 423772 39584 423824 39636
rect 195612 39516 195664 39568
rect 368480 39516 368532 39568
rect 395344 39516 395396 39568
rect 437480 39516 437532 39568
rect 212540 39448 212592 39500
rect 232688 39448 232740 39500
rect 283564 39448 283616 39500
rect 466460 39448 466512 39500
rect 221832 39380 221884 39432
rect 259552 39380 259604 39432
rect 276848 39380 276900 39432
rect 495440 39380 495492 39432
rect 18604 39312 18656 39364
rect 113824 39312 113876 39364
rect 171140 39312 171192 39364
rect 456984 39312 457036 39364
rect 282920 38224 282972 38276
rect 325700 38224 325752 38276
rect 302240 38156 302292 38208
rect 426440 38156 426492 38208
rect 199844 38088 199896 38140
rect 350632 38088 350684 38140
rect 394148 38088 394200 38140
rect 440240 38088 440292 38140
rect 276664 38020 276716 38072
rect 498200 38020 498252 38072
rect 168472 37952 168524 38004
rect 456800 37952 456852 38004
rect 27620 37884 27672 37936
rect 111248 37884 111300 37936
rect 162676 37884 162728 37936
rect 510620 37884 510672 37936
rect 296168 36864 296220 36916
rect 410064 36864 410116 36916
rect 206928 36796 206980 36848
rect 322940 36796 322992 36848
rect 176660 36728 176712 36780
rect 350540 36728 350592 36780
rect 367744 36728 367796 36780
rect 557540 36728 557592 36780
rect 141424 36660 141476 36712
rect 249064 36660 249116 36712
rect 280988 36660 281040 36712
rect 481640 36660 481692 36712
rect 187516 36592 187568 36644
rect 404360 36592 404412 36644
rect 10324 36524 10376 36576
rect 141516 36524 141568 36576
rect 218060 36524 218112 36576
rect 445852 36524 445904 36576
rect 205272 35436 205324 35488
rect 325700 35436 325752 35488
rect 391204 35436 391256 35488
rect 455420 35436 455472 35488
rect 277400 35368 277452 35420
rect 432052 35368 432104 35420
rect 164240 35300 164292 35352
rect 458272 35300 458324 35352
rect 254952 35232 255004 35284
rect 565820 35232 565872 35284
rect 43444 35164 43496 35216
rect 107108 35164 107160 35216
rect 162492 35164 162544 35216
rect 514760 35164 514812 35216
rect 315304 34076 315356 34128
rect 332692 34076 332744 34128
rect 298744 34008 298796 34060
rect 402980 34008 403032 34060
rect 267740 33940 267792 33992
rect 328828 33940 328880 33992
rect 370504 33940 370556 33992
rect 547880 33940 547932 33992
rect 213920 33872 213972 33924
rect 447416 33872 447468 33924
rect 157340 33804 157392 33856
rect 459744 33804 459796 33856
rect 49700 33736 49752 33788
rect 79508 33736 79560 33788
rect 150256 33736 150308 33788
rect 564532 33736 564584 33788
rect 300308 32716 300360 32768
rect 396080 32716 396132 32768
rect 260840 32648 260892 32700
rect 331312 32648 331364 32700
rect 374644 32648 374696 32700
rect 529940 32648 529992 32700
rect 207020 32580 207072 32632
rect 448796 32580 448848 32632
rect 179144 32512 179196 32564
rect 440332 32512 440384 32564
rect 153200 32444 153252 32496
rect 461216 32444 461268 32496
rect 157156 32376 157208 32428
rect 539692 32376 539744 32428
rect 202788 31288 202840 31340
rect 340880 31288 340932 31340
rect 374000 31288 374052 31340
rect 409880 31288 409932 31340
rect 286324 31220 286376 31272
rect 452660 31220 452712 31272
rect 179420 31152 179472 31204
rect 349252 31152 349304 31204
rect 376208 31152 376260 31204
rect 523040 31152 523092 31204
rect 219348 31084 219400 31136
rect 269120 31084 269172 31136
rect 278044 31084 278096 31136
rect 491300 31084 491352 31136
rect 202880 31016 202932 31068
rect 448612 31016 448664 31068
rect 396908 29996 396960 30048
rect 433340 29996 433392 30048
rect 208032 29928 208084 29980
rect 318800 29928 318852 29980
rect 274640 29860 274692 29912
rect 433616 29860 433668 29912
rect 198740 29792 198792 29844
rect 235448 29792 235500 29844
rect 284944 29792 284996 29844
rect 463700 29792 463752 29844
rect 184848 29724 184900 29776
rect 418344 29724 418396 29776
rect 220636 29656 220688 29708
rect 262220 29656 262272 29708
rect 269948 29656 270000 29708
rect 527180 29656 527232 29708
rect 160100 29588 160152 29640
rect 459928 29588 459980 29640
rect 333980 28500 334032 28552
rect 418160 28500 418212 28552
rect 129740 28432 129792 28484
rect 361764 28432 361816 28484
rect 380164 28432 380216 28484
rect 505100 28432 505152 28484
rect 273904 28364 273956 28416
rect 509240 28364 509292 28416
rect 200120 28296 200172 28348
rect 449900 28296 449952 28348
rect 68836 28228 68888 28280
rect 99380 28228 99432 28280
rect 150072 28228 150124 28280
rect 566464 28228 566516 28280
rect 327080 27208 327132 27260
rect 421104 27208 421156 27260
rect 215300 27140 215352 27192
rect 340972 27140 341024 27192
rect 381544 27140 381596 27192
rect 498292 27140 498344 27192
rect 188896 27072 188948 27124
rect 400220 27072 400272 27124
rect 268568 27004 268620 27056
rect 531320 27004 531372 27056
rect 128360 26936 128412 26988
rect 466552 26936 466604 26988
rect 17960 26868 18012 26920
rect 112444 26868 112496 26920
rect 147588 26868 147640 26920
rect 578240 26868 578292 26920
rect 316868 25984 316920 26036
rect 321560 25984 321612 26036
rect 242992 25848 243044 25900
rect 335360 25848 335412 25900
rect 324320 25780 324372 25832
rect 420920 25780 420972 25832
rect 198648 25712 198700 25764
rect 357532 25712 357584 25764
rect 382924 25712 382976 25764
rect 494060 25712 494112 25764
rect 271144 25644 271196 25696
rect 520280 25644 520332 25696
rect 189080 25576 189132 25628
rect 452936 25576 452988 25628
rect 90916 25508 90968 25560
rect 111800 25508 111852 25560
rect 158352 25508 158404 25560
rect 531412 25508 531464 25560
rect 264980 24420 265032 24472
rect 329932 24420 329984 24472
rect 384304 24420 384356 24472
rect 487160 24420 487212 24472
rect 316132 24352 316184 24404
rect 422392 24352 422444 24404
rect 187332 24284 187384 24336
rect 407212 24284 407264 24336
rect 148324 24216 148376 24268
rect 247684 24216 247736 24268
rect 269764 24216 269816 24268
rect 523132 24216 523184 24268
rect 184940 24148 184992 24200
rect 452752 24148 452804 24200
rect 70308 24080 70360 24132
rect 92480 24080 92532 24132
rect 93676 24080 93728 24132
rect 104900 24080 104952 24132
rect 161204 24080 161256 24132
rect 521660 24080 521712 24132
rect 402244 23060 402296 23112
rect 408500 23060 408552 23112
rect 200028 22992 200080 23044
rect 354680 22992 354732 23044
rect 389824 22992 389876 23044
rect 462320 22992 462372 23044
rect 267832 22924 267884 22976
rect 434904 22924 434956 22976
rect 252468 22856 252520 22908
rect 576124 22856 576176 22908
rect 125600 22788 125652 22840
rect 467840 22788 467892 22840
rect 71596 22720 71648 22772
rect 85580 22720 85632 22772
rect 156972 22720 157024 22772
rect 535460 22720 535512 22772
rect 95148 22516 95200 22568
rect 98000 22516 98052 22568
rect 316684 22108 316736 22160
rect 324412 22108 324464 22160
rect 299572 21700 299624 21752
rect 321652 21700 321704 21752
rect 287704 21632 287756 21684
rect 448612 21632 448664 21684
rect 188712 21564 188764 21616
rect 397460 21564 397512 21616
rect 182088 21496 182140 21548
rect 429200 21496 429252 21548
rect 86960 21428 87012 21480
rect 97448 21428 97500 21480
rect 180708 21428 180760 21480
rect 436100 21428 436152 21480
rect 9680 21360 9732 21412
rect 87788 21360 87840 21412
rect 179328 21360 179380 21412
rect 443000 21360 443052 21412
rect 398932 20612 398984 20664
rect 404452 20612 404504 20664
rect 296720 20272 296772 20324
rect 323124 20272 323176 20324
rect 340972 20272 341024 20324
rect 416780 20272 416832 20324
rect 201132 20204 201184 20256
rect 347780 20204 347832 20256
rect 194508 20136 194560 20188
rect 375380 20136 375432 20188
rect 388444 20136 388496 20188
rect 469220 20136 469272 20188
rect 192852 20068 192904 20120
rect 382372 20068 382424 20120
rect 385684 20068 385736 20120
rect 480260 20068 480312 20120
rect 282184 20000 282236 20052
rect 473452 20000 473504 20052
rect 44180 19932 44232 19984
rect 134524 19932 134576 19984
rect 191748 19932 191800 19984
rect 390560 19932 390612 19984
rect 398104 19932 398156 19984
rect 426440 19932 426492 19984
rect 155868 18912 155920 18964
rect 542360 18912 542412 18964
rect 153016 18844 153068 18896
rect 553400 18844 553452 18896
rect 152832 18776 152884 18828
rect 556160 18776 556212 18828
rect 151728 18708 151780 18760
rect 560300 18708 560352 18760
rect 148876 18640 148928 18692
rect 571340 18640 571392 18692
rect 60740 18572 60792 18624
rect 76748 18572 76800 18624
rect 80060 18572 80112 18624
rect 98828 18572 98880 18624
rect 103520 18572 103572 18624
rect 119528 18572 119580 18624
rect 148692 18572 148744 18624
rect 574100 18572 574152 18624
rect 280804 17756 280856 17808
rect 477500 17756 477552 17808
rect 169392 17688 169444 17740
rect 481732 17688 481784 17740
rect 169576 17620 169628 17672
rect 485780 17620 485832 17672
rect 168288 17552 168340 17604
rect 490012 17552 490064 17604
rect 166632 17484 166684 17536
rect 492680 17484 492732 17536
rect 166816 17416 166868 17468
rect 496820 17416 496872 17468
rect 165252 17348 165304 17400
rect 499580 17348 499632 17400
rect 100760 17280 100812 17332
rect 120724 17280 120776 17332
rect 165436 17280 165488 17332
rect 503720 17280 503772 17332
rect 66260 17212 66312 17264
rect 101588 17212 101640 17264
rect 164148 17212 164200 17264
rect 506572 17212 506624 17264
rect 295984 16260 296036 16312
rect 414296 16260 414348 16312
rect 294788 16192 294840 16244
rect 417424 16192 417476 16244
rect 294604 16124 294656 16176
rect 420920 16124 420972 16176
rect 220452 16056 220504 16108
rect 266544 16056 266596 16108
rect 293224 16056 293276 16108
rect 423772 16056 423824 16108
rect 188528 15988 188580 16040
rect 238208 15988 238260 16040
rect 292028 15988 292080 16040
rect 428464 15988 428516 16040
rect 73344 15920 73396 15972
rect 100024 15920 100076 15972
rect 177580 15920 177632 15972
rect 239404 15920 239456 15972
rect 291844 15920 291896 15972
rect 432052 15920 432104 15972
rect 93952 15852 94004 15904
rect 122288 15852 122340 15904
rect 135260 15852 135312 15904
rect 250628 15852 250680 15904
rect 289084 15852 289136 15904
rect 442632 15852 442684 15904
rect 268384 14968 268436 15020
rect 534448 14968 534500 15020
rect 267004 14900 267056 14952
rect 538220 14900 538272 14952
rect 265624 14832 265676 14884
rect 541992 14832 542044 14884
rect 260748 14764 260800 14816
rect 545488 14764 545540 14816
rect 259092 14696 259144 14748
rect 548432 14696 548484 14748
rect 259276 14628 259328 14680
rect 552664 14628 552716 14680
rect 185032 14560 185084 14612
rect 238024 14560 238076 14612
rect 257988 14560 258040 14612
rect 556252 14560 556304 14612
rect 53288 14492 53340 14544
rect 79324 14492 79376 14544
rect 151084 14492 151136 14544
rect 246488 14492 246540 14544
rect 256516 14492 256568 14544
rect 559288 14492 559340 14544
rect 79232 14424 79284 14476
rect 126428 14424 126480 14476
rect 127532 14424 127584 14476
rect 251824 14424 251876 14476
rect 256332 14424 256384 14476
rect 563060 14424 563112 14476
rect 307024 13608 307076 13660
rect 367744 13608 367796 13660
rect 305644 13540 305696 13592
rect 371240 13540 371292 13592
rect 304448 13472 304500 13524
rect 374092 13472 374144 13524
rect 304264 13404 304316 13456
rect 378416 13404 378468 13456
rect 401048 13404 401100 13456
rect 415492 13404 415544 13456
rect 302884 13336 302936 13388
rect 385960 13336 386012 13388
rect 387800 13336 387852 13388
rect 405924 13336 405976 13388
rect 301504 13268 301556 13320
rect 389456 13268 389508 13320
rect 390652 13268 390704 13320
rect 406108 13268 406160 13320
rect 64328 13200 64380 13252
rect 76564 13200 76616 13252
rect 216864 13200 216916 13252
rect 231124 13200 231176 13252
rect 300124 13200 300176 13252
rect 392492 13200 392544 13252
rect 399484 13200 399536 13252
rect 420184 13200 420236 13252
rect 68652 13132 68704 13184
rect 95792 13132 95844 13184
rect 151820 13132 151872 13184
rect 356060 13132 356112 13184
rect 384304 13132 384356 13184
rect 407304 13132 407356 13184
rect 75920 13064 75972 13116
rect 126244 13064 126296 13116
rect 147864 13064 147916 13116
rect 357808 13064 357860 13116
rect 393964 13064 394016 13116
rect 445024 13064 445076 13116
rect 312544 12180 312596 12232
rect 339500 12180 339552 12232
rect 312728 12112 312780 12164
rect 342260 12112 342312 12164
rect 311348 12044 311400 12096
rect 346952 12044 347004 12096
rect 400864 12044 400916 12096
rect 412640 12044 412692 12096
rect 211068 11976 211120 12028
rect 305552 11976 305604 12028
rect 311164 11976 311216 12028
rect 349252 11976 349304 12028
rect 396724 11976 396776 12028
rect 430856 11976 430908 12028
rect 153016 11908 153068 11960
rect 246304 11908 246356 11960
rect 309784 11908 309836 11960
rect 353576 11908 353628 11960
rect 365812 11908 365864 11960
rect 411352 11908 411404 11960
rect 209412 11840 209464 11892
rect 312176 11840 312228 11892
rect 313924 11840 313976 11892
rect 335452 11840 335504 11892
rect 338672 11840 338724 11892
rect 418252 11840 418304 11892
rect 144460 11772 144512 11824
rect 357624 11772 357676 11824
rect 392584 11772 392636 11824
rect 451648 11772 451700 11824
rect 65064 11704 65116 11756
rect 129004 11704 129056 11756
rect 168380 11704 168432 11756
rect 169576 11704 169628 11756
rect 184940 11704 184992 11756
rect 186136 11704 186188 11756
rect 183192 11636 183244 11688
rect 425704 11704 425756 11756
rect 259460 11636 259512 11688
rect 260656 11636 260708 11688
rect 91560 11024 91612 11076
rect 95884 11024 95936 11076
rect 217692 10684 217744 10736
rect 276664 10684 276716 10736
rect 216312 10616 216364 10668
rect 280712 10616 280764 10668
rect 286600 10616 286652 10668
rect 324780 10616 324832 10668
rect 370136 10616 370188 10668
rect 409972 10616 410024 10668
rect 215208 10548 215260 10600
rect 287336 10548 287388 10600
rect 289820 10548 289872 10600
rect 324596 10548 324648 10600
rect 363512 10548 363564 10600
rect 412916 10548 412968 10600
rect 213552 10480 213604 10532
rect 291384 10480 291436 10532
rect 293224 10480 293276 10532
rect 323308 10480 323360 10532
rect 359464 10480 359516 10532
rect 412732 10480 412784 10532
rect 213736 10412 213788 10464
rect 294880 10412 294932 10464
rect 314660 10412 314712 10464
rect 318892 10412 318944 10464
rect 356336 10412 356388 10464
rect 414020 10412 414072 10464
rect 72976 10344 73028 10396
rect 81624 10344 81676 10396
rect 84200 10344 84252 10396
rect 97264 10344 97316 10396
rect 212172 10344 212224 10396
rect 298100 10344 298152 10396
rect 307944 10344 307996 10396
rect 320548 10344 320600 10396
rect 352840 10344 352892 10396
rect 414112 10344 414164 10396
rect 47400 10276 47452 10328
rect 133144 10276 133196 10328
rect 212356 10276 212408 10328
rect 301504 10276 301556 10328
rect 303896 10276 303948 10328
rect 320364 10276 320416 10328
rect 345020 10276 345072 10328
rect 416964 10276 417016 10328
rect 310244 9324 310296 9376
rect 425152 9324 425204 9376
rect 306748 9256 306800 9308
rect 425336 9256 425388 9308
rect 227628 9188 227680 9240
rect 234620 9188 234672 9240
rect 296076 9188 296128 9240
rect 427912 9188 427964 9240
rect 224776 9120 224828 9172
rect 245200 9120 245252 9172
rect 292580 9120 292632 9172
rect 429568 9120 429620 9172
rect 77392 9052 77444 9104
rect 72792 8984 72844 9036
rect 78588 8984 78640 9036
rect 93768 9052 93820 9104
rect 102232 9052 102284 9104
rect 224868 9052 224920 9104
rect 248788 9052 248840 9104
rect 288992 9052 289044 9104
rect 429384 9052 429436 9104
rect 98644 8984 98696 9036
rect 223488 8984 223540 9036
rect 252376 8984 252428 9036
rect 285404 8984 285456 9036
rect 430672 8984 430724 9036
rect 62028 8916 62080 8968
rect 130384 8916 130436 8968
rect 131764 8916 131816 8968
rect 250444 8916 250496 8968
rect 281908 8916 281960 8968
rect 430580 8916 430632 8968
rect 223948 8372 224000 8424
rect 229928 8372 229980 8424
rect 229008 8304 229060 8356
rect 231032 8304 231084 8356
rect 227536 8168 227588 8220
rect 228364 8168 228416 8220
rect 92388 7964 92440 8016
rect 109316 7964 109368 8016
rect 249984 7964 250036 8016
rect 439228 7964 439280 8016
rect 90732 7896 90784 7948
rect 116400 7896 116452 7948
rect 170772 7896 170824 7948
rect 242348 7896 242400 7948
rect 246396 7896 246448 7948
rect 439044 7896 439096 7948
rect 89536 7828 89588 7880
rect 119896 7828 119948 7880
rect 195612 7828 195664 7880
rect 235264 7828 235316 7880
rect 239312 7828 239364 7880
rect 440424 7828 440476 7880
rect 45468 7760 45520 7812
rect 106924 7760 106976 7812
rect 209872 7760 209924 7812
rect 232504 7760 232556 7812
rect 235816 7760 235868 7812
rect 441712 7760 441764 7812
rect 38384 7692 38436 7744
rect 108304 7692 108356 7744
rect 232228 7692 232280 7744
rect 443184 7692 443236 7744
rect 31300 7624 31352 7676
rect 109684 7624 109736 7676
rect 228732 7624 228784 7676
rect 443368 7624 443420 7676
rect 23020 7556 23072 7608
rect 111064 7556 111116 7608
rect 132960 7556 133012 7608
rect 465356 7556 465408 7608
rect 93860 7488 93912 7540
rect 94780 7488 94832 7540
rect 220452 6740 220504 6792
rect 229744 6740 229796 6792
rect 202696 6672 202748 6724
rect 233884 6672 233936 6724
rect 174268 6604 174320 6656
rect 240784 6604 240836 6656
rect 167184 6536 167236 6588
rect 242164 6536 242216 6588
rect 247592 6536 247644 6588
rect 334072 6536 334124 6588
rect 70308 6468 70360 6520
rect 101404 6468 101456 6520
rect 192024 6468 192076 6520
rect 236644 6468 236696 6520
rect 240508 6468 240560 6520
rect 335544 6468 335596 6520
rect 63224 6400 63276 6452
rect 102968 6400 103020 6452
rect 229836 6400 229888 6452
rect 338212 6400 338264 6452
rect 59636 6332 59688 6384
rect 102784 6332 102836 6384
rect 226340 6332 226392 6384
rect 338120 6332 338172 6384
rect 56048 6264 56100 6316
rect 104164 6264 104216 6316
rect 222752 6264 222804 6316
rect 339592 6264 339644 6316
rect 364984 6264 365036 6316
rect 569132 6264 569184 6316
rect 52552 6196 52604 6248
rect 105820 6196 105872 6248
rect 219256 6196 219308 6248
rect 341156 6196 341208 6248
rect 363788 6196 363840 6248
rect 572720 6196 572772 6248
rect 48964 6128 49016 6180
rect 105544 6128 105596 6180
rect 108120 6128 108172 6180
rect 119344 6128 119396 6180
rect 134156 6128 134208 6180
rect 360292 6128 360344 6180
rect 363604 6128 363656 6180
rect 576308 6128 576360 6180
rect 403072 5856 403124 5908
rect 402980 5652 403032 5704
rect 340144 5312 340196 5364
rect 346400 5312 346452 5364
rect 212172 5244 212224 5296
rect 342352 5244 342404 5296
rect 71412 5176 71464 5228
rect 89168 5176 89220 5228
rect 97448 5176 97500 5228
rect 122104 5176 122156 5228
rect 208584 5176 208636 5228
rect 342536 5176 342588 5228
rect 72608 5108 72660 5160
rect 69112 5040 69164 5092
rect 71504 4904 71556 4956
rect 75184 4904 75236 4956
rect 86868 5108 86920 5160
rect 123484 5108 123536 5160
rect 201500 5108 201552 5160
rect 345112 5108 345164 5160
rect 83280 5040 83332 5092
rect 124864 5040 124916 5092
rect 197912 5040 197964 5092
rect 345388 5040 345440 5092
rect 378784 5040 378836 5092
rect 508872 5040 508924 5092
rect 127808 4972 127860 5024
rect 194416 4972 194468 5024
rect 346492 4972 346544 5024
rect 378968 4972 379020 5024
rect 512460 4972 512512 5024
rect 127624 4904 127676 4956
rect 190828 4904 190880 4956
rect 340144 4904 340196 4956
rect 377404 4904 377456 4956
rect 515956 4904 516008 4956
rect 14740 4836 14792 4888
rect 87604 4836 87656 4888
rect 90364 4836 90416 4888
rect 123668 4836 123720 4888
rect 187332 4836 187384 4888
rect 347872 4836 347924 4888
rect 376116 4836 376168 4888
rect 519544 4836 519596 4888
rect 12348 4768 12400 4820
rect 140044 4768 140096 4820
rect 183744 4768 183796 4820
rect 349436 4768 349488 4820
rect 371884 4768 371936 4820
rect 537208 4768 537260 4820
rect 74448 4632 74500 4684
rect 75000 4632 75052 4684
rect 67916 4428 67968 4480
rect 75368 4428 75420 4480
rect 209780 4156 209832 4208
rect 210976 4156 211028 4208
rect 267740 4156 267792 4208
rect 268476 4156 268528 4208
rect 299572 4156 299624 4208
rect 300768 4156 300820 4208
rect 316132 4156 316184 4208
rect 317328 4156 317380 4208
rect 2872 4088 2924 4140
rect 7564 4088 7616 4140
rect 67272 4088 67324 4140
rect 106924 4088 106976 4140
rect 141240 4088 141292 4140
rect 142804 4088 142856 4140
rect 177672 4088 177724 4140
rect 450912 4088 450964 4140
rect 566464 4088 566516 4140
rect 568028 4088 568080 4140
rect 576124 4088 576176 4140
rect 577412 4088 577464 4140
rect 39580 4020 39632 4072
rect 82084 4020 82136 4072
rect 176568 4020 176620 4072
rect 454500 4020 454552 4072
rect 66168 3952 66220 4004
rect 110512 3952 110564 4004
rect 174912 3952 174964 4004
rect 458088 3952 458140 4004
rect 35992 3884 36044 3936
rect 83464 3884 83516 3936
rect 175096 3884 175148 3936
rect 461584 3884 461636 3936
rect 64696 3816 64748 3868
rect 114008 3816 114060 3868
rect 173716 3816 173768 3868
rect 465172 3816 465224 3868
rect 32404 3748 32456 3800
rect 83648 3748 83700 3800
rect 173532 3748 173584 3800
rect 468668 3748 468720 3800
rect 64512 3680 64564 3732
rect 117596 3680 117648 3732
rect 172428 3680 172480 3732
rect 472256 3680 472308 3732
rect 63408 3612 63460 3664
rect 121092 3612 121144 3664
rect 142436 3612 142488 3664
rect 146944 3612 146996 3664
rect 170956 3612 171008 3664
rect 475752 3612 475804 3664
rect 28908 3544 28960 3596
rect 84844 3544 84896 3596
rect 115204 3544 115256 3596
rect 117964 3544 118016 3596
rect 144552 3544 144604 3596
rect 572 3476 624 3528
rect 3424 3476 3476 3528
rect 7656 3476 7708 3528
rect 10324 3476 10376 3528
rect 11152 3476 11204 3528
rect 61384 3476 61436 3528
rect 63316 3476 63368 3528
rect 124680 3476 124732 3528
rect 4068 3408 4120 3460
rect 11704 3408 11756 3460
rect 24216 3408 24268 3460
rect 85028 3408 85080 3460
rect 89628 3408 89680 3460
rect 123484 3408 123536 3460
rect 146208 3544 146260 3596
rect 581000 3544 581052 3596
rect 145932 3476 145984 3528
rect 148324 3476 148376 3528
rect 149520 3476 149572 3528
rect 151084 3476 151136 3528
rect 160100 3476 160152 3528
rect 161296 3476 161348 3528
rect 170864 3476 170916 3528
rect 479340 3476 479392 3528
rect 489920 3476 489972 3528
rect 490748 3476 490800 3528
rect 498200 3476 498252 3528
rect 499028 3476 499080 3528
rect 539600 3476 539652 3528
rect 540428 3476 540480 3528
rect 548524 3476 548576 3528
rect 550272 3476 550324 3528
rect 556160 3476 556212 3528
rect 556988 3476 557040 3528
rect 564440 3476 564492 3528
rect 565268 3476 565320 3528
rect 582196 3408 582248 3460
rect 41880 3340 41932 3392
rect 43444 3340 43496 3392
rect 13544 3272 13596 3324
rect 18604 3272 18656 3324
rect 43076 3272 43128 3324
rect 80980 3340 81032 3392
rect 117228 3340 117280 3392
rect 118792 3340 118844 3392
rect 177948 3340 178000 3392
rect 447416 3340 447468 3392
rect 448612 3340 448664 3392
rect 449808 3340 449860 3392
rect 46664 3272 46716 3324
rect 80704 3272 80756 3324
rect 115848 3272 115900 3324
rect 122288 3272 122340 3324
rect 156604 3272 156656 3324
rect 244924 3272 244976 3324
rect 307760 3272 307812 3324
rect 309048 3272 309100 3324
rect 324412 3272 324464 3324
rect 325608 3272 325660 3324
rect 332600 3272 332652 3324
rect 333888 3272 333940 3324
rect 340972 3272 341024 3324
rect 342168 3272 342220 3324
rect 349252 3272 349304 3324
rect 350448 3272 350500 3324
rect 357532 3272 357584 3324
rect 358728 3272 358780 3324
rect 365812 3272 365864 3324
rect 367008 3272 367060 3324
rect 374092 3272 374144 3324
rect 375288 3272 375340 3324
rect 382372 3272 382424 3324
rect 383568 3272 383620 3324
rect 390652 3272 390704 3324
rect 391848 3272 391900 3324
rect 398840 3272 398892 3324
rect 400128 3272 400180 3324
rect 407212 3272 407264 3324
rect 408408 3272 408460 3324
rect 415492 3272 415544 3324
rect 416688 3272 416740 3324
rect 423772 3272 423824 3324
rect 424968 3272 425020 3324
rect 431960 3272 432012 3324
rect 433248 3272 433300 3324
rect 440240 3272 440292 3324
rect 441528 3272 441580 3324
rect 67456 3204 67508 3256
rect 103336 3204 103388 3256
rect 160100 3204 160152 3256
rect 243544 3204 243596 3256
rect 136456 3136 136508 3188
rect 137284 3136 137336 3188
rect 138848 3136 138900 3188
rect 141424 3136 141476 3188
rect 8760 3000 8812 3052
rect 14464 3000 14516 3052
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 57610 445496 57666 445505
rect 57610 445431 57666 445440
rect 57624 444446 57652 445431
rect 1400 444440 1452 444446
rect 1400 444382 1452 444388
rect 57612 444440 57664 444446
rect 57612 444382 57664 444388
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 584 480 612 3470
rect 542 -960 654 480
rect 1412 354 1440 444382
rect 57610 59936 57666 59945
rect 57610 59871 57666 59880
rect 24860 59696 24912 59702
rect 24860 59638 24912 59644
rect 19340 59628 19392 59634
rect 19340 59570 19392 59576
rect 15200 59560 15252 59566
rect 15200 59502 15252 59508
rect 5540 59492 5592 59498
rect 5540 59434 5592 59440
rect 4160 59424 4212 59430
rect 4160 59366 4212 59372
rect 3424 42084 3476 42090
rect 3424 42026 3476 42032
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 2884 480 2912 4082
rect 3436 3534 3464 42026
rect 4172 16574 4200 59366
rect 5552 16574 5580 59434
rect 7564 58676 7616 58682
rect 7564 58618 7616 58624
rect 4172 16546 5304 16574
rect 5552 16546 6040 16574
rect 3424 3528 3476 3534
rect 3424 3470 3476 3476
rect 4068 3460 4120 3466
rect 4068 3402 4120 3408
rect 4080 480 4108 3402
rect 5276 480 5304 16546
rect 1646 354 1758 480
rect 1412 326 1758 354
rect 1646 -960 1758 326
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6012 354 6040 16546
rect 7576 4146 7604 58618
rect 11704 43444 11756 43450
rect 11704 43386 11756 43392
rect 10324 36576 10376 36582
rect 10324 36518 10376 36524
rect 9680 21412 9732 21418
rect 9680 21354 9732 21360
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7668 480 7696 3470
rect 8760 3052 8812 3058
rect 8760 2994 8812 3000
rect 8772 480 8800 2994
rect 6430 354 6542 480
rect 6012 326 6542 354
rect 6430 -960 6542 326
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 21354
rect 10336 3534 10364 36518
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 11164 480 11192 3470
rect 11716 3466 11744 43386
rect 14464 40724 14516 40730
rect 14464 40666 14516 40672
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 11704 3460 11756 3466
rect 11704 3402 11756 3408
rect 12360 480 12388 4762
rect 13544 3324 13596 3330
rect 13544 3266 13596 3272
rect 13556 480 13584 3266
rect 14476 3058 14504 40666
rect 15212 16574 15240 59502
rect 16580 51740 16632 51746
rect 16580 51682 16632 51688
rect 16592 16574 16620 51682
rect 18604 39364 18656 39370
rect 18604 39306 18656 39312
rect 17960 26920 18012 26926
rect 17960 26862 18012 26868
rect 15212 16546 15976 16574
rect 16592 16546 17080 16574
rect 14740 4888 14792 4894
rect 14740 4830 14792 4836
rect 14464 3052 14516 3058
rect 14464 2994 14516 3000
rect 14752 480 14780 4830
rect 15948 480 15976 16546
rect 17052 480 17080 16546
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 26862
rect 18616 3330 18644 39306
rect 19352 16574 19380 59570
rect 20720 50448 20772 50454
rect 20720 50390 20772 50396
rect 20732 16574 20760 50390
rect 24872 16574 24900 59638
rect 57624 59498 57652 59871
rect 105636 59832 105688 59838
rect 57978 59800 58034 59809
rect 57978 59735 58034 59744
rect 61014 59800 61070 59809
rect 64326 59800 64382 59809
rect 61014 59735 61070 59744
rect 63316 59764 63368 59770
rect 57612 59492 57664 59498
rect 57612 59434 57664 59440
rect 57992 59430 58020 59735
rect 61028 59702 61056 59735
rect 64326 59735 64328 59744
rect 63316 59706 63368 59712
rect 64380 59735 64382 59744
rect 70214 59800 70270 59809
rect 75090 59800 75146 59809
rect 70214 59735 70270 59744
rect 72792 59764 72844 59770
rect 64328 59706 64380 59712
rect 61016 59696 61068 59702
rect 60462 59664 60518 59673
rect 61016 59638 61068 59644
rect 62670 59664 62726 59673
rect 60462 59599 60464 59608
rect 60516 59599 60518 59608
rect 62670 59599 62726 59608
rect 60464 59570 60516 59576
rect 59360 59560 59412 59566
rect 59360 59502 59412 59508
rect 61382 59528 61438 59537
rect 57980 59424 58032 59430
rect 59372 59401 59400 59502
rect 61382 59463 61438 59472
rect 57980 59366 58032 59372
rect 59358 59392 59414 59401
rect 59358 59327 59414 59336
rect 56600 58744 56652 58750
rect 56600 58686 56652 58692
rect 34520 57316 34572 57322
rect 34520 57258 34572 57264
rect 33140 54528 33192 54534
rect 33140 54470 33192 54476
rect 29000 49020 29052 49026
rect 29000 48962 29052 48968
rect 26240 47592 26292 47598
rect 26240 47534 26292 47540
rect 19352 16546 20208 16574
rect 20732 16546 21864 16574
rect 24872 16546 25360 16574
rect 19430 3360 19486 3369
rect 18604 3324 18656 3330
rect 19430 3295 19486 3304
rect 18604 3266 18656 3272
rect 19444 480 19472 3295
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20180 354 20208 16546
rect 21836 480 21864 16546
rect 23020 7608 23072 7614
rect 23020 7550 23072 7556
rect 23032 480 23060 7550
rect 24216 3460 24268 3466
rect 24216 3402 24268 3408
rect 24228 480 24256 3402
rect 25332 480 25360 16546
rect 20598 354 20710 480
rect 20180 326 20710 354
rect 20598 -960 20710 326
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 47534
rect 27620 37936 27672 37942
rect 27620 37878 27672 37884
rect 27632 16574 27660 37878
rect 29012 16574 29040 48962
rect 33152 16574 33180 54470
rect 27632 16546 27752 16574
rect 29012 16546 30144 16574
rect 33152 16546 33640 16574
rect 27724 480 27752 16546
rect 28908 3596 28960 3602
rect 28908 3538 28960 3544
rect 28920 480 28948 3538
rect 30116 480 30144 16546
rect 31300 7676 31352 7682
rect 31300 7618 31352 7624
rect 31312 480 31340 7618
rect 32404 3800 32456 3806
rect 32404 3742 32456 3748
rect 32416 480 32444 3742
rect 33612 480 33640 16546
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34532 354 34560 57258
rect 51080 57248 51132 57254
rect 51080 57190 51132 57196
rect 35900 46232 35952 46238
rect 35900 46174 35952 46180
rect 35912 16574 35940 46174
rect 40040 44872 40092 44878
rect 40040 44814 40092 44820
rect 40052 16574 40080 44814
rect 43444 35216 43496 35222
rect 43444 35158 43496 35164
rect 35912 16546 36768 16574
rect 40052 16546 40264 16574
rect 35992 3936 36044 3942
rect 35992 3878 36044 3884
rect 36004 480 36032 3878
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 38384 7744 38436 7750
rect 38384 7686 38436 7692
rect 38396 480 38424 7686
rect 39580 4072 39632 4078
rect 39580 4014 39632 4020
rect 39592 480 39620 4014
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40236 354 40264 16546
rect 43456 3398 43484 35158
rect 49700 33788 49752 33794
rect 49700 33730 49752 33736
rect 44180 19984 44232 19990
rect 44180 19926 44232 19932
rect 44192 16574 44220 19926
rect 49712 16574 49740 33730
rect 44192 16546 44312 16574
rect 49712 16546 50200 16574
rect 41880 3392 41932 3398
rect 41880 3334 41932 3340
rect 43444 3392 43496 3398
rect 43444 3334 43496 3340
rect 41892 480 41920 3334
rect 43076 3324 43128 3330
rect 43076 3266 43128 3272
rect 43088 480 43116 3266
rect 44284 480 44312 16546
rect 47400 10328 47452 10334
rect 47400 10270 47452 10276
rect 45468 7812 45520 7818
rect 45468 7754 45520 7760
rect 45480 480 45508 7754
rect 46664 3324 46716 3330
rect 46664 3266 46716 3272
rect 46676 480 46704 3266
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47412 354 47440 10270
rect 48964 6180 49016 6186
rect 48964 6122 49016 6128
rect 48976 480 49004 6122
rect 50172 480 50200 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 47830 -960 47942 326
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51092 354 51120 57190
rect 53840 55888 53892 55894
rect 53840 55830 53892 55836
rect 53852 16574 53880 55830
rect 56612 16574 56640 58686
rect 57980 53100 58032 53106
rect 57980 53042 58032 53048
rect 57992 16574 58020 53042
rect 60740 18624 60792 18630
rect 60740 18566 60792 18572
rect 60752 16574 60780 18566
rect 53852 16546 54984 16574
rect 56612 16546 56824 16574
rect 57992 16546 58480 16574
rect 60752 16546 60872 16574
rect 53288 14544 53340 14550
rect 53288 14486 53340 14492
rect 52552 6248 52604 6254
rect 52552 6190 52604 6196
rect 52564 480 52592 6190
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53300 354 53328 14486
rect 54956 480 54984 16546
rect 56048 6316 56100 6322
rect 56048 6258 56100 6264
rect 56060 480 56088 6258
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58452 480 58480 16546
rect 59636 6384 59688 6390
rect 59636 6326 59688 6332
rect 59648 480 59676 6326
rect 60844 480 60872 16546
rect 61396 3534 61424 59463
rect 62684 59401 62712 59599
rect 62670 59392 62726 59401
rect 62670 59327 62726 59336
rect 62028 8968 62080 8974
rect 62028 8910 62080 8916
rect 61384 3528 61436 3534
rect 61384 3470 61436 3476
rect 62040 480 62068 8910
rect 63224 6452 63276 6458
rect 63224 6394 63276 6400
rect 63236 480 63264 6394
rect 63328 3534 63356 59706
rect 69294 59664 69350 59673
rect 67456 59628 67508 59634
rect 69294 59599 69296 59608
rect 67456 59570 67508 59576
rect 69348 59599 69350 59608
rect 70122 59664 70178 59673
rect 70122 59599 70178 59608
rect 69296 59570 69348 59576
rect 64510 59528 64566 59537
rect 64510 59463 64566 59472
rect 66810 59528 66866 59537
rect 66810 59463 66866 59472
rect 63406 59392 63462 59401
rect 63406 59327 63462 59336
rect 63420 3670 63448 59327
rect 64328 13252 64380 13258
rect 64328 13194 64380 13200
rect 63408 3664 63460 3670
rect 63408 3606 63460 3612
rect 63316 3528 63368 3534
rect 63316 3470 63368 3476
rect 64340 480 64368 13194
rect 64524 3738 64552 59463
rect 64694 59392 64750 59401
rect 64694 59327 64750 59336
rect 66166 59392 66222 59401
rect 66166 59327 66222 59336
rect 64708 3874 64736 59327
rect 65064 11756 65116 11762
rect 65064 11698 65116 11704
rect 64696 3868 64748 3874
rect 64696 3810 64748 3816
rect 64512 3732 64564 3738
rect 64512 3674 64564 3680
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 11698
rect 66180 4010 66208 59327
rect 66824 59265 66852 59463
rect 66810 59256 66866 59265
rect 66810 59191 66866 59200
rect 67270 59256 67326 59265
rect 67270 59191 67326 59200
rect 66260 17264 66312 17270
rect 66260 17206 66312 17212
rect 66272 16574 66300 17206
rect 66272 16546 66760 16574
rect 66168 4004 66220 4010
rect 66168 3946 66220 3952
rect 66732 480 66760 16546
rect 67284 4146 67312 59191
rect 67272 4140 67324 4146
rect 67272 4082 67324 4088
rect 67468 3262 67496 59570
rect 68834 59528 68890 59537
rect 68834 59463 68890 59472
rect 68650 59392 68706 59401
rect 68650 59327 68706 59336
rect 68664 13190 68692 59327
rect 68848 28286 68876 59463
rect 70136 59401 70164 59599
rect 70228 59537 70256 59735
rect 79966 59800 80022 59809
rect 75090 59735 75092 59744
rect 72792 59706 72844 59712
rect 75144 59735 75146 59744
rect 78588 59764 78640 59770
rect 75092 59706 75144 59712
rect 79966 59735 79968 59744
rect 78588 59706 78640 59712
rect 80020 59735 80022 59744
rect 84198 59800 84254 59809
rect 93858 59800 93914 59809
rect 84198 59735 84254 59744
rect 92388 59764 92440 59770
rect 79968 59706 80020 59712
rect 70214 59528 70270 59537
rect 70214 59463 70270 59472
rect 70122 59392 70178 59401
rect 70122 59327 70178 59336
rect 70306 59392 70362 59401
rect 70306 59327 70362 59336
rect 68836 28280 68888 28286
rect 68836 28222 68888 28228
rect 70320 24138 70348 59327
rect 71410 59256 71466 59265
rect 71410 59191 71466 59200
rect 70308 24132 70360 24138
rect 70308 24074 70360 24080
rect 68652 13184 68704 13190
rect 68652 13126 68704 13132
rect 70308 6520 70360 6526
rect 70308 6462 70360 6468
rect 69112 5092 69164 5098
rect 69112 5034 69164 5040
rect 67916 4480 67968 4486
rect 67916 4422 67968 4428
rect 67456 3256 67508 3262
rect 67456 3198 67508 3204
rect 67928 480 67956 4422
rect 69124 480 69152 5034
rect 70320 480 70348 6462
rect 71424 5234 71452 59191
rect 71594 59120 71650 59129
rect 71594 59055 71650 59064
rect 71608 22778 71636 59055
rect 71596 22772 71648 22778
rect 71596 22714 71648 22720
rect 72804 9042 72832 59706
rect 76654 59664 76710 59673
rect 75368 59628 75420 59634
rect 76654 59599 76710 59608
rect 77482 59664 77538 59673
rect 77482 59599 77484 59608
rect 75368 59570 75420 59576
rect 74446 59392 74502 59401
rect 74446 59327 74502 59336
rect 72974 58984 73030 58993
rect 72974 58919 73030 58928
rect 72988 10402 73016 58919
rect 73344 15972 73396 15978
rect 73344 15914 73396 15920
rect 72976 10396 73028 10402
rect 72976 10338 73028 10344
rect 72792 9036 72844 9042
rect 72792 8978 72844 8984
rect 71412 5228 71464 5234
rect 71412 5170 71464 5176
rect 72608 5160 72660 5166
rect 72608 5102 72660 5108
rect 71504 4956 71556 4962
rect 71504 4898 71556 4904
rect 71516 480 71544 4898
rect 72620 480 72648 5102
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 15914
rect 74460 4690 74488 59327
rect 75182 59256 75238 59265
rect 75182 59191 75238 59200
rect 75196 4962 75224 59191
rect 75184 4956 75236 4962
rect 75184 4898 75236 4904
rect 74448 4684 74500 4690
rect 74448 4626 74500 4632
rect 75000 4684 75052 4690
rect 75000 4626 75052 4632
rect 75012 480 75040 4626
rect 75380 4486 75408 59570
rect 76562 59528 76618 59537
rect 76562 59463 76618 59472
rect 76576 13258 76604 59463
rect 76668 59401 76696 59599
rect 77536 59599 77538 59608
rect 77484 59570 77536 59576
rect 76654 59392 76710 59401
rect 76654 59327 76710 59336
rect 76838 59392 76894 59401
rect 76838 59327 76894 59336
rect 76852 45554 76880 59327
rect 78600 58750 78628 59706
rect 79322 59664 79378 59673
rect 79322 59599 79378 59608
rect 81622 59664 81678 59673
rect 81622 59599 81678 59608
rect 83278 59664 83334 59673
rect 84106 59664 84162 59673
rect 83278 59599 83334 59608
rect 83476 59622 84106 59650
rect 78588 58744 78640 58750
rect 78588 58686 78640 58692
rect 76760 45526 76880 45554
rect 76760 18630 76788 45526
rect 76748 18624 76800 18630
rect 76748 18566 76800 18572
rect 79336 14550 79364 59599
rect 80702 59528 80758 59537
rect 80702 59463 80758 59472
rect 79506 59392 79562 59401
rect 79506 59327 79562 59336
rect 79520 33794 79548 59327
rect 79508 33788 79560 33794
rect 79508 33730 79560 33736
rect 80060 18624 80112 18630
rect 80060 18566 80112 18572
rect 80072 16574 80100 18566
rect 80072 16546 80652 16574
rect 79324 14544 79376 14550
rect 79324 14486 79376 14492
rect 79232 14476 79284 14482
rect 79232 14418 79284 14424
rect 76564 13252 76616 13258
rect 76564 13194 76616 13200
rect 75920 13116 75972 13122
rect 75920 13058 75972 13064
rect 75368 4480 75420 4486
rect 75368 4422 75420 4428
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 13058
rect 77392 9104 77444 9110
rect 77392 9046 77444 9052
rect 77404 480 77432 9046
rect 78588 9036 78640 9042
rect 78588 8978 78640 8984
rect 78600 480 78628 8978
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79244 354 79272 14418
rect 80624 1034 80652 16546
rect 80716 3330 80744 59463
rect 81636 59401 81664 59599
rect 81622 59392 81678 59401
rect 81622 59327 81678 59336
rect 82084 59016 82136 59022
rect 82084 58958 82136 58964
rect 80888 58540 80940 58546
rect 80888 58482 80940 58488
rect 80900 16574 80928 58482
rect 80900 16546 81020 16574
rect 80992 3398 81020 16546
rect 81624 10396 81676 10402
rect 81624 10338 81676 10344
rect 80980 3392 81032 3398
rect 80980 3334 81032 3340
rect 80704 3324 80756 3330
rect 80704 3266 80756 3272
rect 80624 1006 80928 1034
rect 80900 480 80928 1006
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 10338
rect 82096 4078 82124 58958
rect 83292 58546 83320 59599
rect 83280 58540 83332 58546
rect 83280 58482 83332 58488
rect 83280 5092 83332 5098
rect 83280 5034 83332 5040
rect 82084 4072 82136 4078
rect 82084 4014 82136 4020
rect 83292 480 83320 5034
rect 83476 3942 83504 59622
rect 84106 59599 84162 59608
rect 83646 59392 83702 59401
rect 83646 59327 83702 59336
rect 83464 3936 83516 3942
rect 83464 3878 83516 3884
rect 83660 3806 83688 59327
rect 84212 59022 84240 59735
rect 93858 59735 93860 59744
rect 92388 59706 92440 59712
rect 93912 59735 93914 59744
rect 97354 59800 97410 59809
rect 101402 59800 101458 59809
rect 97354 59735 97410 59744
rect 98644 59764 98696 59770
rect 93860 59706 93912 59712
rect 85762 59664 85818 59673
rect 89074 59664 89130 59673
rect 85762 59599 85818 59608
rect 87604 59628 87656 59634
rect 84842 59528 84898 59537
rect 84842 59463 84898 59472
rect 85028 59492 85080 59498
rect 84200 59016 84252 59022
rect 84200 58958 84252 58964
rect 84200 10396 84252 10402
rect 84200 10338 84252 10344
rect 83648 3800 83700 3806
rect 83648 3742 83700 3748
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 10338
rect 84856 3602 84884 59463
rect 85028 59434 85080 59440
rect 84844 3596 84896 3602
rect 84844 3538 84896 3544
rect 85040 3466 85068 59434
rect 85776 59401 85804 59599
rect 89074 59599 89076 59608
rect 87604 59570 87656 59576
rect 89128 59599 89130 59608
rect 89902 59664 89958 59673
rect 89902 59599 89958 59608
rect 89076 59570 89128 59576
rect 87418 59528 87474 59537
rect 87418 59463 87420 59472
rect 87472 59463 87474 59472
rect 87420 59434 87472 59440
rect 85762 59392 85818 59401
rect 85762 59327 85818 59336
rect 86222 59392 86278 59401
rect 86222 59327 86278 59336
rect 85580 22772 85632 22778
rect 85580 22714 85632 22720
rect 85592 16574 85620 22714
rect 85592 16546 85712 16574
rect 85028 3460 85080 3466
rect 85028 3402 85080 3408
rect 85684 480 85712 16546
rect 86236 3369 86264 59327
rect 86960 21480 87012 21486
rect 86960 21422 87012 21428
rect 86972 16574 87000 21422
rect 86972 16546 87552 16574
rect 86868 5160 86920 5166
rect 86868 5102 86920 5108
rect 86222 3360 86278 3369
rect 86222 3295 86278 3304
rect 86880 480 86908 5102
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87524 354 87552 16546
rect 87616 4894 87644 59570
rect 89626 59528 89682 59537
rect 89536 59492 89588 59498
rect 89626 59463 89682 59472
rect 89536 59434 89588 59440
rect 87786 59256 87842 59265
rect 87786 59191 87842 59200
rect 87800 21418 87828 59191
rect 87788 21412 87840 21418
rect 87788 21354 87840 21360
rect 89548 7886 89576 59434
rect 89536 7880 89588 7886
rect 89536 7822 89588 7828
rect 89168 5228 89220 5234
rect 89168 5170 89220 5176
rect 87604 4888 87656 4894
rect 87604 4830 87656 4836
rect 89180 480 89208 5170
rect 89640 3466 89668 59463
rect 89916 59401 89944 59599
rect 91558 59528 91614 59537
rect 91558 59463 91560 59472
rect 91612 59463 91614 59472
rect 91560 59434 91612 59440
rect 89902 59392 89958 59401
rect 89902 59327 89958 59336
rect 90730 59392 90786 59401
rect 90730 59327 90786 59336
rect 90744 7954 90772 59327
rect 90914 59256 90970 59265
rect 90914 59191 90970 59200
rect 90928 25566 90956 59191
rect 90916 25560 90968 25566
rect 90916 25502 90968 25508
rect 91560 11076 91612 11082
rect 91560 11018 91612 11024
rect 90732 7948 90784 7954
rect 90732 7890 90784 7896
rect 90364 4888 90416 4894
rect 90364 4830 90416 4836
rect 89628 3460 89680 3466
rect 89628 3402 89680 3408
rect 90376 480 90404 4830
rect 91572 480 91600 11018
rect 92400 8022 92428 59706
rect 97368 59702 97396 59735
rect 105634 59800 105636 59809
rect 110328 59832 110380 59838
rect 105688 59800 105690 59809
rect 101402 59735 101404 59744
rect 98644 59706 98696 59712
rect 101456 59735 101458 59744
rect 102784 59764 102836 59770
rect 101404 59706 101456 59712
rect 102784 59706 102836 59712
rect 105544 59764 105596 59770
rect 105634 59735 105690 59744
rect 107198 59800 107254 59809
rect 107198 59735 107254 59744
rect 108026 59800 108082 59809
rect 108026 59735 108028 59744
rect 105544 59706 105596 59712
rect 95884 59696 95936 59702
rect 95422 59664 95478 59673
rect 95884 59638 95936 59644
rect 97356 59696 97408 59702
rect 97356 59638 97408 59644
rect 97446 59664 97502 59673
rect 95422 59599 95478 59608
rect 93766 59528 93822 59537
rect 93766 59463 93822 59472
rect 93674 59392 93730 59401
rect 93674 59327 93730 59336
rect 93688 24138 93716 59327
rect 92480 24132 92532 24138
rect 92480 24074 92532 24080
rect 93676 24132 93728 24138
rect 93676 24074 93728 24080
rect 92388 8016 92440 8022
rect 92388 7958 92440 7964
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92492 354 92520 24074
rect 93780 9110 93808 59463
rect 95436 59401 95464 59599
rect 95422 59392 95478 59401
rect 95422 59327 95478 59336
rect 95146 59256 95202 59265
rect 95146 59191 95202 59200
rect 93858 59120 93914 59129
rect 93858 59055 93914 59064
rect 93768 9104 93820 9110
rect 93768 9046 93820 9052
rect 93872 7546 93900 59055
rect 95160 22574 95188 59191
rect 95148 22568 95200 22574
rect 95148 22510 95200 22516
rect 93952 15904 94004 15910
rect 93952 15846 94004 15852
rect 93860 7540 93912 7546
rect 93860 7482 93912 7488
rect 93964 480 93992 15846
rect 95792 13184 95844 13190
rect 95792 13126 95844 13132
rect 94780 7540 94832 7546
rect 94780 7482 94832 7488
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94792 354 94820 7482
rect 95118 354 95230 480
rect 94792 326 95230 354
rect 95804 354 95832 13126
rect 95896 11082 95924 59638
rect 97446 59599 97502 59608
rect 97354 59392 97410 59401
rect 97354 59327 97410 59336
rect 97368 45554 97396 59327
rect 97276 45526 97396 45554
rect 95884 11076 95936 11082
rect 95884 11018 95936 11024
rect 97276 10402 97304 45526
rect 97460 21486 97488 59599
rect 98000 22568 98052 22574
rect 98000 22510 98052 22516
rect 97448 21480 97500 21486
rect 97448 21422 97500 21428
rect 98012 16574 98040 22510
rect 98012 16546 98224 16574
rect 97264 10396 97316 10402
rect 97264 10338 97316 10344
rect 97448 5228 97500 5234
rect 97448 5170 97500 5176
rect 97460 480 97488 5170
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 98656 9042 98684 59706
rect 99746 59664 99802 59673
rect 99746 59599 99802 59608
rect 98826 59528 98882 59537
rect 98826 59463 98882 59472
rect 98840 18630 98868 59463
rect 99760 59401 99788 59599
rect 101586 59528 101642 59537
rect 101416 59486 101586 59514
rect 99746 59392 99802 59401
rect 99746 59327 99802 59336
rect 100022 59392 100078 59401
rect 100022 59327 100078 59336
rect 99380 28280 99432 28286
rect 99380 28222 99432 28228
rect 98828 18624 98880 18630
rect 98828 18566 98880 18572
rect 99392 16574 99420 28222
rect 99392 16546 99880 16574
rect 98644 9036 98696 9042
rect 98644 8978 98696 8984
rect 99852 480 99880 16546
rect 100036 15978 100064 59327
rect 100760 17332 100812 17338
rect 100760 17274 100812 17280
rect 100024 15972 100076 15978
rect 100024 15914 100076 15920
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 17274
rect 101416 6526 101444 59486
rect 101586 59463 101642 59472
rect 101586 59392 101642 59401
rect 101586 59327 101642 59336
rect 101600 17270 101628 59327
rect 101588 17264 101640 17270
rect 101588 17206 101640 17212
rect 102232 9104 102284 9110
rect 102232 9046 102284 9052
rect 101404 6520 101456 6526
rect 101404 6462 101456 6468
rect 102244 480 102272 9046
rect 102796 6390 102824 59706
rect 103978 59664 104034 59673
rect 103978 59599 104034 59608
rect 103150 59528 103206 59537
rect 103150 59463 103206 59472
rect 103164 45554 103192 59463
rect 103992 59401 104020 59599
rect 103978 59392 104034 59401
rect 103978 59327 104034 59336
rect 104162 59256 104218 59265
rect 104162 59191 104218 59200
rect 102980 45526 103192 45554
rect 102980 6458 103008 45526
rect 103520 18624 103572 18630
rect 103520 18566 103572 18572
rect 103532 16574 103560 18566
rect 103532 16546 104112 16574
rect 102968 6452 103020 6458
rect 102968 6394 103020 6400
rect 102784 6384 102836 6390
rect 102784 6326 102836 6332
rect 103336 3256 103388 3262
rect 103336 3198 103388 3204
rect 103348 480 103376 3198
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 104176 6322 104204 59191
rect 104900 24132 104952 24138
rect 104900 24074 104952 24080
rect 104912 16574 104940 24074
rect 104912 16546 105492 16574
rect 104164 6316 104216 6322
rect 104164 6258 104216 6264
rect 105464 3482 105492 16546
rect 105556 6186 105584 59706
rect 107106 59664 107162 59673
rect 107106 59599 107162 59608
rect 105726 59528 105782 59537
rect 105726 59463 105782 59472
rect 105740 16574 105768 59463
rect 106922 59392 106978 59401
rect 106922 59327 106978 59336
rect 105740 16546 105860 16574
rect 105832 6254 105860 16546
rect 106936 7818 106964 59327
rect 107120 35222 107148 59599
rect 107212 59537 107240 59735
rect 108080 59735 108082 59744
rect 108854 59800 108910 59809
rect 111340 59832 111392 59838
rect 110328 59774 110380 59780
rect 111338 59800 111340 59809
rect 229468 59832 229520 59838
rect 111392 59800 111394 59809
rect 108854 59735 108910 59744
rect 108028 59706 108080 59712
rect 107198 59528 107254 59537
rect 107198 59463 107254 59472
rect 108302 59528 108358 59537
rect 108302 59463 108358 59472
rect 107108 35216 107160 35222
rect 107108 35158 107160 35164
rect 106924 7812 106976 7818
rect 106924 7754 106976 7760
rect 108316 7750 108344 59463
rect 108868 59401 108896 59735
rect 108854 59392 108910 59401
rect 108854 59327 108910 59336
rect 109682 59392 109738 59401
rect 109682 59327 109738 59336
rect 109316 8016 109368 8022
rect 109316 7958 109368 7964
rect 108304 7744 108356 7750
rect 108304 7686 108356 7692
rect 105820 6248 105872 6254
rect 105820 6190 105872 6196
rect 105544 6180 105596 6186
rect 105544 6122 105596 6128
rect 108120 6180 108172 6186
rect 108120 6122 108172 6128
rect 106924 4140 106976 4146
rect 106924 4082 106976 4088
rect 105464 3454 105768 3482
rect 105740 480 105768 3454
rect 106936 480 106964 4082
rect 108132 480 108160 6122
rect 109328 480 109356 7958
rect 109696 7682 109724 59327
rect 110340 57322 110368 59774
rect 111064 59764 111116 59770
rect 111338 59735 111394 59744
rect 113730 59800 113786 59809
rect 116214 59800 116270 59809
rect 113730 59735 113732 59744
rect 111064 59706 111116 59712
rect 113784 59735 113786 59744
rect 114008 59764 114060 59770
rect 113732 59706 113784 59712
rect 122010 59800 122066 59809
rect 116214 59735 116216 59744
rect 114008 59706 114060 59712
rect 116268 59735 116270 59744
rect 119528 59764 119580 59770
rect 116216 59706 116268 59712
rect 122010 59735 122012 59744
rect 119528 59706 119580 59712
rect 122064 59735 122066 59744
rect 123114 59800 123170 59809
rect 126426 59800 126482 59809
rect 123114 59735 123170 59744
rect 124864 59764 124916 59770
rect 122012 59706 122064 59712
rect 110328 57316 110380 57322
rect 110328 57258 110380 57264
rect 110512 54596 110564 54602
rect 110512 54538 110564 54544
rect 109684 7676 109736 7682
rect 109684 7618 109736 7624
rect 110524 6914 110552 54538
rect 111076 7614 111104 59706
rect 111338 59664 111394 59673
rect 111338 59599 111394 59608
rect 111246 59528 111302 59537
rect 111246 59463 111302 59472
rect 111260 37942 111288 59463
rect 111352 59401 111380 59599
rect 113822 59528 113878 59537
rect 113822 59463 113878 59472
rect 111338 59392 111394 59401
rect 111338 59327 111394 59336
rect 112442 59392 112498 59401
rect 112442 59327 112498 59336
rect 111248 37936 111300 37942
rect 111248 37878 111300 37884
rect 112456 26926 112484 59327
rect 113836 39370 113864 59463
rect 114020 40730 114048 59706
rect 114190 59664 114246 59673
rect 117870 59664 117926 59673
rect 114190 59599 114246 59608
rect 117792 59622 117870 59650
rect 114204 59401 114232 59599
rect 117226 59528 117282 59537
rect 117226 59463 117282 59472
rect 114190 59392 114246 59401
rect 114190 59327 114246 59336
rect 115386 59392 115442 59401
rect 115386 59327 115442 59336
rect 115400 45554 115428 59327
rect 115846 59256 115902 59265
rect 115846 59191 115902 59200
rect 115216 45526 115428 45554
rect 115216 43450 115244 45526
rect 115204 43444 115256 43450
rect 115204 43386 115256 43392
rect 114008 40724 114060 40730
rect 114008 40666 114060 40672
rect 113824 39364 113876 39370
rect 113824 39306 113876 39312
rect 112444 26920 112496 26926
rect 112444 26862 112496 26868
rect 111800 25560 111852 25566
rect 111800 25502 111852 25508
rect 111812 16574 111840 25502
rect 111812 16546 112392 16574
rect 111064 7608 111116 7614
rect 111064 7550 111116 7556
rect 110524 6886 111656 6914
rect 110512 4004 110564 4010
rect 110512 3946 110564 3952
rect 110524 480 110552 3946
rect 111628 480 111656 6886
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114008 3868 114060 3874
rect 114008 3810 114060 3816
rect 114020 480 114048 3810
rect 115204 3596 115256 3602
rect 115204 3538 115256 3544
rect 115216 480 115244 3538
rect 115860 3330 115888 59191
rect 116400 7948 116452 7954
rect 116400 7890 116452 7896
rect 115848 3324 115900 3330
rect 115848 3266 115900 3272
rect 116412 480 116440 7890
rect 117240 3398 117268 59463
rect 117792 59401 117820 59622
rect 117870 59599 117926 59608
rect 118148 59628 118200 59634
rect 118148 59570 118200 59576
rect 117778 59392 117834 59401
rect 117778 59327 117834 59336
rect 117962 59392 118018 59401
rect 117962 59327 118018 59336
rect 117596 3732 117648 3738
rect 117596 3674 117648 3680
rect 117228 3392 117280 3398
rect 117228 3334 117280 3340
rect 117608 480 117636 3674
rect 117976 3602 118004 59327
rect 118160 54602 118188 59570
rect 119342 59256 119398 59265
rect 119342 59191 119398 59200
rect 118148 54596 118200 54602
rect 118148 54538 118200 54544
rect 119356 6186 119384 59191
rect 119540 18630 119568 59706
rect 120354 59664 120410 59673
rect 120354 59599 120356 59608
rect 120408 59599 120410 59608
rect 122286 59664 122342 59673
rect 122286 59599 122342 59608
rect 120356 59570 120408 59576
rect 122102 59528 122158 59537
rect 122102 59463 122158 59472
rect 120722 59392 120778 59401
rect 120722 59327 120778 59336
rect 119528 18624 119580 18630
rect 119528 18566 119580 18572
rect 120736 17338 120764 59327
rect 120724 17332 120776 17338
rect 120724 17274 120776 17280
rect 119896 7880 119948 7886
rect 119896 7822 119948 7828
rect 119344 6180 119396 6186
rect 119344 6122 119396 6128
rect 117964 3596 118016 3602
rect 117964 3538 118016 3544
rect 118792 3392 118844 3398
rect 118792 3334 118844 3340
rect 118804 480 118832 3334
rect 119908 480 119936 7822
rect 122116 5234 122144 59463
rect 122300 15910 122328 59599
rect 123128 59401 123156 59735
rect 130198 59800 130254 59809
rect 126426 59735 126428 59744
rect 124864 59706 124916 59712
rect 126480 59735 126482 59744
rect 127624 59764 127676 59770
rect 126428 59706 126480 59712
rect 131026 59800 131082 59809
rect 130198 59735 130200 59744
rect 127624 59706 127676 59712
rect 130252 59735 130254 59744
rect 130672 59758 131026 59786
rect 130200 59706 130252 59712
rect 123298 59664 123354 59673
rect 123298 59599 123354 59608
rect 123114 59392 123170 59401
rect 123312 59378 123340 59599
rect 123666 59392 123722 59401
rect 123312 59350 123666 59378
rect 123114 59327 123170 59336
rect 123666 59327 123722 59336
rect 123484 59288 123536 59294
rect 123484 59230 123536 59236
rect 123666 59256 123722 59265
rect 122288 15904 122340 15910
rect 122288 15846 122340 15852
rect 122104 5228 122156 5234
rect 122104 5170 122156 5176
rect 123496 5166 123524 59230
rect 123666 59191 123722 59200
rect 123484 5160 123536 5166
rect 123484 5102 123536 5108
rect 123680 4894 123708 59191
rect 124876 5098 124904 59706
rect 126242 59664 126298 59673
rect 126164 59622 126242 59650
rect 126164 59294 126192 59622
rect 126242 59599 126298 59608
rect 126426 59664 126482 59673
rect 126426 59599 126482 59608
rect 126242 59392 126298 59401
rect 126242 59327 126298 59336
rect 126152 59288 126204 59294
rect 126152 59230 126204 59236
rect 125600 22840 125652 22846
rect 125600 22782 125652 22788
rect 124864 5092 124916 5098
rect 124864 5034 124916 5040
rect 123668 4888 123720 4894
rect 123668 4830 123720 4836
rect 121092 3664 121144 3670
rect 121092 3606 121144 3612
rect 121104 480 121132 3606
rect 124680 3528 124732 3534
rect 124680 3470 124732 3476
rect 123484 3460 123536 3466
rect 123484 3402 123536 3408
rect 122288 3324 122340 3330
rect 122288 3266 122340 3272
rect 122300 480 122328 3266
rect 123496 480 123524 3402
rect 124692 480 124720 3470
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125612 354 125640 22782
rect 126256 13122 126284 59327
rect 126440 14482 126468 59599
rect 126980 54596 127032 54602
rect 126980 54538 127032 54544
rect 126428 14476 126480 14482
rect 126428 14418 126480 14424
rect 126244 13116 126296 13122
rect 126244 13058 126296 13064
rect 126992 480 127020 54538
rect 127532 14476 127584 14482
rect 127532 14418 127584 14424
rect 127544 3482 127572 14418
rect 127636 4962 127664 59706
rect 128542 59664 128598 59673
rect 128542 59599 128598 59608
rect 130568 59628 130620 59634
rect 127806 59528 127862 59537
rect 127806 59463 127862 59472
rect 127820 5030 127848 59463
rect 128556 59401 128584 59599
rect 130568 59570 130620 59576
rect 130382 59528 130438 59537
rect 130382 59463 130438 59472
rect 128542 59392 128598 59401
rect 128542 59327 128598 59336
rect 129002 59392 129058 59401
rect 129002 59327 129058 59336
rect 128360 26988 128412 26994
rect 128360 26930 128412 26936
rect 128372 16574 128400 26930
rect 128372 16546 128952 16574
rect 127808 5024 127860 5030
rect 127808 4966 127860 4972
rect 127624 4956 127676 4962
rect 127624 4898 127676 4904
rect 127544 3454 128216 3482
rect 128188 480 128216 3454
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 129016 11762 129044 59327
rect 129740 28484 129792 28490
rect 129740 28426 129792 28432
rect 129004 11756 129056 11762
rect 129004 11698 129056 11704
rect 129752 6914 129780 28426
rect 130396 8974 130424 59463
rect 130580 53106 130608 59570
rect 130672 59401 130700 59758
rect 131026 59735 131082 59744
rect 132038 59800 132094 59809
rect 132038 59735 132094 59744
rect 133142 59800 133198 59809
rect 133510 59800 133566 59809
rect 133198 59758 133510 59786
rect 133142 59735 133198 59744
rect 133510 59735 133566 59744
rect 134338 59800 134394 59809
rect 134338 59735 134394 59744
rect 135258 59800 135314 59809
rect 141698 59800 141754 59809
rect 135258 59735 135314 59744
rect 140688 59764 140740 59770
rect 131946 59664 132002 59673
rect 131946 59599 131948 59608
rect 132000 59599 132002 59608
rect 131948 59570 132000 59576
rect 130658 59392 130714 59401
rect 130658 59327 130714 59336
rect 131118 59392 131174 59401
rect 131118 59327 131174 59336
rect 131132 57254 131160 59327
rect 131120 57248 131172 57254
rect 131120 57190 131172 57196
rect 132052 55894 132080 59735
rect 133142 59528 133198 59537
rect 133142 59463 133198 59472
rect 132040 55888 132092 55894
rect 132040 55830 132092 55836
rect 130568 53100 130620 53106
rect 130568 53042 130620 53048
rect 133156 10334 133184 59463
rect 134352 59401 134380 59735
rect 135166 59664 135222 59673
rect 134536 59622 135166 59650
rect 134338 59392 134394 59401
rect 134338 59327 134394 59336
rect 134536 19990 134564 59622
rect 135166 59599 135222 59608
rect 135272 59537 135300 59735
rect 144458 59800 144514 59809
rect 141698 59735 141700 59744
rect 140688 59706 140740 59712
rect 141752 59735 141754 59744
rect 144196 59758 144458 59786
rect 141700 59706 141752 59712
rect 136822 59664 136878 59673
rect 136822 59599 136878 59608
rect 140044 59628 140096 59634
rect 135258 59528 135314 59537
rect 135258 59463 135314 59472
rect 135902 59528 135958 59537
rect 135902 59463 135958 59472
rect 134706 59256 134762 59265
rect 134706 59191 134762 59200
rect 134720 44878 134748 59191
rect 135916 46238 135944 59463
rect 136836 59401 136864 59599
rect 140044 59570 140096 59576
rect 139306 59528 139362 59537
rect 139306 59463 139362 59472
rect 139320 59430 139348 59463
rect 138112 59424 138164 59430
rect 136822 59392 136878 59401
rect 136822 59327 136878 59336
rect 137374 59392 137430 59401
rect 137374 59327 137430 59336
rect 138110 59392 138112 59401
rect 139308 59424 139360 59430
rect 138164 59392 138166 59401
rect 139308 59366 139360 59372
rect 138110 59327 138166 59336
rect 136086 59256 136142 59265
rect 136086 59191 136142 59200
rect 136100 54534 136128 59191
rect 136088 54528 136140 54534
rect 136088 54470 136140 54476
rect 137284 50380 137336 50386
rect 137284 50322 137336 50328
rect 136640 49156 136692 49162
rect 136640 49098 136692 49104
rect 135904 46232 135956 46238
rect 135904 46174 135956 46180
rect 134708 44872 134760 44878
rect 134708 44814 134760 44820
rect 134524 19984 134576 19990
rect 134524 19926 134576 19932
rect 136652 16574 136680 49098
rect 136652 16546 137232 16574
rect 135260 15904 135312 15910
rect 135260 15846 135312 15852
rect 133144 10328 133196 10334
rect 133144 10270 133196 10276
rect 130384 8968 130436 8974
rect 130384 8910 130436 8916
rect 131764 8968 131816 8974
rect 131764 8910 131816 8916
rect 129752 6886 130608 6914
rect 130580 480 130608 6886
rect 131776 480 131804 8910
rect 132960 7608 133012 7614
rect 132960 7550 133012 7556
rect 132972 480 133000 7550
rect 134156 6180 134208 6186
rect 134156 6122 134208 6128
rect 134168 480 134196 6122
rect 135272 480 135300 15846
rect 136456 3188 136508 3194
rect 136456 3130 136508 3136
rect 136468 480 136496 3130
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 137296 3194 137324 50322
rect 137388 49026 137416 59327
rect 138662 59256 138718 59265
rect 138662 59191 138718 59200
rect 137376 49020 137428 49026
rect 137376 48962 137428 48968
rect 138676 47598 138704 59191
rect 138846 59120 138902 59129
rect 138846 59055 138902 59064
rect 138860 50454 138888 59055
rect 138848 50448 138900 50454
rect 138848 50390 138900 50396
rect 138664 47592 138716 47598
rect 138664 47534 138716 47540
rect 139400 40724 139452 40730
rect 139400 40666 139452 40672
rect 139412 16574 139440 40666
rect 139412 16546 139624 16574
rect 137284 3188 137336 3194
rect 137284 3130 137336 3136
rect 138848 3188 138900 3194
rect 138848 3130 138900 3136
rect 138860 480 138888 3130
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 140056 4826 140084 59570
rect 140700 51746 140728 59706
rect 141698 59664 141754 59673
rect 141698 59599 141700 59608
rect 141752 59599 141754 59608
rect 141700 59570 141752 59576
rect 141514 59528 141570 59537
rect 141514 59463 141570 59472
rect 140688 51740 140740 51746
rect 140688 51682 140740 51688
rect 141424 36712 141476 36718
rect 141424 36654 141476 36660
rect 140044 4820 140096 4826
rect 140044 4762 140096 4768
rect 141240 4140 141292 4146
rect 141240 4082 141292 4088
rect 141252 480 141280 4082
rect 141436 3194 141464 36654
rect 141528 36582 141556 59463
rect 144196 59401 144224 59758
rect 144458 59735 144514 59744
rect 145838 59800 145894 59809
rect 145838 59735 145894 59744
rect 148690 59800 148746 59809
rect 151910 59800 151966 59809
rect 148690 59735 148746 59744
rect 150072 59764 150124 59770
rect 144550 59664 144606 59673
rect 144550 59599 144606 59608
rect 142894 59392 142950 59401
rect 142894 59327 142950 59336
rect 144182 59392 144238 59401
rect 144182 59327 144238 59336
rect 142066 59256 142122 59265
rect 142066 59191 142122 59200
rect 142080 58682 142108 59191
rect 142068 58676 142120 58682
rect 142068 58618 142120 58624
rect 142804 42220 142856 42226
rect 142804 42162 142856 42168
rect 141516 36576 141568 36582
rect 141516 36518 141568 36524
rect 142816 4146 142844 42162
rect 142908 42090 142936 59327
rect 143540 51808 143592 51814
rect 143540 51750 143592 51756
rect 142896 42084 142948 42090
rect 142896 42026 142948 42032
rect 142804 4140 142856 4146
rect 142804 4082 142856 4088
rect 142436 3664 142488 3670
rect 142436 3606 142488 3612
rect 141424 3188 141476 3194
rect 141424 3130 141476 3136
rect 142448 480 142476 3606
rect 143552 480 143580 51750
rect 144460 11824 144512 11830
rect 144460 11766 144512 11772
rect 144472 3482 144500 11766
rect 144564 3602 144592 59599
rect 145852 59537 145880 59735
rect 144734 59528 144790 59537
rect 144734 59463 144790 59472
rect 145838 59528 145894 59537
rect 145838 59463 145894 59472
rect 144748 16574 144776 59463
rect 146206 59392 146262 59401
rect 146206 59327 146262 59336
rect 144748 16546 144868 16574
rect 144552 3596 144604 3602
rect 144552 3538 144604 3544
rect 144472 3454 144776 3482
rect 144748 480 144776 3454
rect 144840 3369 144868 16546
rect 146220 3602 146248 59327
rect 148704 58954 148732 59735
rect 158166 59800 158222 59809
rect 151910 59735 151912 59744
rect 150072 59706 150124 59712
rect 151964 59735 151966 59744
rect 157156 59764 157208 59770
rect 151912 59706 151964 59712
rect 158166 59735 158168 59744
rect 157156 59706 157208 59712
rect 158220 59735 158222 59744
rect 164054 59800 164110 59809
rect 173346 59800 173402 59809
rect 164054 59735 164110 59744
rect 172428 59764 172480 59770
rect 158168 59706 158220 59712
rect 149978 59528 150034 59537
rect 149978 59463 150034 59472
rect 148874 59256 148930 59265
rect 148874 59191 148930 59200
rect 147588 58948 147640 58954
rect 147588 58890 147640 58896
rect 148692 58948 148744 58954
rect 148692 58890 148744 58896
rect 146300 53100 146352 53106
rect 146300 53042 146352 53048
rect 146312 16574 146340 53042
rect 146944 50448 146996 50454
rect 146944 50390 146996 50396
rect 146312 16546 146892 16574
rect 146208 3596 146260 3602
rect 146208 3538 146260 3544
rect 145932 3528 145984 3534
rect 145932 3470 145984 3476
rect 146864 3482 146892 16546
rect 146956 3670 146984 50390
rect 147600 26926 147628 58890
rect 148692 58404 148744 58410
rect 148692 58346 148744 58352
rect 147588 26920 147640 26926
rect 147588 26862 147640 26868
rect 148324 24268 148376 24274
rect 148324 24210 148376 24216
rect 147864 13116 147916 13122
rect 147864 13058 147916 13064
rect 146944 3664 146996 3670
rect 146944 3606 146996 3612
rect 144826 3360 144882 3369
rect 144826 3295 144882 3304
rect 145944 480 145972 3470
rect 146864 3454 147168 3482
rect 147140 480 147168 3454
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 147876 354 147904 13058
rect 148336 3534 148364 24210
rect 148704 18630 148732 58346
rect 148888 18698 148916 59191
rect 149992 58410 150020 59463
rect 149980 58404 150032 58410
rect 149980 58346 150032 58352
rect 150084 28286 150112 59706
rect 151634 59664 151690 59673
rect 150256 59628 150308 59634
rect 151634 59599 151636 59608
rect 150256 59570 150308 59576
rect 151688 59599 151690 59608
rect 152830 59664 152886 59673
rect 152830 59599 152886 59608
rect 154946 59664 155002 59673
rect 154946 59599 155002 59608
rect 151636 59570 151688 59576
rect 150268 33794 150296 59570
rect 151726 59528 151782 59537
rect 151726 59463 151782 59472
rect 150440 49020 150492 49026
rect 150440 48962 150492 48968
rect 150256 33788 150308 33794
rect 150256 33730 150308 33736
rect 150072 28280 150124 28286
rect 150072 28222 150124 28228
rect 148876 18692 148928 18698
rect 148876 18634 148928 18640
rect 148692 18624 148744 18630
rect 148692 18566 148744 18572
rect 150452 16574 150480 48962
rect 151740 18766 151768 59463
rect 152844 18834 152872 59599
rect 154302 59528 154358 59537
rect 154302 59463 154358 59472
rect 153014 59392 153070 59401
rect 153014 59327 153070 59336
rect 153028 18902 153056 59327
rect 154316 46238 154344 59463
rect 154960 59401 154988 59599
rect 156970 59528 157026 59537
rect 156970 59463 157026 59472
rect 154946 59392 155002 59401
rect 154946 59327 155002 59336
rect 155866 59392 155922 59401
rect 155866 59327 155922 59336
rect 154580 47728 154632 47734
rect 154580 47670 154632 47676
rect 154304 46232 154356 46238
rect 154304 46174 154356 46180
rect 153200 32496 153252 32502
rect 153200 32438 153252 32444
rect 153016 18896 153068 18902
rect 153016 18838 153068 18844
rect 152832 18828 152884 18834
rect 152832 18770 152884 18776
rect 151728 18760 151780 18766
rect 151728 18702 151780 18708
rect 153212 16574 153240 32438
rect 154592 16574 154620 47670
rect 155880 18970 155908 59327
rect 156984 22778 157012 59463
rect 157168 32434 157196 59706
rect 157246 59664 157302 59673
rect 157246 59599 157302 59608
rect 157614 59664 157670 59673
rect 157614 59599 157670 59608
rect 162766 59664 162822 59673
rect 162766 59599 162822 59608
rect 157260 58682 157288 59599
rect 157628 59401 157656 59599
rect 158350 59528 158406 59537
rect 158350 59463 158406 59472
rect 161202 59528 161258 59537
rect 161202 59463 161258 59472
rect 157614 59392 157670 59401
rect 157614 59327 157670 59336
rect 157248 58676 157300 58682
rect 157248 58618 157300 58624
rect 157340 33856 157392 33862
rect 157340 33798 157392 33804
rect 157156 32428 157208 32434
rect 157156 32370 157208 32376
rect 156972 22772 157024 22778
rect 156972 22714 157024 22720
rect 155868 18964 155920 18970
rect 155868 18906 155920 18912
rect 157352 16574 157380 33798
rect 158364 25566 158392 59463
rect 158626 59392 158682 59401
rect 158626 59327 158682 59336
rect 158640 51746 158668 59327
rect 158628 51740 158680 51746
rect 158628 51682 158680 51688
rect 158720 43648 158772 43654
rect 158720 43590 158772 43596
rect 158352 25560 158404 25566
rect 158352 25502 158404 25508
rect 158732 16574 158760 43590
rect 160100 29640 160152 29646
rect 160100 29582 160152 29588
rect 150452 16546 150664 16574
rect 153212 16546 153792 16574
rect 154592 16546 155448 16574
rect 157352 16546 157840 16574
rect 158732 16546 158944 16574
rect 148324 3528 148376 3534
rect 148324 3470 148376 3476
rect 149520 3528 149572 3534
rect 149520 3470 149572 3476
rect 149532 480 149560 3470
rect 150636 480 150664 16546
rect 151084 14544 151136 14550
rect 151084 14486 151136 14492
rect 151096 3534 151124 14486
rect 151820 13184 151872 13190
rect 151820 13126 151872 13132
rect 151084 3528 151136 3534
rect 151084 3470 151136 3476
rect 151832 480 151860 13126
rect 153016 11960 153068 11966
rect 153016 11902 153068 11908
rect 153028 480 153056 11902
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16546
rect 155420 480 155448 16546
rect 156604 3324 156656 3330
rect 156604 3266 156656 3272
rect 156616 480 156644 3266
rect 157812 480 157840 16546
rect 158916 480 158944 16546
rect 160112 3534 160140 29582
rect 161216 24138 161244 59463
rect 162490 59392 162546 59401
rect 162490 59327 162546 59336
rect 161480 46368 161532 46374
rect 161480 46310 161532 46316
rect 161204 24132 161256 24138
rect 161204 24074 161256 24080
rect 161492 16574 161520 46310
rect 162504 35222 162532 59327
rect 162674 59256 162730 59265
rect 162674 59191 162730 59200
rect 162688 37942 162716 59191
rect 162780 55894 162808 59599
rect 162860 58812 162912 58818
rect 162860 58754 162912 58760
rect 162768 55888 162820 55894
rect 162768 55830 162820 55836
rect 162676 37936 162728 37942
rect 162676 37878 162728 37884
rect 162492 35216 162544 35222
rect 162492 35158 162544 35164
rect 162872 16574 162900 58754
rect 164068 57254 164096 59735
rect 183742 59800 183798 59809
rect 173346 59735 173348 59744
rect 172428 59706 172480 59712
rect 173400 59735 173402 59744
rect 182088 59764 182140 59770
rect 173348 59706 173400 59712
rect 183742 59735 183744 59744
rect 182088 59706 182140 59712
rect 183796 59735 183798 59744
rect 185398 59800 185454 59809
rect 185398 59735 185454 59744
rect 186226 59800 186282 59809
rect 194414 59800 194470 59809
rect 186226 59735 186282 59744
rect 192852 59764 192904 59770
rect 183744 59706 183796 59712
rect 164790 59664 164846 59673
rect 166446 59664 166502 59673
rect 164790 59599 164846 59608
rect 165436 59628 165488 59634
rect 164146 59528 164202 59537
rect 164146 59463 164202 59472
rect 164056 57248 164108 57254
rect 164056 57190 164108 57196
rect 164160 17270 164188 59463
rect 164804 59401 164832 59599
rect 166446 59599 166448 59608
rect 165436 59570 165488 59576
rect 166500 59599 166502 59608
rect 167274 59664 167330 59673
rect 167274 59599 167330 59608
rect 166448 59570 166500 59576
rect 164790 59392 164846 59401
rect 164790 59327 164846 59336
rect 165250 59392 165306 59401
rect 165250 59327 165306 59336
rect 164240 35352 164292 35358
rect 164240 35294 164292 35300
rect 164148 17264 164200 17270
rect 164148 17206 164200 17212
rect 164252 16574 164280 35294
rect 165264 17406 165292 59327
rect 165252 17400 165304 17406
rect 165252 17342 165304 17348
rect 165448 17338 165476 59570
rect 166814 59528 166870 59537
rect 166632 59492 166684 59498
rect 166814 59463 166870 59472
rect 166632 59434 166684 59440
rect 165620 44940 165672 44946
rect 165620 44882 165672 44888
rect 165436 17332 165488 17338
rect 165436 17274 165488 17280
rect 165632 16574 165660 44882
rect 166644 17542 166672 59434
rect 166632 17536 166684 17542
rect 166632 17478 166684 17484
rect 166828 17474 166856 59463
rect 167288 59401 167316 59599
rect 168930 59528 168986 59537
rect 171414 59528 171470 59537
rect 168930 59463 168932 59472
rect 168984 59463 168986 59472
rect 169392 59492 169444 59498
rect 168932 59434 168984 59440
rect 171414 59463 171416 59472
rect 169392 59434 169444 59440
rect 171468 59463 171470 59472
rect 171416 59434 171468 59440
rect 167274 59392 167330 59401
rect 167274 59327 167330 59336
rect 168286 59392 168342 59401
rect 168286 59327 168342 59336
rect 168300 17610 168328 59327
rect 168380 47864 168432 47870
rect 168380 47806 168432 47812
rect 168288 17604 168340 17610
rect 168288 17546 168340 17552
rect 166816 17468 166868 17474
rect 166816 17410 166868 17416
rect 161492 16546 162072 16574
rect 162872 16546 163728 16574
rect 164252 16546 164464 16574
rect 165632 16546 166120 16574
rect 160100 3528 160152 3534
rect 160100 3470 160152 3476
rect 161296 3528 161348 3534
rect 161296 3470 161348 3476
rect 160100 3256 160152 3262
rect 160100 3198 160152 3204
rect 160112 480 160140 3198
rect 161308 480 161336 3470
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 16546
rect 163700 480 163728 16546
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164436 354 164464 16546
rect 166092 480 166120 16546
rect 168392 11762 168420 47806
rect 168472 38004 168524 38010
rect 168472 37946 168524 37952
rect 168380 11756 168432 11762
rect 168380 11698 168432 11704
rect 168484 6914 168512 37946
rect 169404 17746 169432 59434
rect 170770 59392 170826 59401
rect 170770 59327 170826 59336
rect 169574 59256 169630 59265
rect 169574 59191 169630 59200
rect 169392 17740 169444 17746
rect 169392 17682 169444 17688
rect 169588 17678 169616 59191
rect 169576 17672 169628 17678
rect 169576 17614 169628 17620
rect 170784 16574 170812 59327
rect 170954 59120 171010 59129
rect 170954 59055 171010 59064
rect 170784 16546 170904 16574
rect 169576 11756 169628 11762
rect 169576 11698 169628 11704
rect 168392 6886 168512 6914
rect 167184 6588 167236 6594
rect 167184 6530 167236 6536
rect 167196 480 167224 6530
rect 168392 480 168420 6886
rect 169588 480 169616 11698
rect 170772 7948 170824 7954
rect 170772 7890 170824 7896
rect 170784 480 170812 7890
rect 170876 3534 170904 16546
rect 170968 3670 170996 59055
rect 171140 39364 171192 39370
rect 171140 39306 171192 39312
rect 171152 16574 171180 39306
rect 171152 16546 172008 16574
rect 170956 3664 171008 3670
rect 170956 3606 171008 3612
rect 170864 3528 170916 3534
rect 170864 3470 170916 3476
rect 171980 480 172008 16546
rect 172440 3738 172468 59706
rect 173530 59664 173586 59673
rect 175462 59664 175518 59673
rect 173530 59599 173586 59608
rect 174912 59628 174964 59634
rect 172520 56160 172572 56166
rect 172520 56102 172572 56108
rect 172532 16574 172560 56102
rect 172532 16546 172744 16574
rect 172428 3732 172480 3738
rect 172428 3674 172480 3680
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 173544 3806 173572 59599
rect 175462 59599 175518 59608
rect 177118 59664 177174 59673
rect 177118 59599 177120 59608
rect 174912 59570 174964 59576
rect 173714 59392 173770 59401
rect 173714 59327 173770 59336
rect 173728 3874 173756 59327
rect 174268 6656 174320 6662
rect 174268 6598 174320 6604
rect 173716 3868 173768 3874
rect 173716 3810 173768 3816
rect 173532 3800 173584 3806
rect 173532 3742 173584 3748
rect 174280 480 174308 6598
rect 174924 4010 174952 59570
rect 175094 59528 175150 59537
rect 175094 59463 175150 59472
rect 174912 4004 174964 4010
rect 174912 3946 174964 3952
rect 175108 3942 175136 59463
rect 175476 59401 175504 59599
rect 177172 59599 177174 59608
rect 177946 59664 178002 59673
rect 177946 59599 178002 59608
rect 177120 59570 177172 59576
rect 177670 59528 177726 59537
rect 177670 59463 177726 59472
rect 175462 59392 175518 59401
rect 175462 59327 175518 59336
rect 176566 59392 176622 59401
rect 176566 59327 176622 59336
rect 175280 43512 175332 43518
rect 175280 43454 175332 43460
rect 175292 16574 175320 43454
rect 175292 16546 175504 16574
rect 175096 3936 175148 3942
rect 175096 3878 175148 3884
rect 175476 480 175504 16546
rect 176580 4078 176608 59327
rect 176660 36780 176712 36786
rect 176660 36722 176712 36728
rect 176568 4072 176620 4078
rect 176568 4014 176620 4020
rect 176672 480 176700 36722
rect 177580 15972 177632 15978
rect 177580 15914 177632 15920
rect 177592 3482 177620 15914
rect 177684 4146 177712 59463
rect 177960 59401 177988 59599
rect 180430 59528 180486 59537
rect 179328 59492 179380 59498
rect 180430 59463 180432 59472
rect 179328 59434 179380 59440
rect 180484 59463 180486 59472
rect 180432 59434 180484 59440
rect 177946 59392 178002 59401
rect 177946 59327 178002 59336
rect 177854 59256 177910 59265
rect 177854 59191 177910 59200
rect 179142 59256 179198 59265
rect 179142 59191 179198 59200
rect 177868 16574 177896 59191
rect 178040 40792 178092 40798
rect 178040 40734 178092 40740
rect 178052 16574 178080 40734
rect 179156 32570 179184 59191
rect 179144 32564 179196 32570
rect 179144 32506 179196 32512
rect 179340 21418 179368 59434
rect 180706 59392 180762 59401
rect 181074 59392 181130 59401
rect 180706 59327 180762 59336
rect 180812 59350 181074 59378
rect 179420 31204 179472 31210
rect 179420 31146 179472 31152
rect 179328 21412 179380 21418
rect 179328 21354 179380 21360
rect 179432 16574 179460 31146
rect 180720 21486 180748 59327
rect 180812 59265 180840 59350
rect 181074 59327 181130 59336
rect 180798 59256 180854 59265
rect 180798 59191 180854 59200
rect 181994 59120 182050 59129
rect 181994 59055 182050 59064
rect 180800 54528 180852 54534
rect 180800 54470 180852 54476
rect 180708 21480 180760 21486
rect 180708 21422 180760 21428
rect 180812 16574 180840 54470
rect 182008 43586 182036 59055
rect 181996 43580 182048 43586
rect 181996 43522 182048 43528
rect 182100 21554 182128 59706
rect 184846 59528 184902 59537
rect 184846 59463 184902 59472
rect 183190 59256 183246 59265
rect 183190 59191 183246 59200
rect 182180 42084 182232 42090
rect 182180 42026 182232 42032
rect 182088 21548 182140 21554
rect 182088 21490 182140 21496
rect 177868 16546 177988 16574
rect 178052 16546 178632 16574
rect 179432 16546 180288 16574
rect 180812 16546 181024 16574
rect 177672 4140 177724 4146
rect 177672 4082 177724 4088
rect 177592 3454 177896 3482
rect 177868 480 177896 3454
rect 177960 3398 177988 16546
rect 177948 3392 178000 3398
rect 177948 3334 178000 3340
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173134 -960 173246 326
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 180260 480 180288 16546
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 42026
rect 183204 11694 183232 59191
rect 183374 59120 183430 59129
rect 183374 59055 183430 59064
rect 183388 51882 183416 59055
rect 183376 51876 183428 51882
rect 183376 51818 183428 51824
rect 184860 29782 184888 59463
rect 185412 59401 185440 59735
rect 185950 59664 186006 59673
rect 185950 59599 186006 59608
rect 185398 59392 185454 59401
rect 185398 59327 185454 59336
rect 185964 47598 185992 59599
rect 186240 59537 186268 59735
rect 194414 59735 194416 59744
rect 192852 59706 192904 59712
rect 194468 59735 194470 59744
rect 195242 59800 195298 59809
rect 202786 59800 202842 59809
rect 195242 59735 195298 59744
rect 199844 59764 199896 59770
rect 194416 59706 194468 59712
rect 187882 59664 187938 59673
rect 187882 59599 187938 59608
rect 186226 59528 186282 59537
rect 186226 59463 186282 59472
rect 187330 59528 187386 59537
rect 187330 59463 187386 59472
rect 186134 59392 186190 59401
rect 186134 59327 186190 59336
rect 186148 49094 186176 59327
rect 186136 49088 186188 49094
rect 186136 49030 186188 49036
rect 185952 47592 186004 47598
rect 185952 47534 186004 47540
rect 184848 29776 184900 29782
rect 184848 29718 184900 29724
rect 187344 24342 187372 59463
rect 187896 59401 187924 59599
rect 190274 59528 190330 59537
rect 188896 59492 188948 59498
rect 190274 59463 190276 59472
rect 188896 59434 188948 59440
rect 190328 59463 190330 59472
rect 190552 59492 190604 59498
rect 190276 59434 190328 59440
rect 190552 59434 190604 59440
rect 188712 59424 188764 59430
rect 187882 59392 187938 59401
rect 188712 59366 188764 59372
rect 187882 59327 187938 59336
rect 187514 59256 187570 59265
rect 187514 59191 187570 59200
rect 187528 36650 187556 59191
rect 187516 36644 187568 36650
rect 187516 36586 187568 36592
rect 187332 24336 187384 24342
rect 187332 24278 187384 24284
rect 184940 24200 184992 24206
rect 184940 24142 184992 24148
rect 184952 11762 184980 24142
rect 188724 21622 188752 59366
rect 188908 27130 188936 59434
rect 190564 59401 190592 59434
rect 190550 59392 190606 59401
rect 190550 59327 190606 59336
rect 190366 59256 190422 59265
rect 190366 59191 190422 59200
rect 190380 57458 190408 59191
rect 191746 59120 191802 59129
rect 191746 59055 191802 59064
rect 190368 57452 190420 57458
rect 190368 57394 190420 57400
rect 188896 27124 188948 27130
rect 188896 27066 188948 27072
rect 189080 25628 189132 25634
rect 189080 25570 189132 25576
rect 188712 21616 188764 21622
rect 188712 21558 188764 21564
rect 189092 16574 189120 25570
rect 191760 19990 191788 59055
rect 192864 20126 192892 59706
rect 194506 59664 194562 59673
rect 194506 59599 194562 59608
rect 194414 59528 194470 59537
rect 194414 59463 194470 59472
rect 193034 59256 193090 59265
rect 193034 59191 193090 59200
rect 193048 40934 193076 59191
rect 193220 58744 193272 58750
rect 193220 58686 193272 58692
rect 193036 40928 193088 40934
rect 193036 40870 193088 40876
rect 192852 20120 192904 20126
rect 192852 20062 192904 20068
rect 191748 19984 191800 19990
rect 191748 19926 191800 19932
rect 189092 16546 189304 16574
rect 188528 16040 188580 16046
rect 188528 15982 188580 15988
rect 185032 14612 185084 14618
rect 185032 14554 185084 14560
rect 184940 11756 184992 11762
rect 184940 11698 184992 11704
rect 183192 11688 183244 11694
rect 183192 11630 183244 11636
rect 185044 6914 185072 14554
rect 186136 11756 186188 11762
rect 186136 11698 186188 11704
rect 184952 6886 185072 6914
rect 183744 4820 183796 4826
rect 183744 4762 183796 4768
rect 183756 480 183784 4762
rect 184952 480 184980 6886
rect 186148 480 186176 11698
rect 187332 4888 187384 4894
rect 187332 4830 187384 4836
rect 187344 480 187372 4830
rect 188540 480 188568 15982
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189276 354 189304 16546
rect 192024 6520 192076 6526
rect 192024 6462 192076 6468
rect 190828 4956 190880 4962
rect 190828 4898 190880 4904
rect 190840 480 190868 4898
rect 192036 480 192064 6462
rect 193232 480 193260 58686
rect 194428 56098 194456 59463
rect 194416 56092 194468 56098
rect 194416 56034 194468 56040
rect 194520 20194 194548 59599
rect 195256 59401 195284 59735
rect 199844 59706 199896 59712
rect 200212 59764 200264 59770
rect 200212 59706 200264 59712
rect 201316 59764 201368 59770
rect 209410 59800 209466 59809
rect 202786 59735 202788 59744
rect 201316 59706 201368 59712
rect 202840 59735 202842 59744
rect 208216 59764 208268 59770
rect 202788 59706 202840 59712
rect 209410 59735 209412 59744
rect 208216 59706 208268 59712
rect 209464 59735 209466 59744
rect 211710 59800 211766 59809
rect 215850 59800 215906 59809
rect 211710 59735 211766 59744
rect 213552 59764 213604 59770
rect 209412 59706 209464 59712
rect 195794 59664 195850 59673
rect 197082 59664 197138 59673
rect 195794 59599 195850 59608
rect 197004 59622 197082 59650
rect 195242 59392 195298 59401
rect 195242 59327 195298 59336
rect 195610 59392 195666 59401
rect 195610 59327 195666 59336
rect 195624 39574 195652 59327
rect 195808 42294 195836 59599
rect 197004 59401 197032 59622
rect 197082 59599 197138 59608
rect 197082 59528 197138 59537
rect 197082 59463 197138 59472
rect 196990 59392 197046 59401
rect 196990 59327 197046 59336
rect 195980 57316 196032 57322
rect 195980 57258 196032 57264
rect 195796 42288 195848 42294
rect 195796 42230 195848 42236
rect 195612 39568 195664 39574
rect 195612 39510 195664 39516
rect 194508 20188 194560 20194
rect 194508 20130 194560 20136
rect 195992 16574 196020 57258
rect 197096 53242 197124 59463
rect 197266 59392 197322 59401
rect 197266 59327 197322 59336
rect 197084 53236 197136 53242
rect 197084 53178 197136 53184
rect 197280 45014 197308 59327
rect 198646 59256 198702 59265
rect 198646 59191 198702 59200
rect 197268 45008 197320 45014
rect 197268 44950 197320 44956
rect 198660 25770 198688 59191
rect 199856 38146 199884 59706
rect 200224 59537 200252 59706
rect 201038 59664 201094 59673
rect 201038 59599 201094 59608
rect 200026 59528 200082 59537
rect 200026 59463 200082 59472
rect 200210 59528 200266 59537
rect 200210 59463 200266 59472
rect 199844 38140 199896 38146
rect 199844 38082 199896 38088
rect 198740 29844 198792 29850
rect 198740 29786 198792 29792
rect 198648 25764 198700 25770
rect 198648 25706 198700 25712
rect 195992 16546 196848 16574
rect 195612 7880 195664 7886
rect 195612 7822 195664 7828
rect 194416 5024 194468 5030
rect 194416 4966 194468 4972
rect 194428 480 194456 4966
rect 195624 480 195652 7822
rect 196820 480 196848 16546
rect 197912 5092 197964 5098
rect 197912 5034 197964 5040
rect 197924 480 197952 5034
rect 189694 354 189806 480
rect 189276 326 189806 354
rect 189694 -960 189806 326
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 29786
rect 200040 23050 200068 59463
rect 201052 59401 201080 59599
rect 201038 59392 201094 59401
rect 201038 59327 201094 59336
rect 201222 59392 201278 59401
rect 201222 59327 201278 59336
rect 201236 45554 201264 59327
rect 201144 45526 201264 45554
rect 200120 28348 200172 28354
rect 200120 28290 200172 28296
rect 200028 23044 200080 23050
rect 200028 22986 200080 22992
rect 200132 16574 200160 28290
rect 201144 20262 201172 45526
rect 201328 43790 201356 59706
rect 204166 59664 204222 59673
rect 204166 59599 204222 59608
rect 206098 59664 206154 59673
rect 206098 59599 206154 59608
rect 202786 59528 202842 59537
rect 202786 59463 202842 59472
rect 201316 43784 201368 43790
rect 201316 43726 201368 43732
rect 202800 31346 202828 59463
rect 203982 59392 204038 59401
rect 203982 59327 204038 59336
rect 203996 50658 204024 59327
rect 203984 50652 204036 50658
rect 203984 50594 204036 50600
rect 204180 47938 204208 59599
rect 205454 59528 205510 59537
rect 205272 59492 205324 59498
rect 205454 59463 205510 59472
rect 205272 59434 205324 59440
rect 204260 50516 204312 50522
rect 204260 50458 204312 50464
rect 204168 47932 204220 47938
rect 204168 47874 204220 47880
rect 202788 31340 202840 31346
rect 202788 31282 202840 31288
rect 202880 31068 202932 31074
rect 202880 31010 202932 31016
rect 201132 20256 201184 20262
rect 201132 20198 201184 20204
rect 202892 16574 202920 31010
rect 204272 16574 204300 50458
rect 205284 35494 205312 59434
rect 205468 54806 205496 59463
rect 206112 59401 206140 59599
rect 207570 59528 207626 59537
rect 207570 59463 207572 59472
rect 207624 59463 207626 59472
rect 207572 59434 207624 59440
rect 206098 59392 206154 59401
rect 206098 59327 206154 59336
rect 206926 59392 206982 59401
rect 206926 59327 206982 59336
rect 205456 54800 205508 54806
rect 205456 54742 205508 54748
rect 205640 53304 205692 53310
rect 205640 53246 205692 53252
rect 205272 35488 205324 35494
rect 205272 35430 205324 35436
rect 205652 16574 205680 53246
rect 206940 36854 206968 59327
rect 208030 59256 208086 59265
rect 208030 59191 208086 59200
rect 206928 36848 206980 36854
rect 206928 36790 206980 36796
rect 207020 32632 207072 32638
rect 207020 32574 207072 32580
rect 200132 16546 200344 16574
rect 202892 16546 203472 16574
rect 204272 16546 205128 16574
rect 205652 16546 206232 16574
rect 200316 480 200344 16546
rect 202696 6724 202748 6730
rect 202696 6666 202748 6672
rect 201500 5160 201552 5166
rect 201500 5102 201552 5108
rect 201512 480 201540 5102
rect 202708 480 202736 6666
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 16546
rect 205100 480 205128 16546
rect 206204 480 206232 16546
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 32574
rect 208044 29986 208072 59191
rect 208228 49366 208256 59706
rect 211066 59664 211122 59673
rect 211066 59599 211122 59608
rect 209410 59528 209466 59537
rect 209410 59463 209466 59472
rect 208216 49360 208268 49366
rect 208216 49302 208268 49308
rect 208032 29980 208084 29986
rect 208032 29922 208084 29928
rect 209424 11898 209452 59463
rect 209594 59256 209650 59265
rect 209594 59191 209650 59200
rect 209608 42430 209636 59191
rect 209780 55956 209832 55962
rect 209780 55898 209832 55904
rect 209596 42424 209648 42430
rect 209596 42366 209648 42372
rect 209412 11892 209464 11898
rect 209412 11834 209464 11840
rect 208584 5228 208636 5234
rect 208584 5170 208636 5176
rect 208596 480 208624 5170
rect 209792 4214 209820 55898
rect 211080 12034 211108 59599
rect 211724 59401 211752 59735
rect 215850 59735 215852 59744
rect 213552 59706 213604 59712
rect 215904 59735 215906 59744
rect 223210 59800 223266 59809
rect 229006 59800 229062 59809
rect 223210 59735 223266 59744
rect 228376 59758 229006 59786
rect 215852 59706 215904 59712
rect 212354 59528 212410 59537
rect 212354 59463 212410 59472
rect 211710 59392 211766 59401
rect 211710 59327 211766 59336
rect 212170 59392 212226 59401
rect 212170 59327 212226 59336
rect 211068 12028 211120 12034
rect 211068 11970 211120 11976
rect 212184 10402 212212 59327
rect 212172 10396 212224 10402
rect 212172 10338 212224 10344
rect 212368 10334 212396 59463
rect 212540 39500 212592 39506
rect 212540 39442 212592 39448
rect 212552 16574 212580 39442
rect 212552 16546 213408 16574
rect 212356 10328 212408 10334
rect 212356 10270 212408 10276
rect 209872 7812 209924 7818
rect 209872 7754 209924 7760
rect 209780 4208 209832 4214
rect 209780 4150 209832 4156
rect 209884 3482 209912 7754
rect 212172 5296 212224 5302
rect 212172 5238 212224 5244
rect 210976 4208 211028 4214
rect 210976 4150 211028 4156
rect 209792 3454 209912 3482
rect 209792 480 209820 3454
rect 210988 480 211016 4150
rect 212184 480 212212 5238
rect 213380 480 213408 16546
rect 213564 10538 213592 59706
rect 219162 59664 219218 59673
rect 217692 59628 217744 59634
rect 219162 59599 219164 59608
rect 217692 59570 217744 59576
rect 219216 59599 219218 59608
rect 219990 59664 220046 59673
rect 219990 59599 220046 59608
rect 219164 59570 219216 59576
rect 216494 59528 216550 59537
rect 216494 59463 216550 59472
rect 215206 59392 215262 59401
rect 215206 59327 215262 59336
rect 216310 59392 216366 59401
rect 216310 59327 216366 59336
rect 213734 59256 213790 59265
rect 213734 59191 213790 59200
rect 213552 10532 213604 10538
rect 213552 10474 213604 10480
rect 213748 10470 213776 59191
rect 213920 33924 213972 33930
rect 213920 33866 213972 33872
rect 213932 16574 213960 33866
rect 213932 16546 214512 16574
rect 213736 10464 213788 10470
rect 213736 10406 213788 10412
rect 214484 480 214512 16546
rect 215220 10606 215248 59327
rect 215300 27192 215352 27198
rect 215300 27134 215352 27140
rect 215208 10600 215260 10606
rect 215208 10542 215260 10548
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 27134
rect 216324 10674 216352 59327
rect 216508 39642 216536 59463
rect 216496 39636 216548 39642
rect 216496 39578 216548 39584
rect 216864 13252 216916 13258
rect 216864 13194 216916 13200
rect 216312 10668 216364 10674
rect 216312 10610 216364 10616
rect 216876 480 216904 13194
rect 217704 10742 217732 59570
rect 219346 59528 219402 59537
rect 219346 59463 219402 59472
rect 217874 59256 217930 59265
rect 217874 59191 217930 59200
rect 217888 45082 217916 59191
rect 217876 45076 217928 45082
rect 217876 45018 217928 45024
rect 218060 36576 218112 36582
rect 218060 36518 218112 36524
rect 217692 10736 217744 10742
rect 217692 10678 217744 10684
rect 218072 480 218100 36518
rect 219360 31142 219388 59463
rect 220004 59401 220032 59599
rect 222014 59528 222070 59537
rect 222014 59463 222070 59472
rect 219990 59392 220046 59401
rect 219990 59327 220046 59336
rect 221922 59392 221978 59401
rect 221922 59327 221978 59336
rect 220450 59256 220506 59265
rect 220450 59191 220506 59200
rect 219348 31136 219400 31142
rect 219348 31078 219400 31084
rect 220464 16114 220492 59191
rect 220634 59120 220690 59129
rect 220634 59055 220690 59064
rect 220648 29714 220676 59055
rect 221936 45554 221964 59327
rect 222028 53174 222056 59463
rect 223224 59401 223252 59735
rect 227628 59628 227680 59634
rect 227628 59570 227680 59576
rect 224866 59528 224922 59537
rect 226522 59528 226578 59537
rect 224866 59463 224922 59472
rect 225984 59486 226522 59514
rect 223210 59392 223266 59401
rect 223210 59327 223266 59336
rect 223486 59392 223542 59401
rect 223486 59327 223542 59336
rect 224774 59392 224830 59401
rect 224774 59327 224830 59336
rect 222016 53168 222068 53174
rect 222016 53110 222068 53116
rect 221844 45526 221964 45554
rect 220820 44872 220872 44878
rect 220820 44814 220872 44820
rect 220636 29708 220688 29714
rect 220636 29650 220688 29656
rect 220832 16574 220860 44814
rect 221844 39438 221872 45526
rect 221832 39432 221884 39438
rect 221832 39374 221884 39380
rect 220832 16546 221136 16574
rect 220452 16108 220504 16114
rect 220452 16050 220504 16056
rect 220452 6792 220504 6798
rect 220452 6734 220504 6740
rect 219256 6248 219308 6254
rect 219256 6190 219308 6196
rect 219268 480 219296 6190
rect 220464 480 220492 6734
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221108 354 221136 16546
rect 223500 9042 223528 59327
rect 224788 9178 224816 59327
rect 224776 9172 224828 9178
rect 224776 9114 224828 9120
rect 224880 9110 224908 59463
rect 225984 59401 226012 59486
rect 226522 59463 226578 59472
rect 225970 59392 226026 59401
rect 225970 59327 226026 59336
rect 226154 59392 226210 59401
rect 226154 59327 226210 59336
rect 225970 59256 226026 59265
rect 225970 59191 226026 59200
rect 225984 53378 226012 59191
rect 226168 54670 226196 59327
rect 226156 54664 226208 54670
rect 226156 54606 226208 54612
rect 225972 53372 226024 53378
rect 225972 53314 226024 53320
rect 224960 46300 225012 46306
rect 224960 46242 225012 46248
rect 224972 16574 225000 46242
rect 224972 16546 225184 16574
rect 224868 9104 224920 9110
rect 224868 9046 224920 9052
rect 223488 9036 223540 9042
rect 223488 8978 223540 8984
rect 223948 8424 224000 8430
rect 223948 8366 224000 8372
rect 222752 6316 222804 6322
rect 222752 6258 222804 6264
rect 222764 480 222792 6258
rect 223960 480 223988 8366
rect 225156 480 225184 16546
rect 227640 9246 227668 59570
rect 227628 9240 227680 9246
rect 227628 9182 227680 9188
rect 228376 8226 228404 59758
rect 229006 59735 229062 59744
rect 229466 59800 229468 59809
rect 230664 59832 230716 59838
rect 229520 59800 229522 59809
rect 229466 59735 229522 59744
rect 230662 59800 230664 59809
rect 240508 59832 240560 59838
rect 230716 59800 230718 59809
rect 234802 59800 234858 59809
rect 230662 59735 230718 59744
rect 232504 59764 232556 59770
rect 234802 59735 234804 59744
rect 232504 59706 232556 59712
rect 234856 59735 234858 59744
rect 235630 59800 235686 59809
rect 238850 59800 238906 59809
rect 235630 59735 235686 59744
rect 238024 59764 238076 59770
rect 234804 59706 234856 59712
rect 229006 59664 229062 59673
rect 229006 59599 229008 59608
rect 229060 59599 229062 59608
rect 229008 59570 229060 59576
rect 229006 59528 229062 59537
rect 229006 59463 229062 59472
rect 229020 8362 229048 59463
rect 229926 59392 229982 59401
rect 229926 59327 229982 59336
rect 229742 59256 229798 59265
rect 229742 59191 229798 59200
rect 229008 8356 229060 8362
rect 229008 8298 229060 8304
rect 227536 8220 227588 8226
rect 227536 8162 227588 8168
rect 228364 8220 228416 8226
rect 228364 8162 228416 8168
rect 226340 6384 226392 6390
rect 226340 6326 226392 6332
rect 226352 480 226380 6326
rect 227548 480 227576 8162
rect 228732 7676 228784 7682
rect 228732 7618 228784 7624
rect 228744 480 228772 7618
rect 229756 6798 229784 59191
rect 229940 8430 229968 59327
rect 231122 59120 231178 59129
rect 231122 59055 231178 59064
rect 231136 13258 231164 59055
rect 231124 13252 231176 13258
rect 231124 13194 231176 13200
rect 229928 8424 229980 8430
rect 229928 8366 229980 8372
rect 231032 8356 231084 8362
rect 231032 8298 231084 8304
rect 229744 6792 229796 6798
rect 229744 6734 229796 6740
rect 229836 6452 229888 6458
rect 229836 6394 229888 6400
rect 229848 480 229876 6394
rect 231044 480 231072 8298
rect 232516 7818 232544 59706
rect 232686 59664 232742 59673
rect 232686 59599 232742 59608
rect 234802 59664 234858 59673
rect 234802 59599 234858 59608
rect 232700 39506 232728 59599
rect 234066 59528 234122 59537
rect 234066 59463 234122 59472
rect 233882 59392 233938 59401
rect 233882 59327 233938 59336
rect 233240 57520 233292 57526
rect 233240 57462 233292 57468
rect 232688 39500 232740 39506
rect 232688 39442 232740 39448
rect 233252 16574 233280 57462
rect 233252 16546 233464 16574
rect 232504 7812 232556 7818
rect 232504 7754 232556 7760
rect 232228 7744 232280 7750
rect 232228 7686 232280 7692
rect 232240 480 232268 7686
rect 233436 480 233464 16546
rect 233896 6730 233924 59327
rect 234080 53310 234108 59463
rect 234816 59401 234844 59599
rect 235644 59537 235672 59735
rect 240506 59800 240508 59809
rect 296996 59832 297048 59838
rect 240560 59800 240562 59809
rect 238850 59735 238906 59744
rect 239404 59764 239456 59770
rect 238024 59706 238076 59712
rect 236644 59696 236696 59702
rect 236644 59638 236696 59644
rect 235630 59528 235686 59537
rect 235630 59463 235686 59472
rect 234802 59392 234858 59401
rect 234802 59327 234858 59336
rect 235446 59392 235502 59401
rect 235446 59327 235502 59336
rect 235262 59256 235318 59265
rect 235262 59191 235318 59200
rect 234068 53304 234120 53310
rect 234068 53246 234120 53252
rect 234620 9240 234672 9246
rect 234620 9182 234672 9188
rect 233884 6724 233936 6730
rect 233884 6666 233936 6672
rect 234632 480 234660 9182
rect 235276 7886 235304 59191
rect 235460 29850 235488 59327
rect 236000 52012 236052 52018
rect 236000 51954 236052 51960
rect 235448 29844 235500 29850
rect 235448 29786 235500 29792
rect 236012 16574 236040 51954
rect 236012 16546 236592 16574
rect 235264 7880 235316 7886
rect 235264 7822 235316 7828
rect 235816 7812 235868 7818
rect 235816 7754 235868 7760
rect 235828 480 235856 7754
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 236656 6526 236684 59638
rect 237380 53372 237432 53378
rect 237380 53314 237432 53320
rect 237392 16574 237420 53314
rect 237392 16546 237696 16574
rect 236644 6520 236696 6526
rect 236644 6462 236696 6468
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 16546
rect 238036 14618 238064 59706
rect 238864 59702 238892 59735
rect 240506 59735 240562 59744
rect 242162 59800 242218 59809
rect 245474 59800 245530 59809
rect 242162 59735 242164 59744
rect 239404 59706 239456 59712
rect 242216 59735 242218 59744
rect 244188 59764 244240 59770
rect 242164 59706 242216 59712
rect 250534 59800 250590 59809
rect 245474 59735 245476 59744
rect 244188 59706 244240 59712
rect 245528 59735 245530 59744
rect 249064 59764 249116 59770
rect 245476 59706 245528 59712
rect 250534 59735 250590 59744
rect 251270 59800 251326 59809
rect 252282 59800 252338 59809
rect 251270 59735 251272 59744
rect 249064 59706 249116 59712
rect 238852 59696 238904 59702
rect 238852 59638 238904 59644
rect 238298 59528 238354 59537
rect 238298 59463 238354 59472
rect 238312 45554 238340 59463
rect 238220 45526 238340 45554
rect 238220 16046 238248 45526
rect 238208 16040 238260 16046
rect 238208 15982 238260 15988
rect 239416 15978 239444 59706
rect 242346 59528 242402 59537
rect 242346 59463 242402 59472
rect 239586 59392 239642 59401
rect 239586 59327 239642 59336
rect 239600 54534 239628 59327
rect 240782 59256 240838 59265
rect 240782 59191 240838 59200
rect 239588 54528 239640 54534
rect 239588 54470 239640 54476
rect 239404 15972 239456 15978
rect 239404 15914 239456 15920
rect 238024 14612 238076 14618
rect 238024 14554 238076 14560
rect 239312 7880 239364 7886
rect 239312 7822 239364 7828
rect 239324 480 239352 7822
rect 240796 6662 240824 59191
rect 242162 59120 242218 59129
rect 242162 59055 242218 59064
rect 241520 54664 241572 54670
rect 241520 54606 241572 54612
rect 241532 16574 241560 54606
rect 241532 16546 241744 16574
rect 240784 6656 240836 6662
rect 240784 6598 240836 6604
rect 240508 6520 240560 6526
rect 240508 6462 240560 6468
rect 240520 480 240548 6462
rect 241716 480 241744 16546
rect 242176 6594 242204 59055
rect 242360 7954 242388 59463
rect 243542 59256 243598 59265
rect 243542 59191 243598 59200
rect 242900 47796 242952 47802
rect 242900 47738 242952 47744
rect 242348 7948 242400 7954
rect 242348 7890 242400 7896
rect 242164 6588 242216 6594
rect 242164 6530 242216 6536
rect 242912 480 242940 47738
rect 242992 25900 243044 25906
rect 242992 25842 243044 25848
rect 243004 16574 243032 25842
rect 243004 16546 243492 16574
rect 243464 3074 243492 16546
rect 243556 3262 243584 59191
rect 244200 58818 244228 59706
rect 245474 59664 245530 59673
rect 248878 59664 248934 59673
rect 245474 59599 245530 59608
rect 246488 59628 246540 59634
rect 244922 59528 244978 59537
rect 244922 59463 244978 59472
rect 244188 58812 244240 58818
rect 244188 58754 244240 58760
rect 244936 3330 244964 59463
rect 245488 59401 245516 59599
rect 248878 59599 248880 59608
rect 246488 59570 246540 59576
rect 248932 59599 248934 59608
rect 248880 59570 248932 59576
rect 246304 59492 246356 59498
rect 246304 59434 246356 59440
rect 245474 59392 245530 59401
rect 245474 59327 245530 59336
rect 246316 11966 246344 59434
rect 246500 14550 246528 59570
rect 247868 59560 247920 59566
rect 247868 59502 247920 59508
rect 247958 59528 248014 59537
rect 247682 59392 247738 59401
rect 247682 59327 247738 59336
rect 247696 24274 247724 59327
rect 247880 50454 247908 59502
rect 247958 59463 247960 59472
rect 248012 59463 248014 59472
rect 247960 59434 248012 59440
rect 247868 50448 247920 50454
rect 247868 50390 247920 50396
rect 249076 36718 249104 59706
rect 249614 59664 249670 59673
rect 249614 59599 249670 59608
rect 249628 59401 249656 59599
rect 250548 59566 250576 59735
rect 251324 59735 251326 59744
rect 252020 59758 252282 59786
rect 251272 59706 251324 59712
rect 250626 59664 250682 59673
rect 250626 59599 250682 59608
rect 250536 59560 250588 59566
rect 250442 59528 250498 59537
rect 250536 59502 250588 59508
rect 250442 59463 250498 59472
rect 249614 59392 249670 59401
rect 249614 59327 249670 59336
rect 249064 36712 249116 36718
rect 249064 36654 249116 36660
rect 247684 24268 247736 24274
rect 247684 24210 247736 24216
rect 246488 14544 246540 14550
rect 246488 14486 246540 14492
rect 246304 11960 246356 11966
rect 246304 11902 246356 11908
rect 245200 9172 245252 9178
rect 245200 9114 245252 9120
rect 244924 3324 244976 3330
rect 244924 3266 244976 3272
rect 243544 3256 243596 3262
rect 243544 3198 243596 3204
rect 243464 3046 244136 3074
rect 244108 480 244136 3046
rect 245212 480 245240 9114
rect 248788 9104 248840 9110
rect 248788 9046 248840 9052
rect 246396 7948 246448 7954
rect 246396 7890 246448 7896
rect 246408 480 246436 7890
rect 247592 6588 247644 6594
rect 247592 6530 247644 6536
rect 247604 480 247632 6530
rect 248800 480 248828 9046
rect 250456 8974 250484 59463
rect 250640 15910 250668 59599
rect 252020 59537 252048 59758
rect 252282 59735 252338 59744
rect 254582 59800 254638 59809
rect 254582 59735 254638 59744
rect 267462 59800 267518 59809
rect 267462 59735 267464 59744
rect 252006 59528 252062 59537
rect 252006 59463 252062 59472
rect 252282 59528 252338 59537
rect 252282 59463 252338 59472
rect 251180 58948 251232 58954
rect 251180 58890 251232 58896
rect 250628 15904 250680 15910
rect 250628 15846 250680 15852
rect 250444 8968 250496 8974
rect 250444 8910 250496 8916
rect 249984 8016 250036 8022
rect 249984 7958 250036 7964
rect 249996 480 250024 7958
rect 251192 480 251220 58890
rect 252296 45554 252324 59463
rect 254596 59401 254624 59735
rect 267516 59735 267518 59744
rect 269854 59800 269910 59809
rect 270682 59800 270738 59809
rect 269854 59735 269910 59744
rect 269948 59764 270000 59770
rect 267464 59706 267516 59712
rect 269868 59702 269896 59735
rect 278042 59800 278098 59809
rect 270682 59735 270684 59744
rect 269948 59706 270000 59712
rect 270736 59735 270738 59744
rect 271880 59764 271932 59770
rect 270684 59706 270736 59712
rect 271880 59706 271932 59712
rect 277216 59764 277268 59770
rect 277216 59706 277268 59712
rect 277860 59764 277912 59770
rect 278042 59735 278098 59744
rect 278870 59800 278926 59809
rect 278870 59735 278926 59744
rect 281354 59800 281410 59809
rect 283010 59800 283066 59809
rect 281410 59758 281764 59786
rect 281354 59735 281410 59744
rect 277860 59706 277912 59712
rect 269856 59696 269908 59702
rect 257802 59664 257858 59673
rect 256332 59628 256384 59634
rect 257802 59599 257804 59608
rect 256332 59570 256384 59576
rect 257856 59599 257858 59608
rect 258630 59664 258686 59673
rect 261114 59664 261170 59673
rect 258630 59599 258686 59608
rect 259092 59628 259144 59634
rect 257804 59570 257856 59576
rect 255134 59528 255190 59537
rect 255134 59463 255190 59472
rect 254582 59392 254638 59401
rect 254582 59327 254638 59336
rect 254950 59392 255006 59401
rect 254950 59327 255006 59336
rect 252466 59256 252522 59265
rect 252466 59191 252522 59200
rect 253846 59256 253902 59265
rect 253846 59191 253902 59200
rect 251836 45526 252324 45554
rect 251836 14482 251864 45526
rect 252480 22914 252508 59191
rect 252560 54664 252612 54670
rect 252560 54606 252612 54612
rect 252468 22908 252520 22914
rect 252468 22850 252520 22856
rect 252572 16574 252600 54606
rect 253860 54534 253888 59191
rect 253848 54528 253900 54534
rect 253848 54470 253900 54476
rect 253940 41064 253992 41070
rect 253940 41006 253992 41012
rect 253952 16574 253980 41006
rect 254964 35290 254992 59327
rect 255148 43450 255176 59463
rect 255320 53168 255372 53174
rect 255320 53110 255372 53116
rect 255136 43444 255188 43450
rect 255136 43386 255188 43392
rect 254952 35284 255004 35290
rect 254952 35226 255004 35232
rect 255332 16574 255360 53110
rect 252572 16546 253520 16574
rect 253952 16546 254256 16574
rect 255332 16546 255912 16574
rect 251824 14476 251876 14482
rect 251824 14418 251876 14424
rect 252376 9036 252428 9042
rect 252376 8978 252428 8984
rect 252388 480 252416 8978
rect 253492 480 253520 16546
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 255884 480 255912 16546
rect 256344 14482 256372 59570
rect 257986 59528 258042 59537
rect 257986 59463 258042 59472
rect 256514 59256 256570 59265
rect 256514 59191 256570 59200
rect 256528 14550 256556 59191
rect 256700 49224 256752 49230
rect 256700 49166 256752 49172
rect 256516 14544 256568 14550
rect 256516 14486 256568 14492
rect 256332 14476 256384 14482
rect 256332 14418 256384 14424
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 256712 354 256740 49166
rect 258000 14618 258028 59463
rect 258644 59401 258672 59599
rect 261114 59599 261116 59608
rect 259092 59570 259144 59576
rect 261168 59599 261170 59608
rect 265714 59664 265770 59673
rect 269856 59638 269908 59644
rect 265714 59599 265770 59608
rect 261116 59570 261168 59576
rect 258630 59392 258686 59401
rect 258630 59327 258686 59336
rect 258080 53372 258132 53378
rect 258080 53314 258132 53320
rect 258092 16574 258120 53314
rect 258092 16546 258304 16574
rect 257988 14612 258040 14618
rect 257988 14554 258040 14560
rect 258276 480 258304 16546
rect 259104 14754 259132 59570
rect 260746 59528 260802 59537
rect 260746 59463 260802 59472
rect 259274 59256 259330 59265
rect 259274 59191 259330 59200
rect 259092 14748 259144 14754
rect 259092 14690 259144 14696
rect 259288 14686 259316 59191
rect 259460 53168 259512 53174
rect 259460 53110 259512 53116
rect 259276 14680 259328 14686
rect 259276 14622 259328 14628
rect 259472 11694 259500 53110
rect 259552 39432 259604 39438
rect 259552 39374 259604 39380
rect 259460 11688 259512 11694
rect 259460 11630 259512 11636
rect 259564 6914 259592 39374
rect 260760 14822 260788 59463
rect 265728 59401 265756 59599
rect 267002 59528 267058 59537
rect 267002 59463 267058 59472
rect 269762 59528 269818 59537
rect 269762 59463 269818 59472
rect 265530 59392 265586 59401
rect 265530 59327 265586 59336
rect 265714 59392 265770 59401
rect 265714 59327 265770 59336
rect 263600 51944 263652 51950
rect 263600 51886 263652 51892
rect 260840 32700 260892 32706
rect 260840 32642 260892 32648
rect 260852 16574 260880 32642
rect 262220 29708 262272 29714
rect 262220 29650 262272 29656
rect 262232 16574 262260 29650
rect 263612 16574 263640 51886
rect 265544 51074 265572 59327
rect 265544 51046 265664 51074
rect 264980 24472 265032 24478
rect 264980 24414 265032 24420
rect 260852 16546 261800 16574
rect 262232 16546 262536 16574
rect 263612 16546 264192 16574
rect 260748 14816 260800 14822
rect 260748 14758 260800 14764
rect 260656 11688 260708 11694
rect 260656 11630 260708 11636
rect 259472 6886 259592 6914
rect 259472 480 259500 6886
rect 260668 480 260696 11630
rect 261772 480 261800 16546
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 264164 480 264192 16546
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 264992 354 265020 24414
rect 265636 14890 265664 51046
rect 266544 16108 266596 16114
rect 266544 16050 266596 16056
rect 265624 14884 265676 14890
rect 265624 14826 265676 14832
rect 266556 480 266584 16050
rect 267016 14958 267044 59463
rect 268566 59392 268622 59401
rect 268566 59327 268622 59336
rect 268382 59256 268438 59265
rect 268382 59191 268438 59200
rect 267740 33992 267792 33998
rect 267740 33934 267792 33940
rect 267004 14952 267056 14958
rect 267004 14894 267056 14900
rect 267752 4214 267780 33934
rect 267832 22976 267884 22982
rect 267832 22918 267884 22924
rect 267740 4208 267792 4214
rect 267740 4150 267792 4156
rect 267844 3482 267872 22918
rect 268396 15026 268424 59191
rect 268580 27062 268608 59327
rect 269120 31136 269172 31142
rect 269120 31078 269172 31084
rect 268568 27056 268620 27062
rect 268568 26998 268620 27004
rect 269132 16574 269160 31078
rect 269776 24274 269804 59463
rect 269960 29714 269988 59706
rect 270682 59664 270738 59673
rect 270682 59599 270738 59608
rect 270696 51074 270724 59599
rect 271892 58818 271920 59706
rect 272524 59696 272576 59702
rect 272524 59638 272576 59644
rect 276386 59664 276442 59673
rect 272246 59528 272302 59537
rect 272246 59463 272248 59472
rect 272300 59463 272302 59472
rect 272248 59434 272300 59440
rect 271880 58812 271932 58818
rect 271880 58754 271932 58760
rect 270696 51046 271184 51074
rect 270500 43716 270552 43722
rect 270500 43658 270552 43664
rect 269948 29708 270000 29714
rect 269948 29650 270000 29656
rect 269764 24268 269816 24274
rect 269764 24210 269816 24216
rect 270512 16574 270540 43658
rect 271156 25702 271184 51046
rect 271880 45212 271932 45218
rect 271880 45154 271932 45160
rect 271144 25696 271196 25702
rect 271144 25638 271196 25644
rect 271892 16574 271920 45154
rect 272536 42158 272564 59638
rect 276386 59599 276442 59608
rect 273902 59528 273958 59537
rect 273260 59492 273312 59498
rect 273902 59463 273904 59472
rect 273260 59434 273312 59440
rect 273956 59463 273958 59472
rect 273904 59434 273956 59440
rect 273272 57390 273300 59434
rect 276400 59401 276428 59599
rect 277228 59537 277256 59706
rect 277214 59528 277270 59537
rect 276664 59492 276716 59498
rect 277214 59463 277270 59472
rect 276664 59434 276716 59440
rect 276386 59392 276442 59401
rect 276386 59327 276442 59336
rect 273718 59256 273774 59265
rect 273718 59191 273774 59200
rect 274638 59256 274694 59265
rect 274638 59191 274694 59200
rect 273260 57384 273312 57390
rect 273260 57326 273312 57332
rect 273732 55214 273760 59191
rect 274652 56030 274680 59191
rect 274640 56024 274692 56030
rect 274640 55966 274692 55972
rect 273732 55186 273944 55214
rect 273260 45076 273312 45082
rect 273260 45018 273312 45024
rect 272524 42152 272576 42158
rect 272524 42094 272576 42100
rect 269132 16546 270080 16574
rect 270512 16546 270816 16574
rect 271892 16546 272472 16574
rect 268384 15020 268436 15026
rect 268384 14962 268436 14968
rect 268476 4208 268528 4214
rect 268476 4150 268528 4156
rect 267752 3454 267872 3482
rect 267752 480 267780 3454
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268488 354 268516 4150
rect 270052 480 270080 16546
rect 268814 354 268926 480
rect 268488 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 270788 354 270816 16546
rect 272444 480 272472 16546
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273272 354 273300 45018
rect 273916 28422 273944 55186
rect 276020 46504 276072 46510
rect 276020 46446 276072 46452
rect 274640 29912 274692 29918
rect 274640 29854 274692 29860
rect 273904 28416 273956 28422
rect 273904 28358 273956 28364
rect 274652 16574 274680 29854
rect 274652 16546 274864 16574
rect 274836 480 274864 16546
rect 276032 480 276060 46446
rect 276676 38078 276704 59434
rect 276846 59256 276902 59265
rect 276846 59191 276902 59200
rect 276860 39438 276888 59191
rect 277872 55214 277900 59706
rect 278056 59537 278084 59735
rect 278884 59537 278912 59735
rect 279422 59664 279478 59673
rect 279422 59599 279478 59608
rect 280342 59664 280398 59673
rect 280342 59599 280344 59608
rect 278042 59528 278098 59537
rect 278042 59463 278098 59472
rect 278870 59528 278926 59537
rect 278870 59463 278926 59472
rect 277950 59392 278006 59401
rect 278006 59350 278176 59378
rect 277950 59327 278006 59336
rect 277872 55186 278084 55214
rect 276848 39432 276900 39438
rect 276848 39374 276900 39380
rect 276664 38072 276716 38078
rect 276664 38014 276716 38020
rect 277400 35420 277452 35426
rect 277400 35362 277452 35368
rect 277412 16574 277440 35362
rect 278056 31142 278084 55186
rect 278148 50454 278176 59350
rect 278136 50448 278188 50454
rect 278136 50390 278188 50396
rect 279436 47666 279464 59599
rect 280396 59599 280398 59608
rect 280344 59570 280396 59576
rect 281736 59537 281764 59758
rect 286322 59800 286378 59809
rect 283010 59735 283012 59744
rect 283064 59735 283066 59744
rect 284300 59764 284352 59770
rect 283012 59706 283064 59712
rect 286322 59735 286378 59744
rect 287150 59800 287206 59809
rect 287150 59735 287206 59744
rect 287886 59800 287942 59809
rect 291750 59800 291806 59809
rect 287886 59735 287888 59744
rect 284300 59706 284352 59712
rect 282184 59628 282236 59634
rect 282184 59570 282236 59576
rect 280802 59528 280858 59537
rect 280802 59463 280858 59472
rect 281722 59528 281778 59537
rect 281722 59463 281778 59472
rect 279424 47660 279476 47666
rect 279424 47602 279476 47608
rect 278780 39704 278832 39710
rect 278780 39646 278832 39652
rect 278044 31136 278096 31142
rect 278044 31078 278096 31084
rect 278792 16574 278820 39646
rect 280816 17814 280844 59463
rect 280986 59392 281042 59401
rect 280986 59327 281042 59336
rect 281000 36718 281028 59327
rect 280988 36712 281040 36718
rect 280988 36654 281040 36660
rect 282196 20058 282224 59570
rect 283010 59528 283066 59537
rect 283010 59463 283066 59472
rect 282366 59256 282422 59265
rect 282366 59191 282422 59200
rect 282380 40866 282408 59191
rect 283024 51074 283052 59463
rect 284312 54738 284340 59706
rect 286336 59702 286364 59735
rect 286324 59696 286376 59702
rect 286324 59638 286376 59644
rect 286322 59528 286378 59537
rect 286322 59463 286378 59472
rect 284942 59256 284998 59265
rect 284942 59191 284998 59200
rect 284300 54732 284352 54738
rect 284300 54674 284352 54680
rect 283024 51046 283604 51074
rect 282368 40860 282420 40866
rect 282368 40802 282420 40808
rect 283576 39506 283604 51046
rect 284300 39636 284352 39642
rect 284300 39578 284352 39584
rect 283564 39500 283616 39506
rect 283564 39442 283616 39448
rect 282920 38276 282972 38282
rect 282920 38218 282972 38224
rect 282184 20052 282236 20058
rect 282184 19994 282236 20000
rect 280804 17808 280856 17814
rect 280804 17750 280856 17756
rect 282932 16574 282960 38218
rect 277412 16546 278360 16574
rect 278792 16546 279096 16574
rect 282932 16546 283144 16574
rect 276664 10736 276716 10742
rect 276664 10678 276716 10684
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276676 354 276704 10678
rect 278332 480 278360 16546
rect 277094 354 277206 480
rect 276676 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280712 10668 280764 10674
rect 280712 10610 280764 10616
rect 280724 480 280752 10610
rect 281908 8968 281960 8974
rect 281908 8910 281960 8916
rect 281920 480 281948 8910
rect 283116 480 283144 16546
rect 284312 480 284340 39578
rect 284956 29850 284984 59191
rect 286336 31278 286364 59463
rect 287164 59401 287192 59735
rect 287940 59735 287942 59744
rect 290648 59764 290700 59770
rect 287888 59706 287940 59712
rect 291750 59735 291806 59744
rect 293406 59800 293462 59809
rect 293406 59735 293462 59744
rect 293682 59800 293738 59809
rect 293682 59735 293684 59744
rect 290648 59706 290700 59712
rect 288440 59696 288492 59702
rect 287702 59664 287758 59673
rect 288440 59638 288492 59644
rect 289542 59664 289598 59673
rect 287702 59599 287758 59608
rect 287150 59392 287206 59401
rect 287150 59327 287206 59336
rect 286506 59256 286562 59265
rect 286506 59191 286562 59200
rect 286520 50590 286548 59191
rect 286508 50584 286560 50590
rect 286508 50526 286560 50532
rect 286324 31272 286376 31278
rect 286324 31214 286376 31220
rect 284944 29844 284996 29850
rect 284944 29786 284996 29792
rect 287716 21690 287744 59599
rect 288452 53310 288480 59638
rect 289542 59599 289598 59608
rect 289556 59401 289584 59599
rect 290462 59528 290518 59537
rect 290462 59463 290518 59472
rect 289082 59392 289138 59401
rect 289082 59327 289138 59336
rect 289542 59392 289598 59401
rect 289542 59327 289598 59336
rect 288440 53304 288492 53310
rect 288440 53246 288492 53252
rect 287704 21684 287756 21690
rect 287704 21626 287756 21632
rect 289096 15910 289124 59327
rect 290476 45082 290504 59463
rect 290660 49298 290688 59706
rect 291764 58546 291792 59735
rect 292026 59664 292082 59673
rect 292026 59599 292082 59608
rect 291842 59392 291898 59401
rect 291842 59327 291898 59336
rect 291752 58540 291804 58546
rect 291752 58482 291804 58488
rect 290648 49292 290700 49298
rect 290648 49234 290700 49240
rect 290464 45076 290516 45082
rect 290464 45018 290516 45024
rect 291856 15978 291884 59327
rect 292040 16046 292068 59599
rect 293420 58546 293448 59735
rect 293736 59735 293738 59744
rect 294418 59800 294474 59809
rect 296994 59800 296996 59809
rect 298928 59832 298980 59838
rect 297048 59800 297050 59809
rect 294418 59735 294474 59744
rect 295984 59764 296036 59770
rect 293684 59706 293736 59712
rect 294432 59401 294460 59735
rect 295984 59706 296036 59712
rect 296536 59764 296588 59770
rect 380072 59832 380124 59838
rect 298928 59774 298980 59780
rect 300306 59800 300362 59809
rect 296994 59735 297050 59744
rect 298744 59764 298796 59770
rect 296536 59706 296588 59712
rect 298744 59706 298796 59712
rect 294418 59392 294474 59401
rect 294418 59327 294474 59336
rect 294510 58984 294566 58993
rect 294510 58919 294566 58928
rect 293224 58540 293276 58546
rect 293224 58482 293276 58488
rect 293408 58540 293460 58546
rect 293408 58482 293460 58488
rect 293236 16114 293264 58482
rect 294524 55214 294552 58919
rect 294788 58540 294840 58546
rect 294788 58482 294840 58488
rect 294524 55186 294644 55214
rect 294616 16182 294644 55186
rect 294800 16250 294828 58482
rect 295996 16318 296024 59706
rect 296548 59673 296576 59706
rect 296534 59664 296590 59673
rect 296534 59599 296590 59608
rect 296994 59528 297050 59537
rect 296994 59463 297050 59472
rect 296166 59392 296222 59401
rect 296166 59327 296222 59336
rect 296180 36922 296208 59327
rect 297008 46442 297036 59463
rect 296996 46436 297048 46442
rect 296996 46378 297048 46384
rect 296168 36916 296220 36922
rect 296168 36858 296220 36864
rect 298756 34066 298784 59706
rect 298940 52086 298968 59774
rect 300306 59735 300362 59744
rect 301134 59800 301190 59809
rect 301134 59735 301190 59744
rect 301962 59800 302018 59809
rect 305918 59800 305974 59809
rect 301962 59735 301964 59744
rect 300320 59702 300348 59735
rect 300308 59696 300360 59702
rect 300308 59638 300360 59644
rect 300122 59528 300178 59537
rect 300122 59463 300178 59472
rect 298928 52080 298980 52086
rect 298928 52022 298980 52028
rect 299480 42356 299532 42362
rect 299480 42298 299532 42304
rect 298744 34060 298796 34066
rect 298744 34002 298796 34008
rect 296720 20324 296772 20330
rect 296720 20266 296772 20272
rect 296732 16574 296760 20266
rect 296732 16546 297312 16574
rect 295984 16312 296036 16318
rect 295984 16254 296036 16260
rect 294788 16244 294840 16250
rect 294788 16186 294840 16192
rect 294604 16176 294656 16182
rect 294604 16118 294656 16124
rect 293224 16108 293276 16114
rect 293224 16050 293276 16056
rect 292028 16040 292080 16046
rect 292028 15982 292080 15988
rect 291844 15972 291896 15978
rect 291844 15914 291896 15920
rect 289084 15904 289136 15910
rect 289084 15846 289136 15852
rect 286600 10668 286652 10674
rect 286600 10610 286652 10616
rect 285404 9036 285456 9042
rect 285404 8978 285456 8984
rect 285416 480 285444 8978
rect 286612 480 286640 10610
rect 287336 10600 287388 10606
rect 287336 10542 287388 10548
rect 289820 10600 289872 10606
rect 289820 10542 289872 10548
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 354 287376 10542
rect 288992 9104 289044 9110
rect 288992 9046 289044 9052
rect 289004 480 289032 9046
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 289832 354 289860 10542
rect 291384 10532 291436 10538
rect 291384 10474 291436 10480
rect 293224 10532 293276 10538
rect 293224 10474 293276 10480
rect 291396 480 291424 10474
rect 292580 9172 292632 9178
rect 292580 9114 292632 9120
rect 292592 480 292620 9114
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 10474
rect 294880 10464 294932 10470
rect 294880 10406 294932 10412
rect 294892 480 294920 10406
rect 296076 9240 296128 9246
rect 296076 9182 296128 9188
rect 296088 480 296116 9182
rect 297284 480 297312 16546
rect 298100 10396 298152 10402
rect 298100 10338 298152 10344
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 354 298140 10338
rect 299492 3482 299520 42298
rect 299572 21752 299624 21758
rect 299572 21694 299624 21700
rect 299584 4214 299612 21694
rect 300136 13258 300164 59463
rect 301148 59401 301176 59735
rect 302016 59735 302018 59744
rect 304264 59764 304316 59770
rect 301964 59706 302016 59712
rect 305918 59735 305974 59744
rect 312634 59800 312690 59809
rect 312634 59735 312690 59744
rect 314290 59800 314346 59809
rect 316774 59800 316830 59809
rect 314290 59735 314292 59744
rect 304264 59706 304316 59712
rect 302884 59696 302936 59702
rect 301502 59664 301558 59673
rect 302884 59638 302936 59644
rect 301502 59599 301558 59608
rect 300306 59392 300362 59401
rect 300306 59327 300362 59336
rect 301134 59392 301190 59401
rect 301134 59327 301190 59336
rect 300320 32774 300348 59327
rect 300308 32768 300360 32774
rect 300308 32710 300360 32716
rect 301516 13326 301544 59599
rect 302240 38208 302292 38214
rect 302240 38150 302292 38156
rect 301504 13320 301556 13326
rect 301504 13262 301556 13268
rect 300124 13252 300176 13258
rect 300124 13194 300176 13200
rect 301504 10328 301556 10334
rect 301504 10270 301556 10276
rect 299572 4208 299624 4214
rect 299572 4150 299624 4156
rect 300768 4208 300820 4214
rect 300768 4150 300820 4156
rect 299492 3454 299704 3482
rect 299676 480 299704 3454
rect 300780 480 300808 4150
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 10270
rect 302252 6914 302280 38150
rect 302896 13394 302924 59638
rect 303066 59256 303122 59265
rect 303066 59191 303122 59200
rect 303080 41002 303108 59191
rect 303068 40996 303120 41002
rect 303068 40938 303120 40944
rect 304276 13462 304304 59706
rect 304354 59664 304410 59673
rect 304354 59599 304410 59608
rect 304368 59401 304396 59599
rect 305642 59528 305698 59537
rect 305642 59463 305698 59472
rect 304354 59392 304410 59401
rect 304354 59327 304410 59336
rect 304446 59256 304502 59265
rect 304446 59191 304502 59200
rect 304460 13530 304488 59191
rect 305656 13598 305684 59463
rect 305932 59129 305960 59735
rect 312544 59696 312596 59702
rect 306010 59664 306066 59673
rect 310150 59664 310206 59673
rect 306010 59599 306012 59608
rect 306064 59599 306066 59608
rect 307208 59628 307260 59634
rect 306012 59570 306064 59576
rect 310150 59599 310152 59608
rect 307208 59570 307260 59576
rect 310204 59599 310206 59608
rect 312542 59664 312544 59673
rect 312596 59664 312598 59673
rect 312542 59599 312598 59608
rect 310152 59570 310204 59576
rect 306838 59392 306894 59401
rect 306838 59327 306840 59336
rect 306892 59327 306894 59336
rect 306840 59298 306892 59304
rect 307022 59256 307078 59265
rect 307022 59191 307078 59200
rect 305918 59120 305974 59129
rect 305918 59055 305974 59064
rect 307036 13666 307064 59191
rect 307220 45150 307248 59570
rect 308494 59528 308550 59537
rect 312542 59528 312598 59537
rect 308494 59463 308496 59472
rect 308548 59463 308550 59472
rect 311164 59492 311216 59498
rect 308496 59434 308548 59440
rect 312542 59463 312598 59472
rect 311164 59434 311216 59440
rect 308404 59356 308456 59362
rect 308404 59298 308456 59304
rect 310520 59356 310572 59362
rect 310520 59298 310572 59304
rect 308416 46578 308444 59298
rect 309782 59256 309838 59265
rect 309782 59191 309838 59200
rect 308586 59120 308642 59129
rect 308586 59055 308642 59064
rect 308600 53446 308628 59055
rect 308588 53440 308640 53446
rect 308588 53382 308640 53388
rect 308404 46572 308456 46578
rect 308404 46514 308456 46520
rect 307208 45144 307260 45150
rect 307208 45086 307260 45092
rect 307760 42424 307812 42430
rect 307760 42366 307812 42372
rect 307024 13660 307076 13666
rect 307024 13602 307076 13608
rect 305644 13592 305696 13598
rect 305644 13534 305696 13540
rect 304448 13524 304500 13530
rect 304448 13466 304500 13472
rect 304264 13456 304316 13462
rect 304264 13398 304316 13404
rect 302884 13388 302936 13394
rect 302884 13330 302936 13336
rect 305552 12028 305604 12034
rect 305552 11970 305604 11976
rect 303896 10328 303948 10334
rect 303896 10270 303948 10276
rect 302252 6886 303200 6914
rect 303172 480 303200 6886
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 10270
rect 305564 480 305592 11970
rect 306748 9308 306800 9314
rect 306748 9250 306800 9256
rect 306760 480 306788 9250
rect 307772 3330 307800 42366
rect 309796 11966 309824 59191
rect 309784 11960 309836 11966
rect 309784 11902 309836 11908
rect 307944 10396 307996 10402
rect 307944 10338 307996 10344
rect 307760 3324 307812 3330
rect 307760 3266 307812 3272
rect 307956 480 307984 10338
rect 310244 9376 310296 9382
rect 310244 9318 310296 9324
rect 309048 3324 309100 3330
rect 309048 3266 309100 3272
rect 309060 480 309088 3266
rect 310256 480 310284 9318
rect 310532 6914 310560 59298
rect 311176 12034 311204 59434
rect 311346 59392 311402 59401
rect 311346 59327 311402 59336
rect 311360 12102 311388 59327
rect 312556 12238 312584 59463
rect 312648 59401 312676 59735
rect 314344 59735 314346 59744
rect 316684 59764 316736 59770
rect 314292 59706 314344 59712
rect 316774 59735 316830 59744
rect 316958 59800 317014 59809
rect 316958 59735 317014 59744
rect 320822 59800 320878 59809
rect 324134 59800 324190 59809
rect 320822 59735 320824 59744
rect 316684 59706 316736 59712
rect 313924 59696 313976 59702
rect 313924 59638 313976 59644
rect 312728 59628 312780 59634
rect 312728 59570 312780 59576
rect 312634 59392 312690 59401
rect 312634 59327 312690 59336
rect 312544 12232 312596 12238
rect 312544 12174 312596 12180
rect 312740 12170 312768 59570
rect 313280 39636 313332 39642
rect 313280 39578 313332 39584
rect 313292 16574 313320 39578
rect 313292 16546 313872 16574
rect 312728 12164 312780 12170
rect 312728 12106 312780 12112
rect 311348 12096 311400 12102
rect 311348 12038 311400 12044
rect 311164 12028 311216 12034
rect 311164 11970 311216 11976
rect 312176 11892 312228 11898
rect 312176 11834 312228 11840
rect 310532 6886 311480 6914
rect 311452 480 311480 6886
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 354 312216 11834
rect 313844 480 313872 16546
rect 313936 11898 313964 59638
rect 314290 59528 314346 59537
rect 314346 59486 314700 59514
rect 314290 59463 314346 59472
rect 314672 57594 314700 59486
rect 315302 59256 315358 59265
rect 315302 59191 315358 59200
rect 314660 57588 314712 57594
rect 314660 57530 314712 57536
rect 315316 34134 315344 59191
rect 316040 49360 316092 49366
rect 316040 49302 316092 49308
rect 315304 34128 315356 34134
rect 315304 34070 315356 34076
rect 313924 11892 313976 11898
rect 313924 11834 313976 11840
rect 314660 10464 314712 10470
rect 314660 10406 314712 10412
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314672 354 314700 10406
rect 316052 3482 316080 49302
rect 316132 24404 316184 24410
rect 316132 24346 316184 24352
rect 316144 4214 316172 24346
rect 316696 22166 316724 59706
rect 316788 59401 316816 59735
rect 316774 59392 316830 59401
rect 316972 59362 317000 59735
rect 320876 59735 320878 59744
rect 323124 59764 323176 59770
rect 320824 59706 320876 59712
rect 324134 59735 324190 59744
rect 324962 59800 325018 59809
rect 330298 59800 330354 59809
rect 324962 59735 324964 59744
rect 323124 59706 323176 59712
rect 317418 59664 317474 59673
rect 317418 59599 317474 59608
rect 322478 59664 322534 59673
rect 322478 59599 322534 59608
rect 316774 59327 316830 59336
rect 316960 59356 317012 59362
rect 316960 59298 317012 59304
rect 316866 59256 316922 59265
rect 316866 59191 316922 59200
rect 316880 26042 316908 59191
rect 316868 26036 316920 26042
rect 316868 25978 316920 25984
rect 316684 22160 316736 22166
rect 316684 22102 316736 22108
rect 317432 16574 317460 59599
rect 320362 59528 320418 59537
rect 320362 59463 320418 59472
rect 318890 59256 318946 59265
rect 318890 59191 318946 59200
rect 318800 29980 318852 29986
rect 318800 29922 318852 29928
rect 317432 16546 318104 16574
rect 316132 4208 316184 4214
rect 316132 4150 316184 4156
rect 317328 4208 317380 4214
rect 317328 4150 317380 4156
rect 316052 3454 316264 3482
rect 316236 480 316264 3454
rect 317340 480 317368 4150
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 318812 6914 318840 29922
rect 318904 10470 318932 59191
rect 320180 58880 320232 58886
rect 320180 58822 320232 58828
rect 318892 10464 318944 10470
rect 318892 10406 318944 10412
rect 320192 6914 320220 58822
rect 320376 10334 320404 59463
rect 322492 59401 322520 59599
rect 320546 59392 320602 59401
rect 320546 59327 320602 59336
rect 321650 59392 321706 59401
rect 321650 59327 321706 59336
rect 322478 59392 322534 59401
rect 322478 59327 322534 59336
rect 320560 10402 320588 59327
rect 321560 26036 321612 26042
rect 321560 25978 321612 25984
rect 321572 16574 321600 25978
rect 321664 21758 321692 59327
rect 322940 36848 322992 36854
rect 322940 36790 322992 36796
rect 321652 21752 321704 21758
rect 321652 21694 321704 21700
rect 321572 16546 322152 16574
rect 320548 10396 320600 10402
rect 320548 10338 320600 10344
rect 320364 10328 320416 10334
rect 320364 10270 320416 10276
rect 318812 6886 319760 6914
rect 320192 6886 320496 6914
rect 319732 480 319760 6886
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 6886
rect 322124 480 322152 16546
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 322952 354 322980 36790
rect 323136 20330 323164 59706
rect 323306 59528 323362 59537
rect 323306 59463 323362 59472
rect 323124 20324 323176 20330
rect 323124 20266 323176 20272
rect 323320 10538 323348 59463
rect 324148 59401 324176 59735
rect 325016 59735 325018 59744
rect 327356 59764 327408 59770
rect 324964 59706 325016 59712
rect 330298 59735 330354 59744
rect 334898 59800 334954 59809
rect 339038 59800 339094 59809
rect 334898 59735 334900 59744
rect 327356 59706 327408 59712
rect 324778 59664 324834 59673
rect 324778 59599 324834 59608
rect 324134 59392 324190 59401
rect 324134 59327 324190 59336
rect 324594 59256 324650 59265
rect 324594 59191 324650 59200
rect 324320 25832 324372 25838
rect 324320 25774 324372 25780
rect 323308 10532 323360 10538
rect 323308 10474 323360 10480
rect 324332 3210 324360 25774
rect 324412 22160 324464 22166
rect 324412 22102 324464 22108
rect 324424 3330 324452 22102
rect 324608 10606 324636 59191
rect 324792 10674 324820 59599
rect 325790 59392 325846 59401
rect 325790 59327 325792 59336
rect 325844 59327 325846 59336
rect 327172 59356 327224 59362
rect 325792 59298 325844 59304
rect 327172 59298 327224 59304
rect 325698 59256 325754 59265
rect 325698 59191 325754 59200
rect 325712 38282 325740 59191
rect 327184 46510 327212 59298
rect 327172 46504 327224 46510
rect 327172 46446 327224 46452
rect 327368 39710 327396 59706
rect 329102 59528 329158 59537
rect 329102 59463 329104 59472
rect 329156 59463 329158 59472
rect 329104 59434 329156 59440
rect 329930 59392 329986 59401
rect 329930 59327 329986 59336
rect 328826 59256 328882 59265
rect 328826 59191 328882 59200
rect 328642 59120 328698 59129
rect 328642 59055 328698 59064
rect 328460 57588 328512 57594
rect 328460 57530 328512 57536
rect 327356 39704 327408 39710
rect 327356 39646 327408 39652
rect 325700 38276 325752 38282
rect 325700 38218 325752 38224
rect 325700 35488 325752 35494
rect 325700 35430 325752 35436
rect 325712 16574 325740 35430
rect 327080 27260 327132 27266
rect 327080 27202 327132 27208
rect 327092 16574 327120 27202
rect 328472 16574 328500 57530
rect 328656 45218 328684 59055
rect 328644 45212 328696 45218
rect 328644 45154 328696 45160
rect 328840 33998 328868 59191
rect 329840 54800 329892 54806
rect 329840 54742 329892 54748
rect 328828 33992 328880 33998
rect 328828 33934 328880 33940
rect 329852 16574 329880 54742
rect 329944 24478 329972 59327
rect 330312 58954 330340 59735
rect 334952 59735 334954 59744
rect 336924 59764 336976 59770
rect 334900 59706 334952 59712
rect 341522 59800 341578 59809
rect 339038 59735 339040 59744
rect 336924 59706 336976 59712
rect 339092 59735 339094 59744
rect 341156 59764 341208 59770
rect 339040 59706 339092 59712
rect 343086 59800 343142 59809
rect 341522 59735 341524 59744
rect 341156 59706 341208 59712
rect 341576 59735 341578 59744
rect 342536 59764 342588 59770
rect 341524 59706 341576 59712
rect 347962 59800 348018 59809
rect 343086 59735 343088 59744
rect 342536 59706 342588 59712
rect 343140 59735 343142 59744
rect 345112 59764 345164 59770
rect 343088 59706 343140 59712
rect 347962 59735 348018 59744
rect 348422 59800 348478 59809
rect 348422 59735 348478 59744
rect 355230 59800 355286 59809
rect 355230 59735 355286 59744
rect 359554 59800 359610 59809
rect 363694 59800 363750 59809
rect 359554 59735 359556 59744
rect 345112 59706 345164 59712
rect 333242 59664 333298 59673
rect 333242 59599 333298 59608
rect 331494 59528 331550 59537
rect 331312 59492 331364 59498
rect 331494 59463 331550 59472
rect 331312 59434 331364 59440
rect 330300 58948 330352 58954
rect 330300 58890 330352 58896
rect 331220 57588 331272 57594
rect 331220 57530 331272 57536
rect 329932 24472 329984 24478
rect 329932 24414 329984 24420
rect 325712 16546 326384 16574
rect 327092 16546 328040 16574
rect 328472 16546 328776 16574
rect 329852 16546 330432 16574
rect 324780 10668 324832 10674
rect 324780 10610 324832 10616
rect 324596 10600 324648 10606
rect 324596 10542 324648 10548
rect 324412 3324 324464 3330
rect 324412 3266 324464 3272
rect 325608 3324 325660 3330
rect 325608 3266 325660 3272
rect 324332 3182 324452 3210
rect 324424 480 324452 3182
rect 325620 480 325648 3266
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 16546
rect 328012 480 328040 16546
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 328748 354 328776 16546
rect 330404 480 330432 16546
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331232 354 331260 57530
rect 331324 32706 331352 59434
rect 331508 53378 331536 59463
rect 333256 59401 333284 59599
rect 334070 59528 334126 59537
rect 334070 59463 334126 59472
rect 332690 59392 332746 59401
rect 332690 59327 332746 59336
rect 333242 59392 333298 59401
rect 333242 59327 333298 59336
rect 331496 53372 331548 53378
rect 331496 53314 331548 53320
rect 332600 50652 332652 50658
rect 332600 50594 332652 50600
rect 331312 32700 331364 32706
rect 331312 32642 331364 32648
rect 332612 3330 332640 50594
rect 332704 41070 332732 59327
rect 332692 41064 332744 41070
rect 332692 41006 332744 41012
rect 332692 34128 332744 34134
rect 332692 34070 332744 34076
rect 332600 3324 332652 3330
rect 332600 3266 332652 3272
rect 332704 480 332732 34070
rect 333980 28552 334032 28558
rect 333980 28494 334032 28500
rect 333888 3324 333940 3330
rect 333888 3266 333940 3272
rect 333900 480 333928 3266
rect 333992 626 334020 28494
rect 334084 6594 334112 59463
rect 335358 59392 335414 59401
rect 335358 59327 335414 59336
rect 335372 57526 335400 59327
rect 335542 59256 335598 59265
rect 335542 59191 335598 59200
rect 335450 59120 335506 59129
rect 335450 59055 335506 59064
rect 335360 57520 335412 57526
rect 335360 57462 335412 57468
rect 335464 45554 335492 59055
rect 335372 45526 335492 45554
rect 335372 25906 335400 45526
rect 335360 25900 335412 25906
rect 335360 25842 335412 25848
rect 335452 11892 335504 11898
rect 335452 11834 335504 11840
rect 334072 6588 334124 6594
rect 334072 6530 334124 6536
rect 335464 3482 335492 11834
rect 335556 6526 335584 59191
rect 336936 52018 336964 59706
rect 338118 59528 338174 59537
rect 338118 59463 338174 59472
rect 340970 59528 341026 59537
rect 340970 59463 341026 59472
rect 336924 52012 336976 52018
rect 336924 51954 336976 51960
rect 336740 47932 336792 47938
rect 336740 47874 336792 47880
rect 336752 16574 336780 47874
rect 336752 16546 337056 16574
rect 335544 6520 335596 6526
rect 335544 6462 335596 6468
rect 335464 3454 336320 3482
rect 333992 598 334664 626
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 598
rect 336292 480 336320 3454
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 338132 6390 338160 59463
rect 338210 59392 338266 59401
rect 338210 59327 338266 59336
rect 339590 59392 339646 59401
rect 339590 59327 339646 59336
rect 338224 6458 338252 59327
rect 339500 12232 339552 12238
rect 339500 12174 339552 12180
rect 338672 11892 338724 11898
rect 338672 11834 338724 11840
rect 338212 6452 338264 6458
rect 338212 6394 338264 6400
rect 338120 6384 338172 6390
rect 338120 6326 338172 6332
rect 338684 480 338712 11834
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339512 354 339540 12174
rect 339604 6322 339632 59327
rect 340880 31340 340932 31346
rect 340880 31282 340932 31288
rect 339592 6316 339644 6322
rect 339592 6258 339644 6264
rect 340144 5364 340196 5370
rect 340144 5306 340196 5312
rect 340156 4962 340184 5306
rect 340144 4956 340196 4962
rect 340144 4898 340196 4904
rect 340892 3210 340920 31282
rect 340984 27198 341012 59463
rect 340972 27192 341024 27198
rect 340972 27134 341024 27140
rect 340972 20324 341024 20330
rect 340972 20266 341024 20272
rect 340984 3330 341012 20266
rect 341168 6254 341196 59706
rect 342350 59392 342406 59401
rect 342350 59327 342406 59336
rect 342260 12164 342312 12170
rect 342260 12106 342312 12112
rect 341156 6248 341208 6254
rect 341156 6190 341208 6196
rect 340972 3324 341024 3330
rect 340972 3266 341024 3272
rect 342168 3324 342220 3330
rect 342168 3266 342220 3272
rect 340892 3182 341012 3210
rect 340984 480 341012 3182
rect 342180 480 342208 3266
rect 342272 626 342300 12106
rect 342364 5302 342392 59327
rect 342352 5296 342404 5302
rect 342352 5238 342404 5244
rect 342548 5234 342576 59706
rect 343638 59528 343694 59537
rect 343638 59463 343694 59472
rect 344742 59528 344798 59537
rect 344742 59463 344744 59472
rect 343652 50522 343680 59463
rect 344796 59463 344798 59472
rect 344744 59434 344796 59440
rect 343640 50516 343692 50522
rect 343640 50458 343692 50464
rect 343640 43784 343692 43790
rect 343640 43726 343692 43732
rect 343652 16574 343680 43726
rect 343652 16546 344600 16574
rect 342536 5228 342588 5234
rect 342536 5170 342588 5176
rect 342272 598 342944 626
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 598
rect 344572 480 344600 16546
rect 345020 10328 345072 10334
rect 345020 10270 345072 10276
rect 345032 490 345060 10270
rect 345124 5166 345152 59706
rect 347976 59537 348004 59735
rect 348054 59664 348110 59673
rect 348054 59599 348110 59608
rect 347962 59528 348018 59537
rect 346492 59492 346544 59498
rect 347962 59463 348018 59472
rect 346492 59434 346544 59440
rect 345294 59392 345350 59401
rect 345294 59327 345350 59336
rect 345308 16574 345336 59327
rect 346398 59256 346454 59265
rect 346398 59191 346454 59200
rect 345308 16546 345428 16574
rect 345112 5160 345164 5166
rect 345112 5102 345164 5108
rect 345400 5098 345428 16546
rect 346412 5370 346440 59191
rect 346400 5364 346452 5370
rect 346400 5306 346452 5312
rect 345388 5092 345440 5098
rect 345388 5034 345440 5040
rect 346504 5030 346532 59434
rect 348068 59401 348096 59599
rect 347870 59392 347926 59401
rect 347870 59327 347926 59336
rect 348054 59392 348110 59401
rect 348054 59327 348110 59336
rect 347780 20256 347832 20262
rect 347780 20198 347832 20204
rect 346952 12096 347004 12102
rect 346952 12038 347004 12044
rect 346492 5024 346544 5030
rect 346492 4966 346544 4972
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345032 462 345336 490
rect 346964 480 346992 12038
rect 347792 3482 347820 20198
rect 347884 4894 347912 59327
rect 348436 56166 348464 59735
rect 354600 59622 355088 59650
rect 349250 59528 349306 59537
rect 349250 59463 349306 59472
rect 351366 59528 351422 59537
rect 351366 59463 351368 59472
rect 349160 56228 349212 56234
rect 349160 56170 349212 56176
rect 348424 56160 348476 56166
rect 348424 56102 348476 56108
rect 347872 4888 347924 4894
rect 347872 4830 347924 4836
rect 347792 3454 348096 3482
rect 348068 480 348096 3454
rect 349172 3210 349200 56170
rect 349264 31210 349292 59463
rect 351420 59463 351422 59472
rect 353576 59492 353628 59498
rect 351368 59434 351420 59440
rect 353576 59434 353628 59440
rect 349434 59392 349490 59401
rect 349434 59327 349490 59336
rect 349252 31204 349304 31210
rect 349252 31146 349304 31152
rect 349252 12028 349304 12034
rect 349252 11970 349304 11976
rect 349264 3330 349292 11970
rect 349448 4826 349476 59327
rect 350538 59256 350594 59265
rect 350538 59191 350594 59200
rect 351918 59256 351974 59265
rect 351918 59191 351974 59200
rect 353390 59256 353446 59265
rect 353390 59191 353446 59200
rect 350552 36786 350580 59191
rect 351932 47870 351960 59191
rect 351920 47864 351972 47870
rect 351920 47806 351972 47812
rect 353404 46374 353432 59191
rect 353392 46368 353444 46374
rect 353392 46310 353444 46316
rect 353588 44946 353616 59434
rect 354600 59401 354628 59622
rect 354954 59528 355010 59537
rect 354876 59486 354954 59514
rect 354586 59392 354642 59401
rect 354586 59327 354642 59336
rect 354876 47734 354904 59486
rect 354954 59463 355010 59472
rect 354864 47728 354916 47734
rect 354864 47670 354916 47676
rect 355060 45554 355088 59622
rect 355244 59401 355272 59735
rect 359608 59735 359610 59744
rect 361764 59764 361816 59770
rect 359556 59706 359608 59712
rect 363694 59735 363696 59744
rect 361764 59706 361816 59712
rect 363748 59735 363750 59744
rect 365166 59800 365222 59809
rect 367006 59800 367062 59809
rect 365166 59735 365222 59744
rect 366364 59764 366416 59770
rect 363696 59706 363748 59712
rect 357070 59664 357126 59673
rect 357070 59599 357126 59608
rect 358910 59664 358966 59673
rect 358910 59599 358966 59608
rect 356058 59528 356114 59537
rect 356058 59463 356114 59472
rect 355230 59392 355286 59401
rect 355230 59327 355286 59336
rect 354968 45526 355088 45554
rect 353576 44940 353628 44946
rect 353576 44882 353628 44888
rect 354968 43654 354996 45526
rect 354956 43648 355008 43654
rect 354956 43590 355008 43596
rect 350632 38140 350684 38146
rect 350632 38082 350684 38088
rect 350540 36780 350592 36786
rect 350540 36722 350592 36728
rect 350644 16574 350672 38082
rect 354680 23044 354732 23050
rect 354680 22986 354732 22992
rect 354692 16574 354720 22986
rect 350644 16546 351224 16574
rect 354692 16546 355272 16574
rect 349436 4820 349488 4826
rect 349436 4762 349488 4768
rect 349252 3324 349304 3330
rect 349252 3266 349304 3272
rect 350448 3324 350500 3330
rect 350448 3266 350500 3272
rect 349172 3182 349292 3210
rect 349264 480 349292 3182
rect 350460 480 350488 3266
rect 345308 354 345336 462
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 353576 11960 353628 11966
rect 353576 11902 353628 11908
rect 352840 10396 352892 10402
rect 352840 10338 352892 10344
rect 352852 480 352880 10338
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 353588 354 353616 11902
rect 355244 480 355272 16546
rect 356072 13190 356100 59463
rect 357084 59401 357112 59599
rect 357622 59528 357678 59537
rect 357622 59463 357678 59472
rect 357070 59392 357126 59401
rect 357070 59327 357126 59336
rect 357440 46572 357492 46578
rect 357440 46514 357492 46520
rect 356060 13184 356112 13190
rect 356060 13126 356112 13132
rect 356336 10464 356388 10470
rect 356336 10406 356388 10412
rect 356348 480 356376 10406
rect 357452 3210 357480 46514
rect 357532 25764 357584 25770
rect 357532 25706 357584 25712
rect 357544 3330 357572 25706
rect 357636 11830 357664 59463
rect 358818 59392 358874 59401
rect 358818 59327 358874 59336
rect 357806 59256 357862 59265
rect 357806 59191 357862 59200
rect 357820 13122 357848 59191
rect 358832 42226 358860 59327
rect 358924 49162 358952 59599
rect 360198 59392 360254 59401
rect 360254 59350 360332 59378
rect 360198 59327 360254 59336
rect 360200 53440 360252 53446
rect 360200 53382 360252 53388
rect 358912 49156 358964 49162
rect 358912 49098 358964 49104
rect 358820 42220 358872 42226
rect 358820 42162 358872 42168
rect 357808 13116 357860 13122
rect 357808 13058 357860 13064
rect 357624 11824 357676 11830
rect 357624 11766 357676 11772
rect 359464 10532 359516 10538
rect 359464 10474 359516 10480
rect 357532 3324 357584 3330
rect 357532 3266 357584 3272
rect 358728 3324 358780 3330
rect 358728 3266 358780 3272
rect 357452 3182 357572 3210
rect 357544 480 357572 3182
rect 358740 480 358768 3266
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 10474
rect 360212 3482 360240 53382
rect 360304 6186 360332 59350
rect 361578 59256 361634 59265
rect 361578 59191 361634 59200
rect 361592 54602 361620 59191
rect 361580 54596 361632 54602
rect 361580 54538 361632 54544
rect 361580 45008 361632 45014
rect 361580 44950 361632 44956
rect 361592 16574 361620 44950
rect 361776 28490 361804 59706
rect 365180 59702 365208 59735
rect 369398 59800 369454 59809
rect 367006 59735 367008 59744
rect 366364 59706 366416 59712
rect 367060 59735 367062 59744
rect 369124 59764 369176 59770
rect 367008 59706 367060 59712
rect 369398 59735 369400 59744
rect 369124 59706 369176 59712
rect 369452 59735 369454 59744
rect 371054 59800 371110 59809
rect 376022 59800 376078 59809
rect 371054 59735 371056 59744
rect 369400 59706 369452 59712
rect 371108 59735 371110 59744
rect 372620 59764 372672 59770
rect 371056 59706 371108 59712
rect 380070 59800 380072 59809
rect 382924 59832 382976 59838
rect 380124 59800 380126 59809
rect 376022 59735 376024 59744
rect 372620 59706 372672 59712
rect 376076 59735 376078 59744
rect 378968 59764 379020 59770
rect 376024 59706 376076 59712
rect 378968 59706 379020 59712
rect 379428 59764 379480 59770
rect 380990 59800 381046 59809
rect 380070 59735 380126 59744
rect 380164 59764 380216 59770
rect 379428 59706 379480 59712
rect 382924 59774 382976 59780
rect 387522 59800 387578 59809
rect 380990 59735 380992 59744
rect 380164 59706 380216 59712
rect 381044 59735 381046 59744
rect 382280 59764 382332 59770
rect 380992 59706 381044 59712
rect 382280 59706 382332 59712
rect 365168 59696 365220 59702
rect 364982 59664 365038 59673
rect 365168 59638 365220 59644
rect 364982 59599 365038 59608
rect 363786 59528 363842 59537
rect 363786 59463 363842 59472
rect 363602 59392 363658 59401
rect 363602 59327 363658 59336
rect 361764 28484 361816 28490
rect 361764 28426 361816 28432
rect 361592 16546 361896 16574
rect 360292 6180 360344 6186
rect 360292 6122 360344 6128
rect 360212 3454 361160 3482
rect 361132 480 361160 3454
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 361868 354 361896 16546
rect 363512 10600 363564 10606
rect 363512 10542 363564 10548
rect 363524 480 363552 10542
rect 363616 6186 363644 59327
rect 363800 6254 363828 59463
rect 364340 45144 364392 45150
rect 364340 45086 364392 45092
rect 364352 16574 364380 45086
rect 364352 16546 364656 16574
rect 363788 6248 363840 6254
rect 363788 6190 363840 6196
rect 363604 6180 363656 6186
rect 363604 6122 363656 6128
rect 364628 480 364656 16546
rect 364996 6322 365024 59599
rect 365720 53236 365772 53242
rect 365720 53178 365772 53184
rect 364984 6316 365036 6322
rect 364984 6258 365036 6264
rect 365732 3210 365760 53178
rect 366376 44946 366404 59706
rect 366548 59696 366600 59702
rect 366548 59638 366600 59644
rect 366560 46374 366588 59638
rect 367742 59256 367798 59265
rect 367798 59214 367968 59242
rect 367742 59191 367798 59200
rect 367742 59120 367798 59129
rect 367742 59055 367798 59064
rect 366548 46368 366600 46374
rect 366548 46310 366600 46316
rect 366364 44940 366416 44946
rect 366364 44882 366416 44888
rect 367756 36786 367784 59055
rect 367940 47734 367968 59214
rect 369136 49162 369164 59706
rect 371332 59696 371384 59702
rect 371054 59664 371110 59673
rect 371110 59622 371280 59650
rect 371332 59638 371384 59644
rect 371054 59599 371110 59608
rect 369950 59528 370006 59537
rect 369950 59463 370006 59472
rect 370686 59528 370742 59537
rect 370686 59463 370742 59472
rect 369964 59401 369992 59463
rect 369950 59392 370006 59401
rect 369950 59327 370006 59336
rect 370502 59392 370558 59401
rect 370502 59327 370558 59336
rect 369124 49156 369176 49162
rect 369124 49098 369176 49104
rect 367928 47728 367980 47734
rect 367928 47670 367980 47676
rect 368480 39568 368532 39574
rect 368480 39510 368532 39516
rect 367744 36780 367796 36786
rect 367744 36722 367796 36728
rect 368492 16574 368520 39510
rect 370516 33998 370544 59327
rect 370700 50522 370728 59463
rect 371252 51074 371280 59622
rect 371344 52018 371372 59638
rect 372632 53242 372660 59706
rect 376022 59664 376078 59673
rect 378506 59664 378562 59673
rect 376022 59599 376024 59608
rect 376076 59599 376078 59608
rect 377404 59628 377456 59634
rect 376024 59570 376076 59576
rect 378506 59599 378562 59608
rect 377404 59570 377456 59576
rect 372710 59528 372766 59537
rect 376022 59528 376078 59537
rect 372710 59463 372712 59472
rect 372764 59463 372766 59472
rect 374000 59492 374052 59498
rect 372712 59434 372764 59440
rect 376022 59463 376078 59472
rect 374000 59434 374052 59440
rect 374012 54602 374040 59434
rect 374642 59256 374698 59265
rect 374642 59191 374698 59200
rect 374000 54596 374052 54602
rect 374000 54538 374052 54544
rect 372620 53236 372672 53242
rect 372620 53178 372672 53184
rect 371332 52012 371384 52018
rect 371332 51954 371384 51960
rect 371252 51046 371924 51074
rect 370688 50516 370740 50522
rect 370688 50458 370740 50464
rect 370504 33992 370556 33998
rect 370504 33934 370556 33940
rect 368492 16546 369440 16574
rect 367744 13660 367796 13666
rect 367744 13602 367796 13608
rect 365812 11960 365864 11966
rect 365812 11902 365864 11908
rect 365824 3330 365852 11902
rect 365812 3324 365864 3330
rect 365812 3266 365864 3272
rect 367008 3324 367060 3330
rect 367008 3266 367060 3272
rect 365732 3182 365852 3210
rect 365824 480 365852 3182
rect 367020 480 367048 3266
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 13602
rect 369412 480 369440 16546
rect 371240 13592 371292 13598
rect 371240 13534 371292 13540
rect 370136 10668 370188 10674
rect 370136 10610 370188 10616
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370148 354 370176 10610
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 371252 354 371280 13534
rect 371896 4826 371924 51046
rect 372620 42288 372672 42294
rect 372620 42230 372672 42236
rect 372632 16574 372660 42230
rect 374656 32706 374684 59191
rect 374644 32700 374696 32706
rect 374644 32642 374696 32648
rect 374000 31340 374052 31346
rect 374000 31282 374052 31288
rect 372632 16546 372936 16574
rect 371884 4820 371936 4826
rect 371884 4762 371936 4768
rect 372908 480 372936 16546
rect 374012 3210 374040 31282
rect 375380 20188 375432 20194
rect 375380 20130 375432 20136
rect 374092 13524 374144 13530
rect 374092 13466 374144 13472
rect 374104 3330 374132 13466
rect 375392 6914 375420 20130
rect 376036 16574 376064 59463
rect 376206 59256 376262 59265
rect 376206 59191 376262 59200
rect 376220 31210 376248 59191
rect 376760 54800 376812 54806
rect 376760 54742 376812 54748
rect 376208 31204 376260 31210
rect 376208 31146 376260 31152
rect 376772 16574 376800 54742
rect 376036 16546 376156 16574
rect 376772 16546 377352 16574
rect 375392 6886 376064 6914
rect 374092 3324 374144 3330
rect 374092 3266 374144 3272
rect 375288 3324 375340 3330
rect 375288 3266 375340 3272
rect 374012 3182 374132 3210
rect 374104 480 374132 3182
rect 375300 480 375328 3266
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 6886
rect 376128 4894 376156 16546
rect 376116 4888 376168 4894
rect 376116 4830 376168 4836
rect 377324 3482 377352 16546
rect 377416 4962 377444 59570
rect 378520 59401 378548 59599
rect 378506 59392 378562 59401
rect 378506 59327 378562 59336
rect 378782 59256 378838 59265
rect 378782 59191 378838 59200
rect 378416 13456 378468 13462
rect 378416 13398 378468 13404
rect 377404 4956 377456 4962
rect 377404 4898 377456 4904
rect 377324 3454 377720 3482
rect 377692 480 377720 3454
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 13398
rect 378796 5098 378824 59191
rect 378784 5092 378836 5098
rect 378784 5034 378836 5040
rect 378980 5030 379008 59706
rect 379440 59537 379468 59706
rect 379426 59528 379482 59537
rect 379426 59463 379482 59472
rect 379520 40928 379572 40934
rect 379520 40870 379572 40876
rect 378968 5024 379020 5030
rect 378968 4966 379020 4972
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 379532 354 379560 40870
rect 380176 28490 380204 59706
rect 380990 59664 381046 59673
rect 380990 59599 381046 59608
rect 380806 59392 380862 59401
rect 380806 59327 380862 59336
rect 380820 56166 380848 59327
rect 380808 56160 380860 56166
rect 380808 56102 380860 56108
rect 381004 55214 381032 59599
rect 382292 57526 382320 59706
rect 382280 57520 382332 57526
rect 382280 57462 382332 57468
rect 381004 55186 381584 55214
rect 380900 50652 380952 50658
rect 380900 50594 380952 50600
rect 380164 28484 380216 28490
rect 380164 28426 380216 28432
rect 380912 16574 380940 50594
rect 381556 27198 381584 55186
rect 382280 40996 382332 41002
rect 382280 40938 382332 40944
rect 381544 27192 381596 27198
rect 381544 27134 381596 27140
rect 380912 16546 381216 16574
rect 381188 480 381216 16546
rect 382292 3210 382320 40938
rect 382936 25770 382964 59774
rect 390006 59800 390062 59809
rect 387522 59735 387524 59744
rect 387576 59735 387578 59744
rect 389824 59764 389876 59770
rect 387524 59706 387576 59712
rect 390006 59735 390062 59744
rect 390834 59800 390890 59809
rect 390834 59735 390890 59744
rect 391662 59800 391718 59809
rect 397458 59800 397514 59809
rect 391662 59735 391664 59744
rect 389824 59706 389876 59712
rect 383198 59664 383254 59673
rect 383198 59599 383254 59608
rect 385866 59664 385922 59673
rect 385866 59599 385922 59608
rect 383212 59401 383240 59599
rect 383474 59528 383530 59537
rect 383530 59486 383700 59514
rect 383474 59463 383530 59472
rect 383198 59392 383254 59401
rect 383198 59327 383254 59336
rect 383672 58954 383700 59486
rect 385880 59401 385908 59599
rect 387246 59528 387302 59537
rect 387246 59463 387302 59472
rect 384118 59392 384174 59401
rect 385866 59392 385922 59401
rect 384118 59327 384120 59336
rect 384172 59327 384174 59336
rect 385684 59356 385736 59362
rect 384120 59298 384172 59304
rect 385866 59327 385922 59336
rect 385684 59298 385736 59304
rect 384302 59256 384358 59265
rect 384302 59191 384358 59200
rect 383660 58948 383712 58954
rect 383660 58890 383712 58896
rect 382924 25764 382976 25770
rect 382924 25706 382976 25712
rect 384316 24478 384344 59191
rect 384304 24472 384356 24478
rect 384304 24414 384356 24420
rect 385696 20126 385724 59298
rect 387062 59256 387118 59265
rect 387062 59191 387118 59200
rect 386420 56092 386472 56098
rect 386420 56034 386472 56040
rect 382372 20120 382424 20126
rect 382372 20062 382424 20068
rect 385684 20120 385736 20126
rect 385684 20062 385736 20068
rect 382384 3330 382412 20062
rect 386432 16574 386460 56034
rect 387076 40934 387104 59191
rect 387260 46510 387288 59463
rect 388626 59392 388682 59401
rect 388626 59327 388682 59336
rect 388442 59256 388498 59265
rect 388442 59191 388498 59200
rect 387248 46504 387300 46510
rect 387248 46446 387300 46452
rect 387064 40928 387116 40934
rect 387064 40870 387116 40876
rect 388456 20194 388484 59191
rect 388640 45014 388668 59327
rect 388628 45008 388680 45014
rect 388628 44950 388680 44956
rect 389836 23050 389864 59706
rect 390020 59702 390048 59735
rect 390008 59696 390060 59702
rect 390008 59638 390060 59644
rect 390006 59528 390062 59537
rect 390006 59463 390062 59472
rect 390020 43654 390048 59463
rect 390848 59401 390876 59735
rect 391716 59735 391718 59744
rect 393964 59764 394016 59770
rect 391664 59706 391716 59712
rect 402334 59800 402390 59809
rect 397458 59735 397460 59744
rect 393964 59706 394016 59712
rect 397512 59735 397514 59744
rect 399484 59764 399536 59770
rect 397460 59706 397512 59712
rect 406474 59800 406530 59809
rect 402334 59735 402336 59744
rect 399484 59706 399536 59712
rect 402388 59735 402390 59744
rect 404452 59764 404504 59770
rect 402336 59706 402388 59712
rect 410614 59800 410670 59809
rect 406474 59735 406476 59744
rect 404452 59706 404504 59712
rect 406528 59735 406530 59744
rect 408500 59764 408552 59770
rect 406476 59706 406528 59712
rect 416870 59800 416926 59809
rect 410614 59735 410616 59744
rect 408500 59706 408552 59712
rect 410668 59735 410670 59744
rect 412824 59764 412876 59770
rect 410616 59706 410668 59712
rect 416870 59735 416926 59744
rect 419538 59800 419594 59809
rect 419538 59735 419594 59744
rect 425518 59800 425574 59809
rect 427082 59800 427138 59809
rect 425518 59735 425520 59744
rect 412824 59706 412876 59712
rect 392584 59696 392636 59702
rect 391202 59664 391258 59673
rect 392584 59638 392636 59644
rect 393318 59664 393374 59673
rect 391202 59599 391258 59608
rect 390834 59392 390890 59401
rect 390834 59327 390890 59336
rect 390008 43648 390060 43654
rect 390008 43590 390060 43596
rect 391216 35494 391244 59599
rect 391204 35488 391256 35494
rect 391204 35430 391256 35436
rect 389824 23044 389876 23050
rect 389824 22986 389876 22992
rect 388444 20188 388496 20194
rect 388444 20130 388496 20136
rect 390560 19984 390612 19990
rect 390560 19926 390612 19932
rect 386432 16546 386736 16574
rect 385960 13388 386012 13394
rect 385960 13330 386012 13336
rect 384304 13184 384356 13190
rect 384304 13126 384356 13132
rect 382372 3324 382424 3330
rect 382372 3266 382424 3272
rect 383568 3324 383620 3330
rect 383568 3266 383620 3272
rect 382292 3182 382412 3210
rect 382384 480 382412 3182
rect 383580 480 383608 3266
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 378846 -960 378958 326
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 13126
rect 385972 480 386000 13330
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 386708 354 386736 16546
rect 387800 13388 387852 13394
rect 387800 13330 387852 13336
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 13330
rect 389456 13320 389508 13326
rect 389456 13262 389508 13268
rect 389468 480 389496 13262
rect 390572 3210 390600 19926
rect 390652 13320 390704 13326
rect 390652 13262 390704 13268
rect 390664 3330 390692 13262
rect 392492 13252 392544 13258
rect 392492 13194 392544 13200
rect 392504 6914 392532 13194
rect 392596 11830 392624 59638
rect 393318 59599 393320 59608
rect 393372 59599 393374 59608
rect 393320 59570 393372 59576
rect 393318 59528 393374 59537
rect 393686 59528 393742 59537
rect 393374 59486 393686 59514
rect 393318 59463 393374 59472
rect 393686 59463 393742 59472
rect 392766 59392 392822 59401
rect 392766 59327 392822 59336
rect 392780 42226 392808 59327
rect 393320 57452 393372 57458
rect 393320 57394 393372 57400
rect 392768 42220 392820 42226
rect 392768 42162 392820 42168
rect 392584 11824 392636 11830
rect 392584 11766 392636 11772
rect 393332 6914 393360 57394
rect 393976 13122 394004 59706
rect 395802 59664 395858 59673
rect 395344 59628 395396 59634
rect 395802 59599 395858 59608
rect 397458 59664 397514 59673
rect 397826 59664 397882 59673
rect 397514 59622 397826 59650
rect 397458 59599 397514 59608
rect 397826 59599 397882 59608
rect 398286 59664 398342 59673
rect 398286 59599 398342 59608
rect 395344 59570 395396 59576
rect 394146 59528 394202 59537
rect 394146 59463 394202 59472
rect 394160 38146 394188 59463
rect 394700 49360 394752 49366
rect 394700 49302 394752 49308
rect 394148 38140 394200 38146
rect 394148 38082 394200 38088
rect 394712 16574 394740 49302
rect 395356 39574 395384 59570
rect 395816 59401 395844 59599
rect 396722 59528 396778 59537
rect 396722 59463 396778 59472
rect 398102 59528 398158 59537
rect 398102 59463 398104 59472
rect 395802 59392 395858 59401
rect 395802 59327 395858 59336
rect 395344 39568 395396 39574
rect 395344 39510 395396 39516
rect 396080 32768 396132 32774
rect 396080 32710 396132 32716
rect 394712 16546 395384 16574
rect 393964 13116 394016 13122
rect 393964 13058 394016 13064
rect 392504 6886 392624 6914
rect 393332 6886 394280 6914
rect 390652 3324 390704 3330
rect 390652 3266 390704 3272
rect 391848 3324 391900 3330
rect 391848 3266 391900 3272
rect 390572 3182 390692 3210
rect 390664 480 390692 3182
rect 391860 480 391888 3266
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 6886
rect 394252 480 394280 6886
rect 395356 480 395384 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 32710
rect 396736 12034 396764 59463
rect 398156 59463 398158 59472
rect 398104 59434 398156 59440
rect 398010 59392 398066 59401
rect 398010 59327 398066 59336
rect 396906 59256 396962 59265
rect 396906 59191 396962 59200
rect 396920 30054 396948 59191
rect 398024 55214 398052 59327
rect 398024 55186 398144 55214
rect 396908 30048 396960 30054
rect 396908 29990 396960 29996
rect 397460 21616 397512 21622
rect 397460 21558 397512 21564
rect 397472 16574 397500 21558
rect 398116 19990 398144 55186
rect 398300 47870 398328 59599
rect 398840 52080 398892 52086
rect 398840 52022 398892 52028
rect 398288 47864 398340 47870
rect 398288 47806 398340 47812
rect 398104 19984 398156 19990
rect 398104 19926 398156 19932
rect 397472 16546 397776 16574
rect 396724 12028 396776 12034
rect 396724 11970 396776 11976
rect 397748 480 397776 16546
rect 398852 3330 398880 52022
rect 398932 20664 398984 20670
rect 398932 20606 398984 20612
rect 398840 3324 398892 3330
rect 398840 3266 398892 3272
rect 398944 480 398972 20606
rect 399496 13258 399524 59706
rect 399942 59664 399998 59673
rect 399942 59599 399998 59608
rect 400770 59664 400826 59673
rect 400770 59599 400826 59608
rect 399956 59401 399984 59599
rect 400784 59401 400812 59599
rect 400862 59528 400918 59537
rect 400862 59463 400918 59472
rect 401048 59492 401100 59498
rect 399942 59392 399998 59401
rect 399942 59327 399998 59336
rect 400770 59392 400826 59401
rect 400770 59327 400826 59336
rect 400220 27124 400272 27130
rect 400220 27066 400272 27072
rect 399484 13252 399536 13258
rect 399484 13194 399536 13200
rect 400232 6914 400260 27066
rect 400876 12102 400904 59463
rect 401048 59434 401100 59440
rect 401060 13462 401088 59434
rect 401598 59392 401654 59401
rect 401598 59327 401654 59336
rect 403070 59392 403126 59401
rect 403070 59327 403126 59336
rect 401612 59022 401640 59327
rect 402242 59256 402298 59265
rect 402242 59191 402298 59200
rect 401600 59016 401652 59022
rect 401600 58958 401652 58964
rect 402256 23118 402284 59191
rect 402980 34060 403032 34066
rect 402980 34002 403032 34008
rect 402244 23112 402296 23118
rect 402244 23054 402296 23060
rect 401048 13456 401100 13462
rect 401048 13398 401100 13404
rect 400864 12096 400916 12102
rect 400864 12038 400916 12044
rect 400232 6886 400904 6914
rect 400128 3324 400180 3330
rect 400128 3266 400180 3272
rect 400140 480 400168 3266
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 6886
rect 402992 5794 403020 34002
rect 403084 5914 403112 59327
rect 404358 59256 404414 59265
rect 404358 59191 404414 59200
rect 404372 49366 404400 59191
rect 404360 49360 404412 49366
rect 404360 49302 404412 49308
rect 404360 36644 404412 36650
rect 404360 36586 404412 36592
rect 403072 5908 403124 5914
rect 403072 5850 403124 5856
rect 402992 5766 403664 5794
rect 402980 5704 403032 5710
rect 402900 5652 402980 5658
rect 402900 5646 403032 5652
rect 402900 5630 403020 5646
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 354 402602 480
rect 402900 354 402928 5630
rect 403636 480 403664 5766
rect 402490 326 402928 354
rect 402490 -960 402602 326
rect 403594 -960 403706 480
rect 404372 354 404400 36586
rect 404464 20670 404492 59706
rect 405922 59528 405978 59537
rect 405922 59463 405978 59472
rect 408130 59528 408186 59537
rect 408130 59463 408132 59472
rect 405740 59016 405792 59022
rect 405740 58958 405792 58964
rect 404452 20664 404504 20670
rect 404452 20606 404504 20612
rect 405752 6914 405780 58958
rect 405936 13394 405964 59463
rect 408184 59463 408186 59472
rect 408132 59434 408184 59440
rect 406106 59392 406162 59401
rect 406106 59327 406162 59336
rect 405924 13388 405976 13394
rect 405924 13330 405976 13336
rect 406120 13326 406148 59327
rect 407302 59256 407358 59265
rect 407302 59191 407358 59200
rect 407120 46436 407172 46442
rect 407120 46378 407172 46384
rect 406108 13320 406160 13326
rect 406108 13262 406160 13268
rect 405752 6886 406056 6914
rect 406028 480 406056 6886
rect 407132 3210 407160 46378
rect 407212 24336 407264 24342
rect 407212 24278 407264 24284
rect 407224 3330 407252 24278
rect 407316 13190 407344 59191
rect 408512 50658 408540 59706
rect 412086 59664 412142 59673
rect 412086 59599 412142 59608
rect 409970 59528 410026 59537
rect 409880 59492 409932 59498
rect 409970 59463 410026 59472
rect 409880 59434 409932 59440
rect 408682 59392 408738 59401
rect 408682 59327 408738 59336
rect 408696 54806 408724 59327
rect 408684 54800 408736 54806
rect 408684 54742 408736 54748
rect 408500 50652 408552 50658
rect 408500 50594 408552 50600
rect 409892 31346 409920 59434
rect 409880 31340 409932 31346
rect 409880 31282 409932 31288
rect 408500 23112 408552 23118
rect 408500 23054 408552 23060
rect 408512 16574 408540 23054
rect 408512 16546 409184 16574
rect 407304 13184 407356 13190
rect 407304 13126 407356 13132
rect 407212 3324 407264 3330
rect 407212 3266 407264 3272
rect 408408 3324 408460 3330
rect 408408 3266 408460 3272
rect 407132 3182 407252 3210
rect 407224 480 407252 3182
rect 408420 480 408448 3266
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 409984 10674 410012 59463
rect 412100 59401 412128 59599
rect 412730 59528 412786 59537
rect 412730 59463 412786 59472
rect 411350 59392 411406 59401
rect 411350 59327 411406 59336
rect 412086 59392 412142 59401
rect 412086 59327 412142 59336
rect 411260 49088 411312 49094
rect 411260 49030 411312 49036
rect 410064 36916 410116 36922
rect 410064 36858 410116 36864
rect 410076 16574 410104 36858
rect 410076 16546 410840 16574
rect 409972 10668 410024 10674
rect 409972 10610 410024 10616
rect 410812 480 410840 16546
rect 411272 6914 411300 49030
rect 411364 11966 411392 59327
rect 412640 12096 412692 12102
rect 412640 12038 412692 12044
rect 411352 11960 411404 11966
rect 411352 11902 411404 11908
rect 411272 6886 411944 6914
rect 411916 480 411944 6886
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 12038
rect 412744 10538 412772 59463
rect 412836 55214 412864 59706
rect 413098 59664 413154 59673
rect 416410 59664 416466 59673
rect 413098 59599 413100 59608
rect 413152 59599 413154 59608
rect 414112 59628 414164 59634
rect 413100 59570 413152 59576
rect 416410 59599 416412 59608
rect 414112 59570 414164 59576
rect 416464 59599 416466 59608
rect 416412 59570 416464 59576
rect 412914 59528 412970 59537
rect 412914 59463 412970 59472
rect 412928 56234 412956 59463
rect 413926 59392 413982 59401
rect 413982 59350 414060 59378
rect 413926 59327 413982 59336
rect 412916 56228 412968 56234
rect 412916 56170 412968 56176
rect 412836 55186 412956 55214
rect 412928 10606 412956 55186
rect 412916 10600 412968 10606
rect 412916 10542 412968 10548
rect 412732 10532 412784 10538
rect 412732 10474 412784 10480
rect 414032 10470 414060 59350
rect 414020 10464 414072 10470
rect 414020 10406 414072 10412
rect 414124 10402 414152 59570
rect 416778 59528 416834 59537
rect 416778 59463 416834 59472
rect 415400 47592 415452 47598
rect 415400 47534 415452 47540
rect 414296 16312 414348 16318
rect 414296 16254 414348 16260
rect 414112 10396 414164 10402
rect 414112 10338 414164 10344
rect 414308 480 414336 16254
rect 415412 3210 415440 47534
rect 416792 20330 416820 59463
rect 416884 57594 416912 59735
rect 418252 59628 418304 59634
rect 418252 59570 418304 59576
rect 416962 59392 417018 59401
rect 416962 59327 417018 59336
rect 418158 59392 418214 59401
rect 418158 59327 418214 59336
rect 416872 57588 416924 57594
rect 416872 57530 416924 57536
rect 416780 20324 416832 20330
rect 416780 20266 416832 20272
rect 415492 13456 415544 13462
rect 415492 13398 415544 13404
rect 415504 3330 415532 13398
rect 416976 10334 417004 59327
rect 418172 28558 418200 59327
rect 418160 28552 418212 28558
rect 418160 28494 418212 28500
rect 417424 16244 417476 16250
rect 417424 16186 417476 16192
rect 416964 10328 417016 10334
rect 416964 10270 417016 10276
rect 415492 3324 415544 3330
rect 415492 3266 415544 3272
rect 416688 3324 416740 3330
rect 416688 3266 416740 3272
rect 415412 3182 415532 3210
rect 415504 480 415532 3182
rect 416700 480 416728 3266
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16186
rect 418264 11898 418292 59570
rect 419552 58886 419580 59735
rect 425572 59735 425574 59744
rect 426532 59764 426584 59770
rect 425520 59706 425572 59712
rect 431222 59800 431278 59809
rect 427082 59735 427084 59744
rect 426532 59706 426584 59712
rect 427136 59735 427138 59744
rect 429568 59764 429620 59770
rect 427084 59706 427136 59712
rect 435454 59800 435510 59809
rect 431222 59735 431224 59744
rect 429568 59706 429620 59712
rect 431276 59735 431278 59744
rect 433616 59764 433668 59770
rect 431224 59706 431276 59712
rect 436926 59800 436982 59809
rect 435510 59758 435680 59786
rect 435454 59735 435510 59744
rect 433616 59706 433668 59712
rect 420918 59664 420974 59673
rect 420918 59599 420974 59608
rect 419540 58880 419592 58886
rect 419540 58822 419592 58828
rect 418344 29776 418396 29782
rect 418344 29718 418396 29724
rect 418356 16574 418384 29718
rect 420932 25838 420960 59599
rect 425334 59528 425390 59537
rect 425334 59463 425390 59472
rect 422390 59392 422446 59401
rect 422390 59327 422446 59336
rect 425150 59392 425206 59401
rect 425150 59327 425206 59336
rect 421102 59256 421158 59265
rect 421102 59191 421158 59200
rect 421116 27266 421144 59191
rect 422300 51876 422352 51882
rect 422300 51818 422352 51824
rect 421104 27260 421156 27266
rect 421104 27202 421156 27208
rect 420920 25832 420972 25838
rect 420920 25774 420972 25780
rect 422312 16574 422340 51818
rect 422404 24410 422432 59327
rect 423770 59256 423826 59265
rect 423770 59191 423826 59200
rect 423680 47864 423732 47870
rect 423680 47806 423732 47812
rect 422392 24404 422444 24410
rect 422392 24346 422444 24352
rect 418356 16546 418568 16574
rect 422312 16546 422616 16574
rect 418252 11892 418304 11898
rect 418252 11834 418304 11840
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 420920 16176 420972 16182
rect 420920 16118 420972 16124
rect 420184 13252 420236 13258
rect 420184 13194 420236 13200
rect 420196 480 420224 13194
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 16118
rect 422588 480 422616 16546
rect 423692 3210 423720 47806
rect 423784 39642 423812 59191
rect 423772 39636 423824 39642
rect 423772 39578 423824 39584
rect 423772 16108 423824 16114
rect 423772 16050 423824 16056
rect 423784 3330 423812 16050
rect 425164 9382 425192 59327
rect 425152 9376 425204 9382
rect 425152 9318 425204 9324
rect 425348 9314 425376 59463
rect 426438 59256 426494 59265
rect 426438 59191 426494 59200
rect 426452 38214 426480 59191
rect 426544 42362 426572 59706
rect 428738 59528 428794 59537
rect 428738 59463 428740 59472
rect 428792 59463 428794 59472
rect 428740 59434 428792 59440
rect 429382 59392 429438 59401
rect 429382 59327 429438 59336
rect 427910 59256 427966 59265
rect 427910 59191 427966 59200
rect 426532 42356 426584 42362
rect 426532 42298 426584 42304
rect 426440 38208 426492 38214
rect 426440 38150 426492 38156
rect 426440 19984 426492 19990
rect 426440 19926 426492 19932
rect 426452 16574 426480 19926
rect 426452 16546 426848 16574
rect 425704 11756 425756 11762
rect 425704 11698 425756 11704
rect 425336 9308 425388 9314
rect 425336 9250 425388 9256
rect 423772 3324 423824 3330
rect 423772 3266 423824 3272
rect 424968 3324 425020 3330
rect 424968 3266 425020 3272
rect 423692 3182 423812 3210
rect 423784 480 423812 3182
rect 424980 480 425008 3266
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 11698
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 16546
rect 427924 9246 427952 59191
rect 429200 21548 429252 21554
rect 429200 21490 429252 21496
rect 428464 16040 428516 16046
rect 428464 15982 428516 15988
rect 427912 9240 427964 9246
rect 427912 9182 427964 9188
rect 428476 480 428504 15982
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429212 354 429240 21490
rect 429396 9110 429424 59327
rect 429580 9178 429608 59706
rect 430578 59528 430634 59537
rect 432050 59528 432106 59537
rect 430578 59463 430634 59472
rect 430672 59492 430724 59498
rect 429568 9172 429620 9178
rect 429568 9114 429620 9120
rect 429384 9104 429436 9110
rect 429384 9046 429436 9052
rect 430592 8974 430620 59463
rect 432050 59463 432052 59472
rect 430672 59434 430724 59440
rect 432104 59463 432106 59472
rect 433432 59492 433484 59498
rect 432052 59434 432104 59440
rect 433432 59434 433484 59440
rect 430684 9042 430712 59434
rect 432050 59392 432106 59401
rect 432050 59327 432106 59336
rect 431960 43580 432012 43586
rect 431960 43522 432012 43528
rect 430856 12028 430908 12034
rect 430856 11970 430908 11976
rect 430672 9036 430724 9042
rect 430672 8978 430724 8984
rect 430580 8968 430632 8974
rect 430580 8910 430632 8916
rect 430868 480 430896 11970
rect 431972 3330 432000 43522
rect 432064 35426 432092 59327
rect 433444 43722 433472 59434
rect 433432 43716 433484 43722
rect 433432 43658 433484 43664
rect 432052 35420 432104 35426
rect 432052 35362 432104 35368
rect 433340 30048 433392 30054
rect 433340 29990 433392 29996
rect 433352 16574 433380 29990
rect 433628 29918 433656 59706
rect 435652 59537 435680 59758
rect 440238 59800 440294 59809
rect 436926 59735 436928 59744
rect 436980 59735 436982 59744
rect 439228 59764 439280 59770
rect 436928 59706 436980 59712
rect 440238 59735 440294 59744
rect 441158 59800 441214 59809
rect 441434 59800 441490 59809
rect 441214 59758 441434 59786
rect 441158 59735 441214 59744
rect 441434 59735 441490 59744
rect 441894 59800 441950 59809
rect 445942 59800 445998 59809
rect 441894 59735 441896 59744
rect 439228 59706 439280 59712
rect 438582 59664 438638 59673
rect 438582 59599 438638 59608
rect 434718 59528 434774 59537
rect 434718 59463 434774 59472
rect 435638 59528 435694 59537
rect 435638 59463 435694 59472
rect 436374 59528 436430 59537
rect 436374 59463 436430 59472
rect 434732 51950 434760 59463
rect 434902 59392 434958 59401
rect 434902 59327 434958 59336
rect 434720 51944 434772 51950
rect 434720 51886 434772 51892
rect 434720 45076 434772 45082
rect 434720 45018 434772 45024
rect 433616 29912 433668 29918
rect 433616 29854 433668 29860
rect 434732 16574 434760 45018
rect 434916 22982 434944 59327
rect 436190 59256 436246 59265
rect 436190 59191 436246 59200
rect 436204 53174 436232 59191
rect 436192 53168 436244 53174
rect 436192 53110 436244 53116
rect 436388 49230 436416 59463
rect 438596 59401 438624 59599
rect 439042 59528 439098 59537
rect 439042 59463 439098 59472
rect 437478 59392 437534 59401
rect 437478 59327 437534 59336
rect 438582 59392 438638 59401
rect 438582 59327 438638 59336
rect 437492 54670 437520 59327
rect 437480 54664 437532 54670
rect 437480 54606 437532 54612
rect 438860 49292 438912 49298
rect 438860 49234 438912 49240
rect 436376 49224 436428 49230
rect 436376 49166 436428 49172
rect 437480 39568 437532 39574
rect 437480 39510 437532 39516
rect 434904 22976 434956 22982
rect 434904 22918 434956 22924
rect 436100 21480 436152 21486
rect 436100 21422 436152 21428
rect 436112 16574 436140 21422
rect 433352 16546 434024 16574
rect 434732 16546 435128 16574
rect 436112 16546 436784 16574
rect 432052 15972 432104 15978
rect 432052 15914 432104 15920
rect 431960 3324 432012 3330
rect 431960 3266 432012 3272
rect 432064 480 432092 15914
rect 433248 3324 433300 3330
rect 433248 3266 433300 3272
rect 433260 480 433288 3266
rect 429630 354 429742 480
rect 429212 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 16546
rect 436756 480 436784 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 39510
rect 438872 6914 438900 49234
rect 439056 7954 439084 59463
rect 439240 8022 439268 59706
rect 440252 59401 440280 59735
rect 441948 59735 441950 59744
rect 443184 59764 443236 59770
rect 441896 59706 441948 59712
rect 445942 59735 445998 59744
rect 446862 59800 446918 59809
rect 449346 59800 449402 59809
rect 446862 59735 446864 59744
rect 443184 59706 443236 59712
rect 440422 59664 440478 59673
rect 440422 59599 440478 59608
rect 440238 59392 440294 59401
rect 440238 59327 440294 59336
rect 440238 59256 440294 59265
rect 440238 59191 440294 59200
rect 440252 47802 440280 59191
rect 440240 47796 440292 47802
rect 440240 47738 440292 47744
rect 440240 38140 440292 38146
rect 440240 38082 440292 38088
rect 439228 8016 439280 8022
rect 439228 7958 439280 7964
rect 439044 7948 439096 7954
rect 439044 7890 439096 7896
rect 438872 6886 439176 6914
rect 439148 480 439176 6886
rect 440252 3330 440280 38082
rect 440332 32564 440384 32570
rect 440332 32506 440384 32512
rect 440240 3324 440292 3330
rect 440240 3266 440292 3272
rect 440344 480 440372 32506
rect 440436 7886 440464 59599
rect 441710 59256 441766 59265
rect 441710 59191 441766 59200
rect 440424 7880 440476 7886
rect 440424 7822 440476 7828
rect 441724 7818 441752 59191
rect 443000 21412 443052 21418
rect 443000 21354 443052 21360
rect 442632 15904 442684 15910
rect 442632 15846 442684 15852
rect 441712 7812 441764 7818
rect 441712 7754 441764 7760
rect 441528 3324 441580 3330
rect 441528 3266 441580 3272
rect 441540 480 441568 3266
rect 442644 480 442672 15846
rect 443012 6914 443040 21354
rect 443196 7750 443224 59706
rect 445850 59664 445906 59673
rect 445850 59599 445906 59608
rect 444378 59528 444434 59537
rect 444378 59463 444434 59472
rect 443366 59256 443422 59265
rect 443366 59191 443422 59200
rect 443184 7744 443236 7750
rect 443184 7686 443236 7692
rect 443380 7682 443408 59191
rect 444392 44878 444420 59463
rect 444470 59392 444526 59401
rect 444470 59327 444526 59336
rect 444484 46306 444512 59327
rect 445760 53304 445812 53310
rect 445760 53246 445812 53252
rect 444472 46300 444524 46306
rect 444472 46242 444524 46248
rect 444380 44872 444432 44878
rect 444380 44814 444432 44820
rect 445024 13116 445076 13122
rect 445024 13058 445076 13064
rect 443368 7676 443420 7682
rect 443368 7618 443420 7624
rect 443012 6886 443408 6914
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 6886
rect 445036 480 445064 13058
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 445772 354 445800 53246
rect 445864 36582 445892 59599
rect 445956 59401 445984 59735
rect 446916 59735 446918 59744
rect 448796 59764 448848 59770
rect 446864 59706 446916 59712
rect 449346 59735 449402 59744
rect 449714 59800 449770 59809
rect 449714 59735 449770 59744
rect 457534 59800 457590 59809
rect 461582 59800 461638 59809
rect 457534 59735 457536 59744
rect 448796 59706 448848 59712
rect 446862 59664 446918 59673
rect 446918 59622 447180 59650
rect 446862 59599 446918 59608
rect 445942 59392 445998 59401
rect 445942 59327 445998 59336
rect 447152 55962 447180 59622
rect 448610 59528 448666 59537
rect 448610 59463 448666 59472
rect 447414 59392 447470 59401
rect 447414 59327 447470 59336
rect 447140 55956 447192 55962
rect 447140 55898 447192 55904
rect 445852 36576 445904 36582
rect 445852 36518 445904 36524
rect 447428 33930 447456 59327
rect 448520 42220 448572 42226
rect 448520 42162 448572 42168
rect 447416 33924 447468 33930
rect 447416 33866 447468 33872
rect 447416 3392 447468 3398
rect 447416 3334 447468 3340
rect 447428 480 447456 3334
rect 448532 3210 448560 42162
rect 448624 31074 448652 59463
rect 448808 32638 448836 59706
rect 449254 59664 449310 59673
rect 449254 59599 449256 59608
rect 449308 59599 449310 59608
rect 449256 59570 449308 59576
rect 449360 59401 449388 59735
rect 449346 59392 449402 59401
rect 449346 59327 449402 59336
rect 449728 58750 449756 59735
rect 457588 59735 457590 59744
rect 459928 59764 459980 59770
rect 457536 59706 457588 59712
rect 461582 59735 461638 59744
rect 464158 59800 464214 59809
rect 464158 59735 464160 59744
rect 459928 59706 459980 59712
rect 453394 59664 453450 59673
rect 449900 59628 449952 59634
rect 453394 59599 453396 59608
rect 449900 59570 449952 59576
rect 453448 59599 453450 59608
rect 455696 59628 455748 59634
rect 453396 59570 453448 59576
rect 455696 59570 455748 59576
rect 449716 58744 449768 58750
rect 449716 58686 449768 58692
rect 448796 32632 448848 32638
rect 448796 32574 448848 32580
rect 448612 31068 448664 31074
rect 448612 31010 448664 31016
rect 449912 28354 449940 59570
rect 455050 59528 455106 59537
rect 455050 59463 455052 59472
rect 455104 59463 455106 59472
rect 455052 59434 455104 59440
rect 455510 59392 455566 59401
rect 455510 59327 455566 59336
rect 451278 59256 451334 59265
rect 451278 59191 451334 59200
rect 452750 59256 452806 59265
rect 452750 59191 452806 59200
rect 454038 59256 454094 59265
rect 454038 59191 454094 59200
rect 451292 57322 451320 59191
rect 451280 57316 451332 57322
rect 451280 57258 451332 57264
rect 452660 31272 452712 31278
rect 452660 31214 452712 31220
rect 449900 28348 449952 28354
rect 449900 28290 449952 28296
rect 448612 21684 448664 21690
rect 448612 21626 448664 21632
rect 448624 3398 448652 21626
rect 452672 16574 452700 31214
rect 452764 24206 452792 59191
rect 452934 59120 452990 59129
rect 452934 59055 452990 59064
rect 452948 25634 452976 59055
rect 454052 42090 454080 59191
rect 455524 43518 455552 59327
rect 455512 43512 455564 43518
rect 455512 43454 455564 43460
rect 454040 42084 454092 42090
rect 454040 42026 454092 42032
rect 455708 40798 455736 59570
rect 456798 59528 456854 59537
rect 459190 59528 459246 59537
rect 456798 59463 456854 59472
rect 456984 59492 457036 59498
rect 455696 40792 455748 40798
rect 455696 40734 455748 40740
rect 456812 38010 456840 59463
rect 459190 59463 459192 59472
rect 456984 59434 457036 59440
rect 459244 59463 459246 59472
rect 459192 59434 459244 59440
rect 456996 39370 457024 59434
rect 458270 59256 458326 59265
rect 458270 59191 458326 59200
rect 459742 59256 459798 59265
rect 459742 59191 459798 59200
rect 457076 50584 457128 50590
rect 457076 50526 457128 50532
rect 456984 39364 457036 39370
rect 456984 39306 457036 39312
rect 456800 38004 456852 38010
rect 456800 37946 456852 37952
rect 455420 35488 455472 35494
rect 455420 35430 455472 35436
rect 452936 25628 452988 25634
rect 452936 25570 452988 25576
rect 452752 24200 452804 24206
rect 452752 24142 452804 24148
rect 455432 16574 455460 35430
rect 452672 16546 453344 16574
rect 455432 16546 455736 16574
rect 451648 11824 451700 11830
rect 451648 11766 451700 11772
rect 450912 4140 450964 4146
rect 450912 4082 450964 4088
rect 448612 3392 448664 3398
rect 448612 3334 448664 3340
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 448532 3182 448652 3210
rect 448624 480 448652 3182
rect 449820 480 449848 3334
rect 450924 480 450952 4082
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 11766
rect 453316 480 453344 16546
rect 454500 4072 454552 4078
rect 454500 4014 454552 4020
rect 454512 480 454540 4014
rect 455708 480 455736 16546
rect 457088 6914 457116 50526
rect 458180 43648 458232 43654
rect 458180 43590 458232 43596
rect 458192 16574 458220 43590
rect 458284 35358 458312 59191
rect 459560 54732 459612 54738
rect 459560 54674 459612 54680
rect 458272 35352 458324 35358
rect 458272 35294 458324 35300
rect 459572 16574 459600 54674
rect 459756 33862 459784 59191
rect 459744 33856 459796 33862
rect 459744 33798 459796 33804
rect 459940 29646 459968 59706
rect 461216 59492 461268 59498
rect 461216 59434 461268 59440
rect 461030 59256 461086 59265
rect 461030 59191 461086 59200
rect 461044 49026 461072 59191
rect 461032 49020 461084 49026
rect 461032 48962 461084 48968
rect 461228 32502 461256 59434
rect 461596 59401 461624 59735
rect 464212 59735 464214 59744
rect 465356 59764 465408 59770
rect 464160 59706 464212 59712
rect 465356 59706 465408 59712
rect 461674 59664 461730 59673
rect 461730 59622 462360 59650
rect 461674 59599 461730 59608
rect 461582 59392 461638 59401
rect 461582 59327 461638 59336
rect 462332 53106 462360 59622
rect 463974 59528 464030 59537
rect 463974 59463 464030 59472
rect 463790 59392 463846 59401
rect 463790 59327 463846 59336
rect 462320 53100 462372 53106
rect 462320 53042 462372 53048
rect 463804 51814 463832 59327
rect 463792 51808 463844 51814
rect 463792 51750 463844 51756
rect 463988 40730 464016 59463
rect 465078 59256 465134 59265
rect 465078 59191 465134 59200
rect 465092 50386 465120 59191
rect 465080 50380 465132 50386
rect 465080 50322 465132 50328
rect 465264 45008 465316 45014
rect 465264 44950 465316 44956
rect 463976 40724 464028 40730
rect 463976 40666 464028 40672
rect 461216 32496 461268 32502
rect 461216 32438 461268 32444
rect 463700 29844 463752 29850
rect 463700 29786 463752 29792
rect 459928 29640 459980 29646
rect 459928 29582 459980 29588
rect 462320 23044 462372 23050
rect 462320 22986 462372 22992
rect 458192 16546 459232 16574
rect 459572 16546 459968 16574
rect 456904 6886 457116 6914
rect 456904 480 456932 6886
rect 458088 4004 458140 4010
rect 458088 3946 458140 3952
rect 458100 480 458128 3946
rect 459204 480 459232 16546
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 461584 3936 461636 3942
rect 461584 3878 461636 3884
rect 461596 480 461624 3878
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 22986
rect 463712 16574 463740 29786
rect 463712 16546 464016 16574
rect 463988 480 464016 16546
rect 465276 6914 465304 44950
rect 465368 7614 465396 59706
rect 467838 59528 467894 59537
rect 467838 59463 467894 59472
rect 466550 59392 466606 59401
rect 466550 59327 466606 59336
rect 466460 39500 466512 39506
rect 466460 39442 466512 39448
rect 466472 16574 466500 39442
rect 466564 26994 466592 59327
rect 466552 26988 466604 26994
rect 466552 26930 466604 26936
rect 467852 22846 467880 59463
rect 483020 58948 483072 58954
rect 483020 58890 483072 58896
rect 473360 46504 473412 46510
rect 473360 46446 473412 46452
rect 470600 40860 470652 40866
rect 470600 40802 470652 40808
rect 467840 22840 467892 22846
rect 467840 22782 467892 22788
rect 469220 20188 469272 20194
rect 469220 20130 469272 20136
rect 469232 16574 469260 20130
rect 466472 16546 467512 16574
rect 469232 16546 469904 16574
rect 465356 7608 465408 7614
rect 465356 7550 465408 7556
rect 465276 6886 465856 6914
rect 465172 3868 465224 3874
rect 465172 3810 465224 3816
rect 465184 480 465212 3810
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 354 465856 6886
rect 467484 480 467512 16546
rect 468668 3800 468720 3806
rect 468668 3742 468720 3748
rect 468680 480 468708 3742
rect 469876 480 469904 16546
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 354 470640 40802
rect 473372 6914 473400 46446
rect 476120 40928 476172 40934
rect 476120 40870 476172 40876
rect 473452 20052 473504 20058
rect 473452 19994 473504 20000
rect 473464 16574 473492 19994
rect 476132 16574 476160 40870
rect 481640 36712 481692 36718
rect 481640 36654 481692 36660
rect 480260 20120 480312 20126
rect 480260 20062 480312 20068
rect 477500 17808 477552 17814
rect 477500 17750 477552 17756
rect 477512 16574 477540 17750
rect 480272 16574 480300 20062
rect 473464 16546 474136 16574
rect 476132 16546 476528 16574
rect 477512 16546 478184 16574
rect 480272 16546 480576 16574
rect 473372 6886 473492 6914
rect 472256 3732 472308 3738
rect 472256 3674 472308 3680
rect 472268 480 472296 3674
rect 473464 480 473492 6886
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 16546
rect 475752 3664 475804 3670
rect 475752 3606 475804 3612
rect 475764 480 475792 3606
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 478156 480 478184 16546
rect 479340 3528 479392 3534
rect 479340 3470 479392 3476
rect 479352 480 479380 3470
rect 480548 480 480576 16546
rect 481652 6914 481680 36654
rect 481732 17740 481784 17746
rect 481732 17682 481784 17688
rect 481744 16574 481772 17682
rect 483032 16574 483060 58890
rect 513380 58812 513432 58818
rect 513380 58754 513432 58760
rect 489920 57520 489972 57526
rect 489920 57462 489972 57468
rect 488540 50448 488592 50454
rect 488540 50390 488592 50396
rect 484400 47660 484452 47666
rect 484400 47602 484452 47608
rect 484412 16574 484440 47602
rect 487160 24472 487212 24478
rect 487160 24414 487212 24420
rect 485780 17672 485832 17678
rect 485780 17614 485832 17620
rect 485792 16574 485820 17614
rect 481744 16546 482416 16574
rect 483032 16546 484072 16574
rect 484412 16546 484808 16574
rect 485792 16546 486464 16574
rect 481652 6886 481772 6914
rect 481744 480 481772 6886
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 354 482416 16546
rect 484044 480 484072 16546
rect 482806 354 482918 480
rect 482388 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 486436 480 486464 16546
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487172 354 487200 24414
rect 488552 16574 488580 50390
rect 488552 16546 488856 16574
rect 488828 480 488856 16546
rect 489932 3534 489960 57462
rect 506480 57384 506532 57390
rect 506480 57326 506532 57332
rect 500960 56160 501012 56166
rect 500960 56102 501012 56108
rect 495440 39432 495492 39438
rect 495440 39374 495492 39380
rect 491300 31136 491352 31142
rect 491300 31078 491352 31084
rect 490012 17604 490064 17610
rect 490012 17546 490064 17552
rect 489920 3528 489972 3534
rect 489920 3470 489972 3476
rect 490024 3346 490052 17546
rect 491312 16574 491340 31078
rect 494060 25764 494112 25770
rect 494060 25706 494112 25712
rect 492680 17536 492732 17542
rect 492680 17478 492732 17484
rect 492692 16574 492720 17478
rect 494072 16574 494100 25706
rect 491312 16546 492352 16574
rect 492692 16546 493088 16574
rect 494072 16546 494744 16574
rect 490748 3528 490800 3534
rect 490748 3470 490800 3476
rect 489932 3318 490052 3346
rect 489932 480 489960 3318
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490760 354 490788 3470
rect 492324 480 492352 16546
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494716 480 494744 16546
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 39374
rect 498200 38072 498252 38078
rect 498200 38014 498252 38020
rect 496820 17468 496872 17474
rect 496820 17410 496872 17416
rect 496832 16574 496860 17410
rect 496832 16546 497136 16574
rect 497108 480 497136 16546
rect 498212 3534 498240 38014
rect 498292 27192 498344 27198
rect 498292 27134 498344 27140
rect 498200 3528 498252 3534
rect 498200 3470 498252 3476
rect 498304 3346 498332 27134
rect 499580 17400 499632 17406
rect 499580 17342 499632 17348
rect 499592 16574 499620 17342
rect 500972 16574 501000 56102
rect 502340 56024 502392 56030
rect 502340 55966 502392 55972
rect 502352 16574 502380 55966
rect 505100 28484 505152 28490
rect 505100 28426 505152 28432
rect 503720 17332 503772 17338
rect 503720 17274 503772 17280
rect 499592 16546 500632 16574
rect 500972 16546 501368 16574
rect 502352 16546 503024 16574
rect 499028 3528 499080 3534
rect 499028 3470 499080 3476
rect 498212 3318 498332 3346
rect 498212 480 498240 3318
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499040 354 499068 3470
rect 500604 480 500632 16546
rect 499366 354 499478 480
rect 499040 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501340 354 501368 16546
rect 502996 480 503024 16546
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503732 354 503760 17274
rect 505112 16574 505140 28426
rect 505112 16546 505416 16574
rect 505388 480 505416 16546
rect 506492 480 506520 57326
rect 510620 37936 510672 37942
rect 510620 37878 510672 37884
rect 509240 28416 509292 28422
rect 509240 28358 509292 28364
rect 506572 17264 506624 17270
rect 506572 17206 506624 17212
rect 506584 16574 506612 17206
rect 509252 16574 509280 28358
rect 510632 16574 510660 37878
rect 506584 16546 507256 16574
rect 509252 16546 509648 16574
rect 510632 16546 511304 16574
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 354 507256 16546
rect 508872 5092 508924 5098
rect 508872 5034 508924 5040
rect 508884 480 508912 5034
rect 507646 354 507758 480
rect 507228 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 511276 480 511304 16546
rect 512460 5024 512512 5030
rect 512460 4966 512512 4972
rect 512472 480 512500 4966
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513392 354 513420 58754
rect 546500 58676 546552 58682
rect 546500 58618 546552 58624
rect 517520 57248 517572 57254
rect 517520 57190 517572 57196
rect 516140 42152 516192 42158
rect 516140 42094 516192 42100
rect 514760 35216 514812 35222
rect 514760 35158 514812 35164
rect 514772 480 514800 35158
rect 516152 16574 516180 42094
rect 517532 16574 517560 57190
rect 524420 55888 524472 55894
rect 524420 55830 524472 55836
rect 523040 31204 523092 31210
rect 523040 31146 523092 31152
rect 520280 25696 520332 25702
rect 520280 25638 520332 25644
rect 516152 16546 517192 16574
rect 517532 16546 517928 16574
rect 515956 4956 516008 4962
rect 515956 4898 516008 4904
rect 515968 480 515996 4898
rect 517164 480 517192 16546
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519544 4888 519596 4894
rect 519544 4830 519596 4836
rect 519556 480 519584 4830
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 25638
rect 521660 24132 521712 24138
rect 521660 24074 521712 24080
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 24074
rect 523052 480 523080 31146
rect 523132 24268 523184 24274
rect 523132 24210 523184 24216
rect 523144 16574 523172 24210
rect 524432 16574 524460 55830
rect 525800 54596 525852 54602
rect 525800 54538 525852 54544
rect 525812 16574 525840 54538
rect 532700 53236 532752 53242
rect 532700 53178 532752 53184
rect 528560 51740 528612 51746
rect 528560 51682 528612 51688
rect 527180 29708 527232 29714
rect 527180 29650 527232 29656
rect 527192 16574 527220 29650
rect 523144 16546 523816 16574
rect 524432 16546 525472 16574
rect 525812 16546 526208 16574
rect 527192 16546 527864 16574
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523788 354 523816 16546
rect 525444 480 525472 16546
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527836 480 527864 16546
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 51682
rect 529940 32700 529992 32706
rect 529940 32642 529992 32648
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 32642
rect 531320 27056 531372 27062
rect 531320 26998 531372 27004
rect 531332 480 531360 26998
rect 531412 25560 531464 25566
rect 531412 25502 531464 25508
rect 531424 16574 531452 25502
rect 532712 16574 532740 53178
rect 539600 52012 539652 52018
rect 539600 51954 539652 51960
rect 535460 22772 535512 22778
rect 535460 22714 535512 22720
rect 535472 16574 535500 22714
rect 531424 16546 532096 16574
rect 532712 16546 533752 16574
rect 535472 16546 536144 16574
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532068 354 532096 16546
rect 533724 480 533752 16546
rect 534448 15020 534500 15026
rect 534448 14962 534500 14968
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 14962
rect 536116 480 536144 16546
rect 538220 14952 538272 14958
rect 538220 14894 538272 14900
rect 537208 4820 537260 4826
rect 537208 4762 537260 4768
rect 537220 480 537248 4762
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 14894
rect 539612 3534 539640 51954
rect 543740 50516 543792 50522
rect 543740 50458 543792 50464
rect 539692 32428 539744 32434
rect 539692 32370 539744 32376
rect 539600 3528 539652 3534
rect 539600 3470 539652 3476
rect 539704 3346 539732 32370
rect 542360 18964 542412 18970
rect 542360 18906 542412 18912
rect 542372 16574 542400 18906
rect 543752 16574 543780 50458
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 541992 14884 542044 14890
rect 541992 14826 542044 14832
rect 540428 3528 540480 3534
rect 540428 3470 540480 3476
rect 539612 3318 539732 3346
rect 539612 480 539640 3318
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540440 354 540468 3470
rect 542004 480 542032 14826
rect 540766 354 540878 480
rect 540440 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545488 14816 545540 14822
rect 545488 14758 545540 14764
rect 545500 480 545528 14758
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 58618
rect 572720 54528 572772 54534
rect 572720 54470 572772 54476
rect 550640 49156 550692 49162
rect 550640 49098 550692 49104
rect 548524 46232 548576 46238
rect 548524 46174 548576 46180
rect 547880 33992 547932 33998
rect 547880 33934 547932 33940
rect 547892 480 547920 33934
rect 548432 14748 548484 14754
rect 548432 14690 548484 14696
rect 548444 490 548472 14690
rect 548536 3534 548564 46174
rect 550652 16574 550680 49098
rect 554780 47728 554832 47734
rect 554780 47670 554832 47676
rect 553400 18896 553452 18902
rect 553400 18838 553452 18844
rect 553412 16574 553440 18838
rect 550652 16546 551048 16574
rect 553412 16546 553808 16574
rect 548524 3528 548576 3534
rect 548524 3470 548576 3476
rect 550272 3528 550324 3534
rect 550272 3470 550324 3476
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548444 462 548656 490
rect 550284 480 550312 3470
rect 548628 354 548656 462
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 552664 14680 552716 14686
rect 552664 14622 552716 14628
rect 552676 480 552704 14622
rect 553780 480 553808 16546
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 47670
rect 561680 46368 561732 46374
rect 561680 46310 561732 46316
rect 557540 36780 557592 36786
rect 557540 36722 557592 36728
rect 556160 18828 556212 18834
rect 556160 18770 556212 18776
rect 556172 3534 556200 18770
rect 557552 16574 557580 36722
rect 560300 18760 560352 18766
rect 560300 18702 560352 18708
rect 560312 16574 560340 18702
rect 561692 16574 561720 46310
rect 564440 44940 564492 44946
rect 564440 44882 564492 44888
rect 557552 16546 558592 16574
rect 560312 16546 560432 16574
rect 561692 16546 562088 16574
rect 556252 14612 556304 14618
rect 556252 14554 556304 14560
rect 556160 3528 556212 3534
rect 556160 3470 556212 3476
rect 556264 3346 556292 14554
rect 556988 3528 557040 3534
rect 556988 3470 557040 3476
rect 556172 3318 556292 3346
rect 556172 480 556200 3318
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 557000 354 557028 3470
rect 558564 480 558592 16546
rect 559288 14544 559340 14550
rect 559288 14486 559340 14492
rect 557326 354 557438 480
rect 557000 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 14486
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 562060 480 562088 16546
rect 563060 14476 563112 14482
rect 563060 14418 563112 14424
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 14418
rect 564452 3534 564480 44882
rect 569960 43444 570012 43450
rect 569960 43386 570012 43392
rect 565820 35284 565872 35290
rect 565820 35226 565872 35232
rect 564532 33788 564584 33794
rect 564532 33730 564584 33736
rect 564440 3528 564492 3534
rect 564440 3470 564492 3476
rect 564544 3346 564572 33730
rect 565832 16574 565860 35226
rect 566464 28280 566516 28286
rect 566464 28222 566516 28228
rect 565832 16546 566412 16574
rect 565268 3528 565320 3534
rect 565268 3470 565320 3476
rect 566384 3482 566412 16546
rect 566476 4146 566504 28222
rect 569972 16574 570000 43386
rect 571340 18692 571392 18698
rect 571340 18634 571392 18640
rect 569972 16546 570368 16574
rect 569132 6316 569184 6322
rect 569132 6258 569184 6264
rect 566464 4140 566516 4146
rect 566464 4082 566516 4088
rect 568028 4140 568080 4146
rect 568028 4082 568080 4088
rect 564452 3318 564572 3346
rect 564452 480 564480 3318
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565280 354 565308 3470
rect 566384 3454 566872 3482
rect 566844 480 566872 3454
rect 568040 480 568068 4082
rect 569144 480 569172 6258
rect 570340 480 570368 16546
rect 565606 354 565718 480
rect 565280 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571352 354 571380 18634
rect 572732 16574 572760 54470
rect 578240 26920 578292 26926
rect 578240 26862 578292 26868
rect 576124 22908 576176 22914
rect 576124 22850 576176 22856
rect 574100 18624 574152 18630
rect 574100 18566 574152 18572
rect 574112 16574 574140 18566
rect 572732 16546 573496 16574
rect 574112 16546 575152 16574
rect 572720 6248 572772 6254
rect 572720 6190 572772 6196
rect 572732 480 572760 6190
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573468 354 573496 16546
rect 575124 480 575152 16546
rect 576136 4146 576164 22850
rect 578252 16574 578280 26862
rect 578252 16546 578648 16574
rect 576308 6180 576360 6186
rect 576308 6122 576360 6128
rect 576124 4140 576176 4146
rect 576124 4082 576176 4088
rect 576320 480 576348 6122
rect 577412 4140 577464 4146
rect 577412 4082 577464 4088
rect 577424 480 577452 4082
rect 578620 480 578648 16546
rect 581000 3596 581052 3602
rect 581000 3538 581052 3544
rect 581012 480 581040 3538
rect 582196 3460 582248 3466
rect 582196 3402 582248 3408
rect 582208 480 582236 3402
rect 583390 3360 583446 3369
rect 583390 3295 583446 3304
rect 583404 480 583432 3295
rect 573886 354 573998 480
rect 573468 326 573998 354
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 57610 445440 57666 445496
rect 57610 59880 57666 59936
rect 57978 59744 58034 59800
rect 61014 59744 61070 59800
rect 64326 59764 64382 59800
rect 64326 59744 64328 59764
rect 64328 59744 64380 59764
rect 64380 59744 64382 59764
rect 70214 59744 70270 59800
rect 60462 59628 60518 59664
rect 60462 59608 60464 59628
rect 60464 59608 60516 59628
rect 60516 59608 60518 59628
rect 62670 59608 62726 59664
rect 61382 59472 61438 59528
rect 59358 59336 59414 59392
rect 19430 3304 19486 3360
rect 62670 59336 62726 59392
rect 69294 59628 69350 59664
rect 69294 59608 69296 59628
rect 69296 59608 69348 59628
rect 69348 59608 69350 59628
rect 70122 59608 70178 59664
rect 64510 59472 64566 59528
rect 66810 59472 66866 59528
rect 63406 59336 63462 59392
rect 64694 59336 64750 59392
rect 66166 59336 66222 59392
rect 66810 59200 66866 59256
rect 67270 59200 67326 59256
rect 68834 59472 68890 59528
rect 68650 59336 68706 59392
rect 75090 59764 75146 59800
rect 75090 59744 75092 59764
rect 75092 59744 75144 59764
rect 75144 59744 75146 59764
rect 79966 59764 80022 59800
rect 79966 59744 79968 59764
rect 79968 59744 80020 59764
rect 80020 59744 80022 59764
rect 84198 59744 84254 59800
rect 70214 59472 70270 59528
rect 70122 59336 70178 59392
rect 70306 59336 70362 59392
rect 71410 59200 71466 59256
rect 71594 59064 71650 59120
rect 76654 59608 76710 59664
rect 77482 59628 77538 59664
rect 77482 59608 77484 59628
rect 77484 59608 77536 59628
rect 77536 59608 77538 59628
rect 74446 59336 74502 59392
rect 72974 58928 73030 58984
rect 75182 59200 75238 59256
rect 76562 59472 76618 59528
rect 76654 59336 76710 59392
rect 76838 59336 76894 59392
rect 79322 59608 79378 59664
rect 81622 59608 81678 59664
rect 83278 59608 83334 59664
rect 80702 59472 80758 59528
rect 79506 59336 79562 59392
rect 81622 59336 81678 59392
rect 84106 59608 84162 59664
rect 83646 59336 83702 59392
rect 93858 59764 93914 59800
rect 93858 59744 93860 59764
rect 93860 59744 93912 59764
rect 93912 59744 93914 59764
rect 97354 59744 97410 59800
rect 85762 59608 85818 59664
rect 84842 59472 84898 59528
rect 89074 59628 89130 59664
rect 89074 59608 89076 59628
rect 89076 59608 89128 59628
rect 89128 59608 89130 59628
rect 89902 59608 89958 59664
rect 87418 59492 87474 59528
rect 87418 59472 87420 59492
rect 87420 59472 87472 59492
rect 87472 59472 87474 59492
rect 85762 59336 85818 59392
rect 86222 59336 86278 59392
rect 86222 3304 86278 3360
rect 89626 59472 89682 59528
rect 87786 59200 87842 59256
rect 91558 59492 91614 59528
rect 91558 59472 91560 59492
rect 91560 59472 91612 59492
rect 91612 59472 91614 59492
rect 89902 59336 89958 59392
rect 90730 59336 90786 59392
rect 90914 59200 90970 59256
rect 101402 59764 101458 59800
rect 105634 59780 105636 59800
rect 105636 59780 105688 59800
rect 105688 59780 105690 59800
rect 101402 59744 101404 59764
rect 101404 59744 101456 59764
rect 101456 59744 101458 59764
rect 105634 59744 105690 59780
rect 107198 59744 107254 59800
rect 108026 59764 108082 59800
rect 108026 59744 108028 59764
rect 108028 59744 108080 59764
rect 108080 59744 108082 59764
rect 95422 59608 95478 59664
rect 93766 59472 93822 59528
rect 93674 59336 93730 59392
rect 95422 59336 95478 59392
rect 95146 59200 95202 59256
rect 93858 59064 93914 59120
rect 97446 59608 97502 59664
rect 97354 59336 97410 59392
rect 99746 59608 99802 59664
rect 98826 59472 98882 59528
rect 99746 59336 99802 59392
rect 100022 59336 100078 59392
rect 101586 59472 101642 59528
rect 101586 59336 101642 59392
rect 103978 59608 104034 59664
rect 103150 59472 103206 59528
rect 103978 59336 104034 59392
rect 104162 59200 104218 59256
rect 107106 59608 107162 59664
rect 105726 59472 105782 59528
rect 106922 59336 106978 59392
rect 108854 59744 108910 59800
rect 111338 59780 111340 59800
rect 111340 59780 111392 59800
rect 111392 59780 111394 59800
rect 107198 59472 107254 59528
rect 108302 59472 108358 59528
rect 108854 59336 108910 59392
rect 109682 59336 109738 59392
rect 111338 59744 111394 59780
rect 113730 59764 113786 59800
rect 113730 59744 113732 59764
rect 113732 59744 113784 59764
rect 113784 59744 113786 59764
rect 116214 59764 116270 59800
rect 116214 59744 116216 59764
rect 116216 59744 116268 59764
rect 116268 59744 116270 59764
rect 122010 59764 122066 59800
rect 122010 59744 122012 59764
rect 122012 59744 122064 59764
rect 122064 59744 122066 59764
rect 123114 59744 123170 59800
rect 111338 59608 111394 59664
rect 111246 59472 111302 59528
rect 113822 59472 113878 59528
rect 111338 59336 111394 59392
rect 112442 59336 112498 59392
rect 114190 59608 114246 59664
rect 117226 59472 117282 59528
rect 114190 59336 114246 59392
rect 115386 59336 115442 59392
rect 115846 59200 115902 59256
rect 117870 59608 117926 59664
rect 117778 59336 117834 59392
rect 117962 59336 118018 59392
rect 119342 59200 119398 59256
rect 120354 59628 120410 59664
rect 120354 59608 120356 59628
rect 120356 59608 120408 59628
rect 120408 59608 120410 59628
rect 122286 59608 122342 59664
rect 122102 59472 122158 59528
rect 120722 59336 120778 59392
rect 126426 59764 126482 59800
rect 126426 59744 126428 59764
rect 126428 59744 126480 59764
rect 126480 59744 126482 59764
rect 130198 59764 130254 59800
rect 130198 59744 130200 59764
rect 130200 59744 130252 59764
rect 130252 59744 130254 59764
rect 123298 59608 123354 59664
rect 123114 59336 123170 59392
rect 123666 59336 123722 59392
rect 123666 59200 123722 59256
rect 126242 59608 126298 59664
rect 126426 59608 126482 59664
rect 126242 59336 126298 59392
rect 128542 59608 128598 59664
rect 127806 59472 127862 59528
rect 130382 59472 130438 59528
rect 128542 59336 128598 59392
rect 129002 59336 129058 59392
rect 131026 59744 131082 59800
rect 132038 59744 132094 59800
rect 133142 59744 133198 59800
rect 133510 59744 133566 59800
rect 134338 59744 134394 59800
rect 135258 59744 135314 59800
rect 131946 59628 132002 59664
rect 131946 59608 131948 59628
rect 131948 59608 132000 59628
rect 132000 59608 132002 59628
rect 130658 59336 130714 59392
rect 131118 59336 131174 59392
rect 133142 59472 133198 59528
rect 134338 59336 134394 59392
rect 135166 59608 135222 59664
rect 141698 59764 141754 59800
rect 141698 59744 141700 59764
rect 141700 59744 141752 59764
rect 141752 59744 141754 59764
rect 136822 59608 136878 59664
rect 135258 59472 135314 59528
rect 135902 59472 135958 59528
rect 134706 59200 134762 59256
rect 139306 59472 139362 59528
rect 136822 59336 136878 59392
rect 137374 59336 137430 59392
rect 138110 59372 138112 59392
rect 138112 59372 138164 59392
rect 138164 59372 138166 59392
rect 138110 59336 138166 59372
rect 136086 59200 136142 59256
rect 138662 59200 138718 59256
rect 138846 59064 138902 59120
rect 141698 59628 141754 59664
rect 141698 59608 141700 59628
rect 141700 59608 141752 59628
rect 141752 59608 141754 59628
rect 141514 59472 141570 59528
rect 144458 59744 144514 59800
rect 145838 59744 145894 59800
rect 148690 59744 148746 59800
rect 144550 59608 144606 59664
rect 142894 59336 142950 59392
rect 144182 59336 144238 59392
rect 142066 59200 142122 59256
rect 144734 59472 144790 59528
rect 145838 59472 145894 59528
rect 146206 59336 146262 59392
rect 151910 59764 151966 59800
rect 151910 59744 151912 59764
rect 151912 59744 151964 59764
rect 151964 59744 151966 59764
rect 158166 59764 158222 59800
rect 158166 59744 158168 59764
rect 158168 59744 158220 59764
rect 158220 59744 158222 59764
rect 164054 59744 164110 59800
rect 149978 59472 150034 59528
rect 148874 59200 148930 59256
rect 144826 3304 144882 3360
rect 151634 59628 151690 59664
rect 151634 59608 151636 59628
rect 151636 59608 151688 59628
rect 151688 59608 151690 59628
rect 152830 59608 152886 59664
rect 154946 59608 155002 59664
rect 151726 59472 151782 59528
rect 154302 59472 154358 59528
rect 153014 59336 153070 59392
rect 156970 59472 157026 59528
rect 154946 59336 155002 59392
rect 155866 59336 155922 59392
rect 157246 59608 157302 59664
rect 157614 59608 157670 59664
rect 162766 59608 162822 59664
rect 158350 59472 158406 59528
rect 161202 59472 161258 59528
rect 157614 59336 157670 59392
rect 158626 59336 158682 59392
rect 162490 59336 162546 59392
rect 162674 59200 162730 59256
rect 173346 59764 173402 59800
rect 173346 59744 173348 59764
rect 173348 59744 173400 59764
rect 173400 59744 173402 59764
rect 183742 59764 183798 59800
rect 183742 59744 183744 59764
rect 183744 59744 183796 59764
rect 183796 59744 183798 59764
rect 185398 59744 185454 59800
rect 186226 59744 186282 59800
rect 164790 59608 164846 59664
rect 164146 59472 164202 59528
rect 166446 59628 166502 59664
rect 166446 59608 166448 59628
rect 166448 59608 166500 59628
rect 166500 59608 166502 59628
rect 167274 59608 167330 59664
rect 164790 59336 164846 59392
rect 165250 59336 165306 59392
rect 166814 59472 166870 59528
rect 168930 59492 168986 59528
rect 168930 59472 168932 59492
rect 168932 59472 168984 59492
rect 168984 59472 168986 59492
rect 171414 59492 171470 59528
rect 171414 59472 171416 59492
rect 171416 59472 171468 59492
rect 171468 59472 171470 59492
rect 167274 59336 167330 59392
rect 168286 59336 168342 59392
rect 170770 59336 170826 59392
rect 169574 59200 169630 59256
rect 170954 59064 171010 59120
rect 173530 59608 173586 59664
rect 175462 59608 175518 59664
rect 177118 59628 177174 59664
rect 177118 59608 177120 59628
rect 177120 59608 177172 59628
rect 177172 59608 177174 59628
rect 173714 59336 173770 59392
rect 175094 59472 175150 59528
rect 177946 59608 178002 59664
rect 177670 59472 177726 59528
rect 175462 59336 175518 59392
rect 176566 59336 176622 59392
rect 180430 59492 180486 59528
rect 180430 59472 180432 59492
rect 180432 59472 180484 59492
rect 180484 59472 180486 59492
rect 177946 59336 178002 59392
rect 177854 59200 177910 59256
rect 179142 59200 179198 59256
rect 180706 59336 180762 59392
rect 181074 59336 181130 59392
rect 180798 59200 180854 59256
rect 181994 59064 182050 59120
rect 184846 59472 184902 59528
rect 183190 59200 183246 59256
rect 183374 59064 183430 59120
rect 185950 59608 186006 59664
rect 185398 59336 185454 59392
rect 194414 59764 194470 59800
rect 194414 59744 194416 59764
rect 194416 59744 194468 59764
rect 194468 59744 194470 59764
rect 195242 59744 195298 59800
rect 187882 59608 187938 59664
rect 186226 59472 186282 59528
rect 187330 59472 187386 59528
rect 186134 59336 186190 59392
rect 190274 59492 190330 59528
rect 190274 59472 190276 59492
rect 190276 59472 190328 59492
rect 190328 59472 190330 59492
rect 187882 59336 187938 59392
rect 187514 59200 187570 59256
rect 190550 59336 190606 59392
rect 190366 59200 190422 59256
rect 191746 59064 191802 59120
rect 194506 59608 194562 59664
rect 194414 59472 194470 59528
rect 193034 59200 193090 59256
rect 202786 59764 202842 59800
rect 202786 59744 202788 59764
rect 202788 59744 202840 59764
rect 202840 59744 202842 59764
rect 209410 59764 209466 59800
rect 209410 59744 209412 59764
rect 209412 59744 209464 59764
rect 209464 59744 209466 59764
rect 211710 59744 211766 59800
rect 195794 59608 195850 59664
rect 195242 59336 195298 59392
rect 195610 59336 195666 59392
rect 197082 59608 197138 59664
rect 197082 59472 197138 59528
rect 196990 59336 197046 59392
rect 197266 59336 197322 59392
rect 198646 59200 198702 59256
rect 201038 59608 201094 59664
rect 200026 59472 200082 59528
rect 200210 59472 200266 59528
rect 201038 59336 201094 59392
rect 201222 59336 201278 59392
rect 204166 59608 204222 59664
rect 206098 59608 206154 59664
rect 202786 59472 202842 59528
rect 203982 59336 204038 59392
rect 205454 59472 205510 59528
rect 207570 59492 207626 59528
rect 207570 59472 207572 59492
rect 207572 59472 207624 59492
rect 207624 59472 207626 59492
rect 206098 59336 206154 59392
rect 206926 59336 206982 59392
rect 208030 59200 208086 59256
rect 211066 59608 211122 59664
rect 209410 59472 209466 59528
rect 209594 59200 209650 59256
rect 215850 59764 215906 59800
rect 215850 59744 215852 59764
rect 215852 59744 215904 59764
rect 215904 59744 215906 59764
rect 223210 59744 223266 59800
rect 212354 59472 212410 59528
rect 211710 59336 211766 59392
rect 212170 59336 212226 59392
rect 219162 59628 219218 59664
rect 219162 59608 219164 59628
rect 219164 59608 219216 59628
rect 219216 59608 219218 59628
rect 219990 59608 220046 59664
rect 216494 59472 216550 59528
rect 215206 59336 215262 59392
rect 216310 59336 216366 59392
rect 213734 59200 213790 59256
rect 219346 59472 219402 59528
rect 217874 59200 217930 59256
rect 222014 59472 222070 59528
rect 219990 59336 220046 59392
rect 221922 59336 221978 59392
rect 220450 59200 220506 59256
rect 220634 59064 220690 59120
rect 224866 59472 224922 59528
rect 223210 59336 223266 59392
rect 223486 59336 223542 59392
rect 224774 59336 224830 59392
rect 226522 59472 226578 59528
rect 225970 59336 226026 59392
rect 226154 59336 226210 59392
rect 225970 59200 226026 59256
rect 229006 59744 229062 59800
rect 229466 59780 229468 59800
rect 229468 59780 229520 59800
rect 229520 59780 229522 59800
rect 229466 59744 229522 59780
rect 230662 59780 230664 59800
rect 230664 59780 230716 59800
rect 230716 59780 230718 59800
rect 230662 59744 230718 59780
rect 234802 59764 234858 59800
rect 234802 59744 234804 59764
rect 234804 59744 234856 59764
rect 234856 59744 234858 59764
rect 235630 59744 235686 59800
rect 229006 59628 229062 59664
rect 229006 59608 229008 59628
rect 229008 59608 229060 59628
rect 229060 59608 229062 59628
rect 229006 59472 229062 59528
rect 229926 59336 229982 59392
rect 229742 59200 229798 59256
rect 231122 59064 231178 59120
rect 232686 59608 232742 59664
rect 234802 59608 234858 59664
rect 234066 59472 234122 59528
rect 233882 59336 233938 59392
rect 238850 59744 238906 59800
rect 240506 59780 240508 59800
rect 240508 59780 240560 59800
rect 240560 59780 240562 59800
rect 235630 59472 235686 59528
rect 234802 59336 234858 59392
rect 235446 59336 235502 59392
rect 235262 59200 235318 59256
rect 240506 59744 240562 59780
rect 242162 59764 242218 59800
rect 242162 59744 242164 59764
rect 242164 59744 242216 59764
rect 242216 59744 242218 59764
rect 245474 59764 245530 59800
rect 245474 59744 245476 59764
rect 245476 59744 245528 59764
rect 245528 59744 245530 59764
rect 250534 59744 250590 59800
rect 251270 59764 251326 59800
rect 251270 59744 251272 59764
rect 251272 59744 251324 59764
rect 251324 59744 251326 59764
rect 238298 59472 238354 59528
rect 242346 59472 242402 59528
rect 239586 59336 239642 59392
rect 240782 59200 240838 59256
rect 242162 59064 242218 59120
rect 243542 59200 243598 59256
rect 245474 59608 245530 59664
rect 244922 59472 244978 59528
rect 248878 59628 248934 59664
rect 248878 59608 248880 59628
rect 248880 59608 248932 59628
rect 248932 59608 248934 59628
rect 245474 59336 245530 59392
rect 247682 59336 247738 59392
rect 247958 59492 248014 59528
rect 247958 59472 247960 59492
rect 247960 59472 248012 59492
rect 248012 59472 248014 59492
rect 249614 59608 249670 59664
rect 250626 59608 250682 59664
rect 250442 59472 250498 59528
rect 249614 59336 249670 59392
rect 252282 59744 252338 59800
rect 254582 59744 254638 59800
rect 267462 59764 267518 59800
rect 267462 59744 267464 59764
rect 267464 59744 267516 59764
rect 267516 59744 267518 59764
rect 252006 59472 252062 59528
rect 252282 59472 252338 59528
rect 269854 59744 269910 59800
rect 270682 59764 270738 59800
rect 270682 59744 270684 59764
rect 270684 59744 270736 59764
rect 270736 59744 270738 59764
rect 278042 59744 278098 59800
rect 278870 59744 278926 59800
rect 281354 59744 281410 59800
rect 257802 59628 257858 59664
rect 257802 59608 257804 59628
rect 257804 59608 257856 59628
rect 257856 59608 257858 59628
rect 258630 59608 258686 59664
rect 255134 59472 255190 59528
rect 254582 59336 254638 59392
rect 254950 59336 255006 59392
rect 252466 59200 252522 59256
rect 253846 59200 253902 59256
rect 257986 59472 258042 59528
rect 256514 59200 256570 59256
rect 261114 59628 261170 59664
rect 261114 59608 261116 59628
rect 261116 59608 261168 59628
rect 261168 59608 261170 59628
rect 265714 59608 265770 59664
rect 258630 59336 258686 59392
rect 260746 59472 260802 59528
rect 259274 59200 259330 59256
rect 267002 59472 267058 59528
rect 269762 59472 269818 59528
rect 265530 59336 265586 59392
rect 265714 59336 265770 59392
rect 268566 59336 268622 59392
rect 268382 59200 268438 59256
rect 270682 59608 270738 59664
rect 272246 59492 272302 59528
rect 272246 59472 272248 59492
rect 272248 59472 272300 59492
rect 272300 59472 272302 59492
rect 276386 59608 276442 59664
rect 273902 59492 273958 59528
rect 273902 59472 273904 59492
rect 273904 59472 273956 59492
rect 273956 59472 273958 59492
rect 277214 59472 277270 59528
rect 276386 59336 276442 59392
rect 273718 59200 273774 59256
rect 274638 59200 274694 59256
rect 276846 59200 276902 59256
rect 279422 59608 279478 59664
rect 280342 59628 280398 59664
rect 280342 59608 280344 59628
rect 280344 59608 280396 59628
rect 280396 59608 280398 59628
rect 278042 59472 278098 59528
rect 278870 59472 278926 59528
rect 277950 59336 278006 59392
rect 283010 59764 283066 59800
rect 283010 59744 283012 59764
rect 283012 59744 283064 59764
rect 283064 59744 283066 59764
rect 286322 59744 286378 59800
rect 287150 59744 287206 59800
rect 287886 59764 287942 59800
rect 287886 59744 287888 59764
rect 287888 59744 287940 59764
rect 287940 59744 287942 59764
rect 280802 59472 280858 59528
rect 281722 59472 281778 59528
rect 280986 59336 281042 59392
rect 283010 59472 283066 59528
rect 282366 59200 282422 59256
rect 286322 59472 286378 59528
rect 284942 59200 284998 59256
rect 291750 59744 291806 59800
rect 293406 59744 293462 59800
rect 293682 59764 293738 59800
rect 293682 59744 293684 59764
rect 293684 59744 293736 59764
rect 293736 59744 293738 59764
rect 287702 59608 287758 59664
rect 287150 59336 287206 59392
rect 286506 59200 286562 59256
rect 289542 59608 289598 59664
rect 290462 59472 290518 59528
rect 289082 59336 289138 59392
rect 289542 59336 289598 59392
rect 292026 59608 292082 59664
rect 291842 59336 291898 59392
rect 294418 59744 294474 59800
rect 296994 59780 296996 59800
rect 296996 59780 297048 59800
rect 297048 59780 297050 59800
rect 296994 59744 297050 59780
rect 294418 59336 294474 59392
rect 294510 58928 294566 58984
rect 296534 59608 296590 59664
rect 296994 59472 297050 59528
rect 296166 59336 296222 59392
rect 300306 59744 300362 59800
rect 301134 59744 301190 59800
rect 301962 59764 302018 59800
rect 301962 59744 301964 59764
rect 301964 59744 302016 59764
rect 302016 59744 302018 59764
rect 300122 59472 300178 59528
rect 305918 59744 305974 59800
rect 312634 59744 312690 59800
rect 314290 59764 314346 59800
rect 314290 59744 314292 59764
rect 314292 59744 314344 59764
rect 314344 59744 314346 59764
rect 301502 59608 301558 59664
rect 300306 59336 300362 59392
rect 301134 59336 301190 59392
rect 303066 59200 303122 59256
rect 304354 59608 304410 59664
rect 305642 59472 305698 59528
rect 304354 59336 304410 59392
rect 304446 59200 304502 59256
rect 306010 59628 306066 59664
rect 306010 59608 306012 59628
rect 306012 59608 306064 59628
rect 306064 59608 306066 59628
rect 310150 59628 310206 59664
rect 310150 59608 310152 59628
rect 310152 59608 310204 59628
rect 310204 59608 310206 59628
rect 312542 59644 312544 59664
rect 312544 59644 312596 59664
rect 312596 59644 312598 59664
rect 312542 59608 312598 59644
rect 306838 59356 306894 59392
rect 306838 59336 306840 59356
rect 306840 59336 306892 59356
rect 306892 59336 306894 59356
rect 307022 59200 307078 59256
rect 305918 59064 305974 59120
rect 308494 59492 308550 59528
rect 308494 59472 308496 59492
rect 308496 59472 308548 59492
rect 308548 59472 308550 59492
rect 312542 59472 312598 59528
rect 309782 59200 309838 59256
rect 308586 59064 308642 59120
rect 311346 59336 311402 59392
rect 316774 59744 316830 59800
rect 316958 59744 317014 59800
rect 320822 59764 320878 59800
rect 320822 59744 320824 59764
rect 320824 59744 320876 59764
rect 320876 59744 320878 59764
rect 312634 59336 312690 59392
rect 314290 59472 314346 59528
rect 315302 59200 315358 59256
rect 316774 59336 316830 59392
rect 324134 59744 324190 59800
rect 324962 59764 325018 59800
rect 324962 59744 324964 59764
rect 324964 59744 325016 59764
rect 325016 59744 325018 59764
rect 317418 59608 317474 59664
rect 322478 59608 322534 59664
rect 316866 59200 316922 59256
rect 320362 59472 320418 59528
rect 318890 59200 318946 59256
rect 320546 59336 320602 59392
rect 321650 59336 321706 59392
rect 322478 59336 322534 59392
rect 323306 59472 323362 59528
rect 330298 59744 330354 59800
rect 334898 59764 334954 59800
rect 334898 59744 334900 59764
rect 334900 59744 334952 59764
rect 334952 59744 334954 59764
rect 324778 59608 324834 59664
rect 324134 59336 324190 59392
rect 324594 59200 324650 59256
rect 325790 59356 325846 59392
rect 325790 59336 325792 59356
rect 325792 59336 325844 59356
rect 325844 59336 325846 59356
rect 325698 59200 325754 59256
rect 329102 59492 329158 59528
rect 329102 59472 329104 59492
rect 329104 59472 329156 59492
rect 329156 59472 329158 59492
rect 329930 59336 329986 59392
rect 328826 59200 328882 59256
rect 328642 59064 328698 59120
rect 339038 59764 339094 59800
rect 339038 59744 339040 59764
rect 339040 59744 339092 59764
rect 339092 59744 339094 59764
rect 341522 59764 341578 59800
rect 341522 59744 341524 59764
rect 341524 59744 341576 59764
rect 341576 59744 341578 59764
rect 343086 59764 343142 59800
rect 343086 59744 343088 59764
rect 343088 59744 343140 59764
rect 343140 59744 343142 59764
rect 347962 59744 348018 59800
rect 348422 59744 348478 59800
rect 355230 59744 355286 59800
rect 359554 59764 359610 59800
rect 359554 59744 359556 59764
rect 359556 59744 359608 59764
rect 359608 59744 359610 59764
rect 333242 59608 333298 59664
rect 331494 59472 331550 59528
rect 334070 59472 334126 59528
rect 332690 59336 332746 59392
rect 333242 59336 333298 59392
rect 335358 59336 335414 59392
rect 335542 59200 335598 59256
rect 335450 59064 335506 59120
rect 338118 59472 338174 59528
rect 340970 59472 341026 59528
rect 338210 59336 338266 59392
rect 339590 59336 339646 59392
rect 342350 59336 342406 59392
rect 343638 59472 343694 59528
rect 344742 59492 344798 59528
rect 344742 59472 344744 59492
rect 344744 59472 344796 59492
rect 344796 59472 344798 59492
rect 348054 59608 348110 59664
rect 347962 59472 348018 59528
rect 345294 59336 345350 59392
rect 346398 59200 346454 59256
rect 347870 59336 347926 59392
rect 348054 59336 348110 59392
rect 349250 59472 349306 59528
rect 351366 59492 351422 59528
rect 351366 59472 351368 59492
rect 351368 59472 351420 59492
rect 351420 59472 351422 59492
rect 349434 59336 349490 59392
rect 350538 59200 350594 59256
rect 351918 59200 351974 59256
rect 353390 59200 353446 59256
rect 354586 59336 354642 59392
rect 354954 59472 355010 59528
rect 363694 59764 363750 59800
rect 363694 59744 363696 59764
rect 363696 59744 363748 59764
rect 363748 59744 363750 59764
rect 365166 59744 365222 59800
rect 357070 59608 357126 59664
rect 358910 59608 358966 59664
rect 356058 59472 356114 59528
rect 355230 59336 355286 59392
rect 357622 59472 357678 59528
rect 357070 59336 357126 59392
rect 358818 59336 358874 59392
rect 357806 59200 357862 59256
rect 360198 59336 360254 59392
rect 361578 59200 361634 59256
rect 367006 59764 367062 59800
rect 367006 59744 367008 59764
rect 367008 59744 367060 59764
rect 367060 59744 367062 59764
rect 369398 59764 369454 59800
rect 369398 59744 369400 59764
rect 369400 59744 369452 59764
rect 369452 59744 369454 59764
rect 371054 59764 371110 59800
rect 371054 59744 371056 59764
rect 371056 59744 371108 59764
rect 371108 59744 371110 59764
rect 376022 59764 376078 59800
rect 380070 59780 380072 59800
rect 380072 59780 380124 59800
rect 380124 59780 380126 59800
rect 376022 59744 376024 59764
rect 376024 59744 376076 59764
rect 376076 59744 376078 59764
rect 380070 59744 380126 59780
rect 380990 59764 381046 59800
rect 380990 59744 380992 59764
rect 380992 59744 381044 59764
rect 381044 59744 381046 59764
rect 364982 59608 365038 59664
rect 363786 59472 363842 59528
rect 363602 59336 363658 59392
rect 367742 59200 367798 59256
rect 367742 59064 367798 59120
rect 371054 59608 371110 59664
rect 369950 59472 370006 59528
rect 370686 59472 370742 59528
rect 369950 59336 370006 59392
rect 370502 59336 370558 59392
rect 376022 59628 376078 59664
rect 376022 59608 376024 59628
rect 376024 59608 376076 59628
rect 376076 59608 376078 59628
rect 378506 59608 378562 59664
rect 372710 59492 372766 59528
rect 372710 59472 372712 59492
rect 372712 59472 372764 59492
rect 372764 59472 372766 59492
rect 376022 59472 376078 59528
rect 374642 59200 374698 59256
rect 376206 59200 376262 59256
rect 378506 59336 378562 59392
rect 378782 59200 378838 59256
rect 379426 59472 379482 59528
rect 380990 59608 381046 59664
rect 380806 59336 380862 59392
rect 387522 59764 387578 59800
rect 387522 59744 387524 59764
rect 387524 59744 387576 59764
rect 387576 59744 387578 59764
rect 390006 59744 390062 59800
rect 390834 59744 390890 59800
rect 391662 59764 391718 59800
rect 391662 59744 391664 59764
rect 391664 59744 391716 59764
rect 391716 59744 391718 59764
rect 383198 59608 383254 59664
rect 385866 59608 385922 59664
rect 383474 59472 383530 59528
rect 383198 59336 383254 59392
rect 387246 59472 387302 59528
rect 384118 59356 384174 59392
rect 384118 59336 384120 59356
rect 384120 59336 384172 59356
rect 384172 59336 384174 59356
rect 385866 59336 385922 59392
rect 384302 59200 384358 59256
rect 387062 59200 387118 59256
rect 388626 59336 388682 59392
rect 388442 59200 388498 59256
rect 390006 59472 390062 59528
rect 397458 59764 397514 59800
rect 397458 59744 397460 59764
rect 397460 59744 397512 59764
rect 397512 59744 397514 59764
rect 402334 59764 402390 59800
rect 402334 59744 402336 59764
rect 402336 59744 402388 59764
rect 402388 59744 402390 59764
rect 406474 59764 406530 59800
rect 406474 59744 406476 59764
rect 406476 59744 406528 59764
rect 406528 59744 406530 59764
rect 410614 59764 410670 59800
rect 410614 59744 410616 59764
rect 410616 59744 410668 59764
rect 410668 59744 410670 59764
rect 416870 59744 416926 59800
rect 419538 59744 419594 59800
rect 425518 59764 425574 59800
rect 425518 59744 425520 59764
rect 425520 59744 425572 59764
rect 425572 59744 425574 59764
rect 391202 59608 391258 59664
rect 390834 59336 390890 59392
rect 393318 59628 393374 59664
rect 393318 59608 393320 59628
rect 393320 59608 393372 59628
rect 393372 59608 393374 59628
rect 393318 59472 393374 59528
rect 393686 59472 393742 59528
rect 392766 59336 392822 59392
rect 395802 59608 395858 59664
rect 397458 59608 397514 59664
rect 397826 59608 397882 59664
rect 398286 59608 398342 59664
rect 394146 59472 394202 59528
rect 396722 59472 396778 59528
rect 398102 59492 398158 59528
rect 398102 59472 398104 59492
rect 398104 59472 398156 59492
rect 398156 59472 398158 59492
rect 395802 59336 395858 59392
rect 398010 59336 398066 59392
rect 396906 59200 396962 59256
rect 399942 59608 399998 59664
rect 400770 59608 400826 59664
rect 400862 59472 400918 59528
rect 399942 59336 399998 59392
rect 400770 59336 400826 59392
rect 401598 59336 401654 59392
rect 403070 59336 403126 59392
rect 402242 59200 402298 59256
rect 404358 59200 404414 59256
rect 405922 59472 405978 59528
rect 408130 59492 408186 59528
rect 408130 59472 408132 59492
rect 408132 59472 408184 59492
rect 408184 59472 408186 59492
rect 406106 59336 406162 59392
rect 407302 59200 407358 59256
rect 412086 59608 412142 59664
rect 409970 59472 410026 59528
rect 408682 59336 408738 59392
rect 412730 59472 412786 59528
rect 411350 59336 411406 59392
rect 412086 59336 412142 59392
rect 413098 59628 413154 59664
rect 413098 59608 413100 59628
rect 413100 59608 413152 59628
rect 413152 59608 413154 59628
rect 416410 59628 416466 59664
rect 416410 59608 416412 59628
rect 416412 59608 416464 59628
rect 416464 59608 416466 59628
rect 412914 59472 412970 59528
rect 413926 59336 413982 59392
rect 416778 59472 416834 59528
rect 416962 59336 417018 59392
rect 418158 59336 418214 59392
rect 427082 59764 427138 59800
rect 427082 59744 427084 59764
rect 427084 59744 427136 59764
rect 427136 59744 427138 59764
rect 431222 59764 431278 59800
rect 431222 59744 431224 59764
rect 431224 59744 431276 59764
rect 431276 59744 431278 59764
rect 435454 59744 435510 59800
rect 420918 59608 420974 59664
rect 425334 59472 425390 59528
rect 422390 59336 422446 59392
rect 425150 59336 425206 59392
rect 421102 59200 421158 59256
rect 423770 59200 423826 59256
rect 426438 59200 426494 59256
rect 428738 59492 428794 59528
rect 428738 59472 428740 59492
rect 428740 59472 428792 59492
rect 428792 59472 428794 59492
rect 429382 59336 429438 59392
rect 427910 59200 427966 59256
rect 430578 59472 430634 59528
rect 432050 59492 432106 59528
rect 432050 59472 432052 59492
rect 432052 59472 432104 59492
rect 432104 59472 432106 59492
rect 432050 59336 432106 59392
rect 436926 59764 436982 59800
rect 436926 59744 436928 59764
rect 436928 59744 436980 59764
rect 436980 59744 436982 59764
rect 440238 59744 440294 59800
rect 441158 59744 441214 59800
rect 441434 59744 441490 59800
rect 441894 59764 441950 59800
rect 441894 59744 441896 59764
rect 441896 59744 441948 59764
rect 441948 59744 441950 59764
rect 438582 59608 438638 59664
rect 434718 59472 434774 59528
rect 435638 59472 435694 59528
rect 436374 59472 436430 59528
rect 434902 59336 434958 59392
rect 436190 59200 436246 59256
rect 439042 59472 439098 59528
rect 437478 59336 437534 59392
rect 438582 59336 438638 59392
rect 445942 59744 445998 59800
rect 446862 59764 446918 59800
rect 446862 59744 446864 59764
rect 446864 59744 446916 59764
rect 446916 59744 446918 59764
rect 440422 59608 440478 59664
rect 440238 59336 440294 59392
rect 440238 59200 440294 59256
rect 441710 59200 441766 59256
rect 445850 59608 445906 59664
rect 444378 59472 444434 59528
rect 443366 59200 443422 59256
rect 444470 59336 444526 59392
rect 449346 59744 449402 59800
rect 449714 59744 449770 59800
rect 457534 59764 457590 59800
rect 457534 59744 457536 59764
rect 457536 59744 457588 59764
rect 457588 59744 457590 59764
rect 446862 59608 446918 59664
rect 445942 59336 445998 59392
rect 448610 59472 448666 59528
rect 447414 59336 447470 59392
rect 449254 59628 449310 59664
rect 449254 59608 449256 59628
rect 449256 59608 449308 59628
rect 449308 59608 449310 59628
rect 449346 59336 449402 59392
rect 461582 59744 461638 59800
rect 464158 59764 464214 59800
rect 464158 59744 464160 59764
rect 464160 59744 464212 59764
rect 464212 59744 464214 59764
rect 453394 59628 453450 59664
rect 453394 59608 453396 59628
rect 453396 59608 453448 59628
rect 453448 59608 453450 59628
rect 455050 59492 455106 59528
rect 455050 59472 455052 59492
rect 455052 59472 455104 59492
rect 455104 59472 455106 59492
rect 455510 59336 455566 59392
rect 451278 59200 451334 59256
rect 452750 59200 452806 59256
rect 454038 59200 454094 59256
rect 452934 59064 452990 59120
rect 456798 59472 456854 59528
rect 459190 59492 459246 59528
rect 459190 59472 459192 59492
rect 459192 59472 459244 59492
rect 459244 59472 459246 59492
rect 458270 59200 458326 59256
rect 459742 59200 459798 59256
rect 461030 59200 461086 59256
rect 461674 59608 461730 59664
rect 461582 59336 461638 59392
rect 463974 59472 464030 59528
rect 463790 59336 463846 59392
rect 465078 59200 465134 59256
rect 467838 59472 467894 59528
rect 466550 59336 466606 59392
rect 583390 3304 583446 3360
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 57605 445498 57671 445501
rect 59494 445498 60076 445508
rect 57605 445496 60076 445498
rect 57605 445440 57610 445496
rect 57666 445448 60076 445496
rect 57666 445440 59554 445448
rect 57605 445438 59554 445440
rect 57605 445435 57671 445438
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 57605 59938 57671 59941
rect 60292 59938 60352 60044
rect 57605 59936 60352 59938
rect 57605 59880 57610 59936
rect 57666 59880 60352 59936
rect 57605 59878 60352 59880
rect 57605 59875 57671 59878
rect 57973 59802 58039 59805
rect 60844 59802 60904 60044
rect 57973 59800 60904 59802
rect 57973 59744 57978 59800
rect 58034 59744 60904 59800
rect 57973 59742 60904 59744
rect 61009 59802 61075 59805
rect 61672 59802 61732 60044
rect 61009 59800 61732 59802
rect 61009 59744 61014 59800
rect 61070 59744 61732 59800
rect 61009 59742 61732 59744
rect 57973 59739 58039 59742
rect 61009 59739 61075 59742
rect 60457 59666 60523 59669
rect 62500 59666 62560 60044
rect 60457 59664 62560 59666
rect 60457 59608 60462 59664
rect 60518 59608 62560 59664
rect 60457 59606 62560 59608
rect 62665 59666 62731 59669
rect 63328 59666 63388 60044
rect 62665 59664 63388 59666
rect 62665 59608 62670 59664
rect 62726 59608 63388 59664
rect 62665 59606 63388 59608
rect 60457 59603 60523 59606
rect 62665 59603 62731 59606
rect 61377 59530 61443 59533
rect 64156 59530 64216 60044
rect 64321 59802 64387 59805
rect 64984 59802 65044 60044
rect 64321 59800 65044 59802
rect 64321 59744 64326 59800
rect 64382 59744 65044 59800
rect 64321 59742 65044 59744
rect 64321 59739 64387 59742
rect 65812 59666 65872 60044
rect 61377 59528 64216 59530
rect 61377 59472 61382 59528
rect 61438 59472 64216 59528
rect 61377 59470 64216 59472
rect 64278 59606 65872 59666
rect 61377 59467 61443 59470
rect 59353 59394 59419 59397
rect 62665 59394 62731 59397
rect 59353 59392 62731 59394
rect 59353 59336 59358 59392
rect 59414 59336 62670 59392
rect 62726 59336 62731 59392
rect 59353 59334 62731 59336
rect 59353 59331 59419 59334
rect 62665 59331 62731 59334
rect 63401 59394 63467 59397
rect 64278 59394 64338 59606
rect 64505 59530 64571 59533
rect 66640 59530 66700 60044
rect 64505 59528 66700 59530
rect 64505 59472 64510 59528
rect 64566 59472 66700 59528
rect 64505 59470 66700 59472
rect 66805 59530 66871 59533
rect 67468 59530 67528 60044
rect 66805 59528 67528 59530
rect 66805 59472 66810 59528
rect 66866 59472 67528 59528
rect 66805 59470 67528 59472
rect 64505 59467 64571 59470
rect 66805 59467 66871 59470
rect 63401 59392 64338 59394
rect 63401 59336 63406 59392
rect 63462 59336 64338 59392
rect 63401 59334 64338 59336
rect 64689 59394 64755 59397
rect 66161 59394 66227 59397
rect 68296 59394 68356 60044
rect 69124 59666 69184 60044
rect 64689 59392 65994 59394
rect 64689 59336 64694 59392
rect 64750 59336 65994 59392
rect 64689 59334 65994 59336
rect 63401 59331 63467 59334
rect 64689 59331 64755 59334
rect 65934 59258 65994 59334
rect 66161 59392 68356 59394
rect 66161 59336 66166 59392
rect 66222 59336 68356 59392
rect 66161 59334 68356 59336
rect 68510 59606 69184 59666
rect 69289 59666 69355 59669
rect 69952 59666 70012 60044
rect 70209 59802 70275 59805
rect 70780 59802 70840 60044
rect 70209 59800 70840 59802
rect 70209 59744 70214 59800
rect 70270 59744 70840 59800
rect 70209 59742 70840 59744
rect 70209 59739 70275 59742
rect 69289 59664 70012 59666
rect 69289 59608 69294 59664
rect 69350 59608 70012 59664
rect 69289 59606 70012 59608
rect 70117 59666 70183 59669
rect 71608 59666 71668 60044
rect 70117 59664 71668 59666
rect 70117 59608 70122 59664
rect 70178 59608 71668 59664
rect 70117 59606 71668 59608
rect 66161 59331 66227 59334
rect 66805 59258 66871 59261
rect 65934 59256 66871 59258
rect 65934 59200 66810 59256
rect 66866 59200 66871 59256
rect 65934 59198 66871 59200
rect 66805 59195 66871 59198
rect 67265 59258 67331 59261
rect 68510 59258 68570 59606
rect 69289 59603 69355 59606
rect 70117 59603 70183 59606
rect 68829 59530 68895 59533
rect 70209 59530 70275 59533
rect 68829 59528 70275 59530
rect 68829 59472 68834 59528
rect 68890 59472 70214 59528
rect 70270 59472 70275 59528
rect 68829 59470 70275 59472
rect 68829 59467 68895 59470
rect 70209 59467 70275 59470
rect 68645 59394 68711 59397
rect 70117 59394 70183 59397
rect 68645 59392 70183 59394
rect 68645 59336 68650 59392
rect 68706 59336 70122 59392
rect 70178 59336 70183 59392
rect 68645 59334 70183 59336
rect 68645 59331 68711 59334
rect 70117 59331 70183 59334
rect 70301 59394 70367 59397
rect 72436 59394 72496 60044
rect 73264 59394 73324 60044
rect 74092 59394 74152 60044
rect 74920 59530 74980 60044
rect 75085 59802 75151 59805
rect 75748 59802 75808 60044
rect 75085 59800 75808 59802
rect 75085 59744 75090 59800
rect 75146 59744 75808 59800
rect 75085 59742 75808 59744
rect 75085 59739 75151 59742
rect 76484 59666 76544 60044
rect 70301 59392 72496 59394
rect 70301 59336 70306 59392
rect 70362 59336 72496 59392
rect 70301 59334 72496 59336
rect 72558 59334 73324 59394
rect 73478 59334 74152 59394
rect 74214 59470 74980 59530
rect 75502 59606 76544 59666
rect 76649 59666 76715 59669
rect 77312 59666 77372 60044
rect 76649 59664 77372 59666
rect 76649 59608 76654 59664
rect 76710 59608 77372 59664
rect 76649 59606 77372 59608
rect 77477 59666 77543 59669
rect 78140 59666 78200 60044
rect 77477 59664 78200 59666
rect 77477 59608 77482 59664
rect 77538 59608 78200 59664
rect 77477 59606 78200 59608
rect 70301 59331 70367 59334
rect 67265 59256 68570 59258
rect 67265 59200 67270 59256
rect 67326 59200 68570 59256
rect 67265 59198 68570 59200
rect 71405 59258 71471 59261
rect 72558 59258 72618 59334
rect 71405 59256 72618 59258
rect 71405 59200 71410 59256
rect 71466 59200 72618 59256
rect 71405 59198 72618 59200
rect 67265 59195 67331 59198
rect 71405 59195 71471 59198
rect 71589 59122 71655 59125
rect 73478 59122 73538 59334
rect 71589 59120 73538 59122
rect 71589 59064 71594 59120
rect 71650 59064 73538 59120
rect 71589 59062 73538 59064
rect 71589 59059 71655 59062
rect 72969 58986 73035 58989
rect 74214 58986 74274 59470
rect 74441 59394 74507 59397
rect 75502 59394 75562 59606
rect 76649 59603 76715 59606
rect 77477 59603 77543 59606
rect 76557 59530 76623 59533
rect 78968 59530 79028 60044
rect 79796 59802 79856 60044
rect 76557 59528 79028 59530
rect 76557 59472 76562 59528
rect 76618 59472 79028 59528
rect 76557 59470 79028 59472
rect 79182 59742 79856 59802
rect 79961 59802 80027 59805
rect 80624 59802 80684 60044
rect 79961 59800 80684 59802
rect 79961 59744 79966 59800
rect 80022 59744 80684 59800
rect 79961 59742 80684 59744
rect 76557 59467 76623 59470
rect 76649 59394 76715 59397
rect 74441 59392 75562 59394
rect 74441 59336 74446 59392
rect 74502 59336 75562 59392
rect 74441 59334 75562 59336
rect 75686 59392 76715 59394
rect 75686 59336 76654 59392
rect 76710 59336 76715 59392
rect 75686 59334 76715 59336
rect 74441 59331 74507 59334
rect 75177 59258 75243 59261
rect 75686 59258 75746 59334
rect 76649 59331 76715 59334
rect 76833 59394 76899 59397
rect 79182 59394 79242 59742
rect 79961 59739 80027 59742
rect 79317 59666 79383 59669
rect 81452 59666 81512 60044
rect 79317 59664 81512 59666
rect 79317 59608 79322 59664
rect 79378 59608 81512 59664
rect 79317 59606 81512 59608
rect 81617 59666 81683 59669
rect 82280 59666 82340 60044
rect 81617 59664 82340 59666
rect 81617 59608 81622 59664
rect 81678 59608 82340 59664
rect 81617 59606 82340 59608
rect 79317 59603 79383 59606
rect 81617 59603 81683 59606
rect 80697 59530 80763 59533
rect 83108 59530 83168 60044
rect 83273 59666 83339 59669
rect 83936 59666 83996 60044
rect 84193 59802 84259 59805
rect 84764 59802 84824 60044
rect 84193 59800 84824 59802
rect 84193 59744 84198 59800
rect 84254 59744 84824 59800
rect 84193 59742 84824 59744
rect 84193 59739 84259 59742
rect 83273 59664 83996 59666
rect 83273 59608 83278 59664
rect 83334 59608 83996 59664
rect 83273 59606 83996 59608
rect 84101 59666 84167 59669
rect 85592 59666 85652 60044
rect 84101 59664 85652 59666
rect 84101 59608 84106 59664
rect 84162 59608 85652 59664
rect 84101 59606 85652 59608
rect 85757 59666 85823 59669
rect 86420 59666 86480 60044
rect 85757 59664 86480 59666
rect 85757 59608 85762 59664
rect 85818 59608 86480 59664
rect 85757 59606 86480 59608
rect 83273 59603 83339 59606
rect 84101 59603 84167 59606
rect 85757 59603 85823 59606
rect 80697 59528 83168 59530
rect 80697 59472 80702 59528
rect 80758 59472 83168 59528
rect 80697 59470 83168 59472
rect 84837 59530 84903 59533
rect 87248 59530 87308 60044
rect 84837 59528 87308 59530
rect 84837 59472 84842 59528
rect 84898 59472 87308 59528
rect 84837 59470 87308 59472
rect 87413 59530 87479 59533
rect 88076 59530 88136 60044
rect 87413 59528 88136 59530
rect 87413 59472 87418 59528
rect 87474 59472 88136 59528
rect 87413 59470 88136 59472
rect 80697 59467 80763 59470
rect 84837 59467 84903 59470
rect 87413 59467 87479 59470
rect 76833 59392 79242 59394
rect 76833 59336 76838 59392
rect 76894 59336 79242 59392
rect 76833 59334 79242 59336
rect 79501 59394 79567 59397
rect 81617 59394 81683 59397
rect 79501 59392 81683 59394
rect 79501 59336 79506 59392
rect 79562 59336 81622 59392
rect 81678 59336 81683 59392
rect 79501 59334 81683 59336
rect 76833 59331 76899 59334
rect 79501 59331 79567 59334
rect 81617 59331 81683 59334
rect 83641 59394 83707 59397
rect 85757 59394 85823 59397
rect 83641 59392 85823 59394
rect 83641 59336 83646 59392
rect 83702 59336 85762 59392
rect 85818 59336 85823 59392
rect 83641 59334 85823 59336
rect 83641 59331 83707 59334
rect 85757 59331 85823 59334
rect 86217 59394 86283 59397
rect 88904 59394 88964 60044
rect 89069 59666 89135 59669
rect 89732 59666 89792 60044
rect 89069 59664 89792 59666
rect 89069 59608 89074 59664
rect 89130 59608 89792 59664
rect 89069 59606 89792 59608
rect 89897 59666 89963 59669
rect 90560 59666 90620 60044
rect 89897 59664 90620 59666
rect 89897 59608 89902 59664
rect 89958 59608 90620 59664
rect 89897 59606 90620 59608
rect 89069 59603 89135 59606
rect 89897 59603 89963 59606
rect 89621 59530 89687 59533
rect 91388 59530 91448 60044
rect 89621 59528 91448 59530
rect 89621 59472 89626 59528
rect 89682 59472 91448 59528
rect 89621 59470 91448 59472
rect 91553 59530 91619 59533
rect 92216 59530 92276 60044
rect 91553 59528 92276 59530
rect 91553 59472 91558 59528
rect 91614 59472 92276 59528
rect 91553 59470 92276 59472
rect 89621 59467 89687 59470
rect 91553 59467 91619 59470
rect 89897 59394 89963 59397
rect 86217 59392 88964 59394
rect 86217 59336 86222 59392
rect 86278 59336 88964 59392
rect 86217 59334 88964 59336
rect 89118 59392 89963 59394
rect 89118 59336 89902 59392
rect 89958 59336 89963 59392
rect 89118 59334 89963 59336
rect 86217 59331 86283 59334
rect 75177 59256 75746 59258
rect 75177 59200 75182 59256
rect 75238 59200 75746 59256
rect 75177 59198 75746 59200
rect 87781 59258 87847 59261
rect 89118 59258 89178 59334
rect 89897 59331 89963 59334
rect 90725 59394 90791 59397
rect 92952 59394 93012 60044
rect 93780 59938 93840 60044
rect 90725 59392 93012 59394
rect 90725 59336 90730 59392
rect 90786 59336 93012 59392
rect 90725 59334 93012 59336
rect 93166 59878 93840 59938
rect 90725 59331 90791 59334
rect 87781 59256 89178 59258
rect 87781 59200 87786 59256
rect 87842 59200 89178 59256
rect 87781 59198 89178 59200
rect 90909 59258 90975 59261
rect 93166 59258 93226 59878
rect 93853 59802 93919 59805
rect 94608 59802 94668 60044
rect 93853 59800 94668 59802
rect 93853 59744 93858 59800
rect 93914 59744 94668 59800
rect 93853 59742 94668 59744
rect 93853 59739 93919 59742
rect 95436 59669 95496 60044
rect 95417 59664 95496 59669
rect 95417 59608 95422 59664
rect 95478 59608 95496 59664
rect 95417 59606 95496 59608
rect 95417 59603 95483 59606
rect 93761 59530 93827 59533
rect 96264 59530 96324 60044
rect 93761 59528 96324 59530
rect 93761 59472 93766 59528
rect 93822 59472 96324 59528
rect 93761 59470 96324 59472
rect 93761 59467 93827 59470
rect 93669 59394 93735 59397
rect 95417 59394 95483 59397
rect 97092 59394 97152 60044
rect 97920 59938 97980 60044
rect 93669 59392 95483 59394
rect 93669 59336 93674 59392
rect 93730 59336 95422 59392
rect 95478 59336 95483 59392
rect 93669 59334 95483 59336
rect 93669 59331 93735 59334
rect 95417 59331 95483 59334
rect 95558 59334 97152 59394
rect 97214 59878 97980 59938
rect 90909 59256 93226 59258
rect 90909 59200 90914 59256
rect 90970 59200 93226 59256
rect 90909 59198 93226 59200
rect 95141 59258 95207 59261
rect 95558 59258 95618 59334
rect 95141 59256 95618 59258
rect 95141 59200 95146 59256
rect 95202 59200 95618 59256
rect 95141 59198 95618 59200
rect 75177 59195 75243 59198
rect 87781 59195 87847 59198
rect 90909 59195 90975 59198
rect 95141 59195 95207 59198
rect 93853 59122 93919 59125
rect 97214 59122 97274 59878
rect 97349 59802 97415 59805
rect 98748 59802 98808 60044
rect 97349 59800 98808 59802
rect 97349 59744 97354 59800
rect 97410 59744 98808 59800
rect 97349 59742 98808 59744
rect 97349 59739 97415 59742
rect 97441 59666 97507 59669
rect 99576 59666 99636 60044
rect 97441 59664 99636 59666
rect 97441 59608 97446 59664
rect 97502 59608 99636 59664
rect 97441 59606 99636 59608
rect 99741 59666 99807 59669
rect 100404 59666 100464 60044
rect 99741 59664 100464 59666
rect 99741 59608 99746 59664
rect 99802 59608 100464 59664
rect 99741 59606 100464 59608
rect 97441 59603 97507 59606
rect 99741 59603 99807 59606
rect 98821 59530 98887 59533
rect 101232 59530 101292 60044
rect 101397 59802 101463 59805
rect 102060 59802 102120 60044
rect 102888 59802 102948 60044
rect 101397 59800 102120 59802
rect 101397 59744 101402 59800
rect 101458 59744 102120 59800
rect 101397 59742 102120 59744
rect 102182 59742 102948 59802
rect 101397 59739 101463 59742
rect 102182 59666 102242 59742
rect 103716 59666 103776 60044
rect 98821 59528 101292 59530
rect 98821 59472 98826 59528
rect 98882 59472 101292 59528
rect 98821 59470 101292 59472
rect 101446 59606 102242 59666
rect 102918 59606 103776 59666
rect 103973 59666 104039 59669
rect 104544 59666 104604 60044
rect 103973 59664 104604 59666
rect 103973 59608 103978 59664
rect 104034 59608 104604 59664
rect 103973 59606 104604 59608
rect 98821 59467 98887 59470
rect 97349 59394 97415 59397
rect 99741 59394 99807 59397
rect 97349 59392 99807 59394
rect 97349 59336 97354 59392
rect 97410 59336 99746 59392
rect 99802 59336 99807 59392
rect 97349 59334 99807 59336
rect 97349 59331 97415 59334
rect 99741 59331 99807 59334
rect 100017 59394 100083 59397
rect 101446 59394 101506 59606
rect 101581 59530 101647 59533
rect 102918 59530 102978 59606
rect 103973 59603 104039 59606
rect 101581 59528 102978 59530
rect 101581 59472 101586 59528
rect 101642 59472 102978 59528
rect 101581 59470 102978 59472
rect 103145 59530 103211 59533
rect 105372 59530 105432 60044
rect 105629 59802 105695 59805
rect 106200 59802 106260 60044
rect 107028 59802 107088 60044
rect 105629 59800 106260 59802
rect 105629 59744 105634 59800
rect 105690 59744 106260 59800
rect 105629 59742 106260 59744
rect 106414 59742 107088 59802
rect 107193 59802 107259 59805
rect 107856 59802 107916 60044
rect 107193 59800 107916 59802
rect 107193 59744 107198 59800
rect 107254 59744 107916 59800
rect 107193 59742 107916 59744
rect 108021 59802 108087 59805
rect 108684 59802 108744 60044
rect 108021 59800 108744 59802
rect 108021 59744 108026 59800
rect 108082 59744 108744 59800
rect 108021 59742 108744 59744
rect 108849 59802 108915 59805
rect 109420 59802 109480 60044
rect 108849 59800 109480 59802
rect 108849 59744 108854 59800
rect 108910 59744 109480 59800
rect 108849 59742 109480 59744
rect 105629 59739 105695 59742
rect 106414 59666 106474 59742
rect 107193 59739 107259 59742
rect 108021 59739 108087 59742
rect 108849 59739 108915 59742
rect 103145 59528 105432 59530
rect 103145 59472 103150 59528
rect 103206 59472 105432 59528
rect 103145 59470 105432 59472
rect 105494 59606 106474 59666
rect 107101 59666 107167 59669
rect 110248 59666 110308 60044
rect 111076 59938 111136 60044
rect 107101 59664 110308 59666
rect 107101 59608 107106 59664
rect 107162 59608 110308 59664
rect 107101 59606 110308 59608
rect 110462 59878 111136 59938
rect 101581 59467 101647 59470
rect 103145 59467 103211 59470
rect 100017 59392 101506 59394
rect 100017 59336 100022 59392
rect 100078 59336 101506 59392
rect 100017 59334 101506 59336
rect 101581 59394 101647 59397
rect 103973 59394 104039 59397
rect 105494 59394 105554 59606
rect 107101 59603 107167 59606
rect 105721 59530 105787 59533
rect 107193 59530 107259 59533
rect 105721 59528 107259 59530
rect 105721 59472 105726 59528
rect 105782 59472 107198 59528
rect 107254 59472 107259 59528
rect 105721 59470 107259 59472
rect 105721 59467 105787 59470
rect 107193 59467 107259 59470
rect 108297 59530 108363 59533
rect 110462 59530 110522 59878
rect 111333 59802 111399 59805
rect 111904 59802 111964 60044
rect 111333 59800 111964 59802
rect 111333 59744 111338 59800
rect 111394 59744 111964 59800
rect 111333 59742 111964 59744
rect 111333 59739 111399 59742
rect 111333 59666 111399 59669
rect 112732 59666 112792 60044
rect 111333 59664 112792 59666
rect 111333 59608 111338 59664
rect 111394 59608 112792 59664
rect 111333 59606 112792 59608
rect 111333 59603 111399 59606
rect 108297 59528 110522 59530
rect 108297 59472 108302 59528
rect 108358 59472 110522 59528
rect 108297 59470 110522 59472
rect 111241 59530 111307 59533
rect 113560 59530 113620 60044
rect 113725 59802 113791 59805
rect 114388 59802 114448 60044
rect 113725 59800 114448 59802
rect 113725 59744 113730 59800
rect 113786 59744 114448 59800
rect 113725 59742 114448 59744
rect 113725 59739 113791 59742
rect 114185 59666 114251 59669
rect 115216 59666 115276 60044
rect 114185 59664 115276 59666
rect 114185 59608 114190 59664
rect 114246 59608 115276 59664
rect 114185 59606 115276 59608
rect 114185 59603 114251 59606
rect 111241 59528 113620 59530
rect 111241 59472 111246 59528
rect 111302 59472 113620 59528
rect 111241 59470 113620 59472
rect 113817 59530 113883 59533
rect 116044 59530 116104 60044
rect 116209 59802 116275 59805
rect 116872 59802 116932 60044
rect 116209 59800 116932 59802
rect 116209 59744 116214 59800
rect 116270 59744 116932 59800
rect 116209 59742 116932 59744
rect 116209 59739 116275 59742
rect 117700 59666 117760 60044
rect 113817 59528 116104 59530
rect 113817 59472 113822 59528
rect 113878 59472 116104 59528
rect 113817 59470 116104 59472
rect 116166 59606 117760 59666
rect 117865 59666 117931 59669
rect 118528 59666 118588 60044
rect 117865 59664 118588 59666
rect 117865 59608 117870 59664
rect 117926 59608 118588 59664
rect 117865 59606 118588 59608
rect 108297 59467 108363 59470
rect 111241 59467 111307 59470
rect 113817 59467 113883 59470
rect 101581 59392 104039 59394
rect 101581 59336 101586 59392
rect 101642 59336 103978 59392
rect 104034 59336 104039 59392
rect 101581 59334 104039 59336
rect 100017 59331 100083 59334
rect 101581 59331 101647 59334
rect 103973 59331 104039 59334
rect 104758 59334 105554 59394
rect 106917 59394 106983 59397
rect 108849 59394 108915 59397
rect 106917 59392 108915 59394
rect 106917 59336 106922 59392
rect 106978 59336 108854 59392
rect 108910 59336 108915 59392
rect 106917 59334 108915 59336
rect 104157 59258 104223 59261
rect 104758 59258 104818 59334
rect 106917 59331 106983 59334
rect 108849 59331 108915 59334
rect 109677 59394 109743 59397
rect 111333 59394 111399 59397
rect 109677 59392 111399 59394
rect 109677 59336 109682 59392
rect 109738 59336 111338 59392
rect 111394 59336 111399 59392
rect 109677 59334 111399 59336
rect 109677 59331 109743 59334
rect 111333 59331 111399 59334
rect 112437 59394 112503 59397
rect 114185 59394 114251 59397
rect 112437 59392 114251 59394
rect 112437 59336 112442 59392
rect 112498 59336 114190 59392
rect 114246 59336 114251 59392
rect 112437 59334 114251 59336
rect 112437 59331 112503 59334
rect 114185 59331 114251 59334
rect 115381 59394 115447 59397
rect 116166 59394 116226 59606
rect 117865 59603 117931 59606
rect 117221 59530 117287 59533
rect 119356 59530 119416 60044
rect 117221 59528 119416 59530
rect 117221 59472 117226 59528
rect 117282 59472 119416 59528
rect 117221 59470 119416 59472
rect 117221 59467 117287 59470
rect 117773 59394 117839 59397
rect 115381 59392 116226 59394
rect 115381 59336 115386 59392
rect 115442 59336 116226 59392
rect 115381 59334 116226 59336
rect 116350 59392 117839 59394
rect 116350 59336 117778 59392
rect 117834 59336 117839 59392
rect 116350 59334 117839 59336
rect 115381 59331 115447 59334
rect 104157 59256 104818 59258
rect 104157 59200 104162 59256
rect 104218 59200 104818 59256
rect 104157 59198 104818 59200
rect 115841 59258 115907 59261
rect 116350 59258 116410 59334
rect 117773 59331 117839 59334
rect 117957 59394 118023 59397
rect 120184 59394 120244 60044
rect 120349 59666 120415 59669
rect 121012 59666 121072 60044
rect 120349 59664 121072 59666
rect 120349 59608 120354 59664
rect 120410 59608 121072 59664
rect 120349 59606 121072 59608
rect 120349 59603 120415 59606
rect 121840 59530 121900 60044
rect 122005 59802 122071 59805
rect 122668 59802 122728 60044
rect 122005 59800 122728 59802
rect 122005 59744 122010 59800
rect 122066 59744 122728 59800
rect 122005 59742 122728 59744
rect 123109 59802 123175 59805
rect 123496 59802 123556 60044
rect 123109 59800 123556 59802
rect 123109 59744 123114 59800
rect 123170 59744 123556 59800
rect 123109 59742 123556 59744
rect 122005 59739 122071 59742
rect 123109 59739 123175 59742
rect 122281 59666 122347 59669
rect 123293 59666 123359 59669
rect 122281 59664 123359 59666
rect 122281 59608 122286 59664
rect 122342 59608 123298 59664
rect 123354 59608 123359 59664
rect 122281 59606 123359 59608
rect 122281 59603 122347 59606
rect 123293 59603 123359 59606
rect 117957 59392 120244 59394
rect 117957 59336 117962 59392
rect 118018 59336 120244 59392
rect 117957 59334 120244 59336
rect 120398 59470 121900 59530
rect 122097 59530 122163 59533
rect 124324 59530 124384 60044
rect 122097 59528 124384 59530
rect 122097 59472 122102 59528
rect 122158 59472 124384 59528
rect 122097 59470 124384 59472
rect 117957 59331 118023 59334
rect 115841 59256 116410 59258
rect 115841 59200 115846 59256
rect 115902 59200 116410 59256
rect 115841 59198 116410 59200
rect 119337 59258 119403 59261
rect 120398 59258 120458 59470
rect 122097 59467 122163 59470
rect 120717 59394 120783 59397
rect 123109 59394 123175 59397
rect 120717 59392 123175 59394
rect 120717 59336 120722 59392
rect 120778 59336 123114 59392
rect 123170 59336 123175 59392
rect 120717 59334 123175 59336
rect 120717 59331 120783 59334
rect 123109 59331 123175 59334
rect 123661 59394 123727 59397
rect 125060 59394 125120 60044
rect 125888 59394 125948 60044
rect 126716 59938 126776 60044
rect 126286 59878 126776 59938
rect 126286 59669 126346 59878
rect 126421 59802 126487 59805
rect 127544 59802 127604 60044
rect 126421 59800 127604 59802
rect 126421 59744 126426 59800
rect 126482 59744 127604 59800
rect 126421 59742 127604 59744
rect 126421 59739 126487 59742
rect 126237 59664 126346 59669
rect 126237 59608 126242 59664
rect 126298 59608 126346 59664
rect 126237 59606 126346 59608
rect 126421 59666 126487 59669
rect 128372 59666 128432 60044
rect 126421 59664 128432 59666
rect 126421 59608 126426 59664
rect 126482 59608 128432 59664
rect 126421 59606 128432 59608
rect 128537 59666 128603 59669
rect 129200 59666 129260 60044
rect 128537 59664 129260 59666
rect 128537 59608 128542 59664
rect 128598 59608 129260 59664
rect 128537 59606 129260 59608
rect 126237 59603 126303 59606
rect 126421 59603 126487 59606
rect 128537 59603 128603 59606
rect 127801 59530 127867 59533
rect 130028 59530 130088 60044
rect 130856 59938 130916 60044
rect 130334 59878 130916 59938
rect 130193 59802 130259 59805
rect 130334 59802 130394 59878
rect 130193 59800 130394 59802
rect 130193 59744 130198 59800
rect 130254 59744 130394 59800
rect 130193 59742 130394 59744
rect 131021 59802 131087 59805
rect 131684 59802 131744 60044
rect 132512 59938 132572 60044
rect 131021 59800 131744 59802
rect 131021 59744 131026 59800
rect 131082 59744 131744 59800
rect 131021 59742 131744 59744
rect 131806 59878 132572 59938
rect 130193 59739 130259 59742
rect 131021 59739 131087 59742
rect 127801 59528 130088 59530
rect 127801 59472 127806 59528
rect 127862 59472 130088 59528
rect 127801 59470 130088 59472
rect 130377 59530 130443 59533
rect 131806 59530 131866 59878
rect 132033 59802 132099 59805
rect 133137 59802 133203 59805
rect 132033 59800 133203 59802
rect 132033 59744 132038 59800
rect 132094 59744 133142 59800
rect 133198 59744 133203 59800
rect 132033 59742 133203 59744
rect 132033 59739 132099 59742
rect 133137 59739 133203 59742
rect 131941 59666 132007 59669
rect 133340 59666 133400 60044
rect 133505 59802 133571 59805
rect 134168 59802 134228 60044
rect 133505 59800 134228 59802
rect 133505 59744 133510 59800
rect 133566 59744 134228 59800
rect 133505 59742 134228 59744
rect 134333 59802 134399 59805
rect 134996 59802 135056 60044
rect 134333 59800 135056 59802
rect 134333 59744 134338 59800
rect 134394 59744 135056 59800
rect 134333 59742 135056 59744
rect 135253 59802 135319 59805
rect 135824 59802 135884 60044
rect 135253 59800 135884 59802
rect 135253 59744 135258 59800
rect 135314 59744 135884 59800
rect 135253 59742 135884 59744
rect 133505 59739 133571 59742
rect 134333 59739 134399 59742
rect 135253 59739 135319 59742
rect 131941 59664 133400 59666
rect 131941 59608 131946 59664
rect 132002 59608 133400 59664
rect 131941 59606 133400 59608
rect 135161 59666 135227 59669
rect 136652 59666 136712 60044
rect 135161 59664 136712 59666
rect 135161 59608 135166 59664
rect 135222 59608 136712 59664
rect 135161 59606 136712 59608
rect 136817 59666 136883 59669
rect 137480 59666 137540 60044
rect 136817 59664 137540 59666
rect 136817 59608 136822 59664
rect 136878 59608 137540 59664
rect 136817 59606 137540 59608
rect 131941 59603 132007 59606
rect 135161 59603 135227 59606
rect 136817 59603 136883 59606
rect 130377 59528 131866 59530
rect 130377 59472 130382 59528
rect 130438 59472 131866 59528
rect 130377 59470 131866 59472
rect 133137 59530 133203 59533
rect 135253 59530 135319 59533
rect 133137 59528 135319 59530
rect 133137 59472 133142 59528
rect 133198 59472 135258 59528
rect 135314 59472 135319 59528
rect 133137 59470 135319 59472
rect 127801 59467 127867 59470
rect 130377 59467 130443 59470
rect 133137 59467 133203 59470
rect 135253 59467 135319 59470
rect 135897 59530 135963 59533
rect 138308 59530 138368 60044
rect 135897 59528 138368 59530
rect 135897 59472 135902 59528
rect 135958 59472 138368 59528
rect 135897 59470 138368 59472
rect 135897 59467 135963 59470
rect 123661 59392 125120 59394
rect 123661 59336 123666 59392
rect 123722 59336 125120 59392
rect 123661 59334 125120 59336
rect 125182 59334 125948 59394
rect 126237 59394 126303 59397
rect 128537 59394 128603 59397
rect 126237 59392 128603 59394
rect 126237 59336 126242 59392
rect 126298 59336 128542 59392
rect 128598 59336 128603 59392
rect 126237 59334 128603 59336
rect 123661 59331 123727 59334
rect 119337 59256 120458 59258
rect 119337 59200 119342 59256
rect 119398 59200 120458 59256
rect 119337 59198 120458 59200
rect 123661 59258 123727 59261
rect 125182 59258 125242 59334
rect 126237 59331 126303 59334
rect 128537 59331 128603 59334
rect 128997 59394 129063 59397
rect 130653 59394 130719 59397
rect 128997 59392 130719 59394
rect 128997 59336 129002 59392
rect 129058 59336 130658 59392
rect 130714 59336 130719 59392
rect 128997 59334 130719 59336
rect 128997 59331 129063 59334
rect 130653 59331 130719 59334
rect 131113 59394 131179 59397
rect 134333 59394 134399 59397
rect 136817 59394 136883 59397
rect 131113 59392 134399 59394
rect 131113 59336 131118 59392
rect 131174 59336 134338 59392
rect 134394 59336 134399 59392
rect 131113 59334 134399 59336
rect 131113 59331 131179 59334
rect 134333 59331 134399 59334
rect 135118 59392 136883 59394
rect 135118 59336 136822 59392
rect 136878 59336 136883 59392
rect 135118 59334 136883 59336
rect 123661 59256 125242 59258
rect 123661 59200 123666 59256
rect 123722 59200 125242 59256
rect 123661 59198 125242 59200
rect 134701 59258 134767 59261
rect 135118 59258 135178 59334
rect 136817 59331 136883 59334
rect 137369 59394 137435 59397
rect 138105 59394 138171 59397
rect 139136 59394 139196 60044
rect 139301 59530 139367 59533
rect 139964 59530 140024 60044
rect 139301 59528 140024 59530
rect 139301 59472 139306 59528
rect 139362 59472 140024 59528
rect 139301 59470 140024 59472
rect 139301 59467 139367 59470
rect 140792 59394 140852 60044
rect 141528 59666 141588 60044
rect 141693 59802 141759 59805
rect 142356 59802 142416 60044
rect 141693 59800 142416 59802
rect 141693 59744 141698 59800
rect 141754 59744 142416 59800
rect 141693 59742 142416 59744
rect 141693 59739 141759 59742
rect 137369 59392 138171 59394
rect 137369 59336 137374 59392
rect 137430 59336 138110 59392
rect 138166 59336 138171 59392
rect 137369 59334 138171 59336
rect 137369 59331 137435 59334
rect 138105 59331 138171 59334
rect 138246 59334 139196 59394
rect 139350 59334 140852 59394
rect 141006 59606 141588 59666
rect 141693 59666 141759 59669
rect 143184 59666 143244 60044
rect 141693 59664 143244 59666
rect 141693 59608 141698 59664
rect 141754 59608 143244 59664
rect 141693 59606 143244 59608
rect 134701 59256 135178 59258
rect 134701 59200 134706 59256
rect 134762 59200 135178 59256
rect 134701 59198 135178 59200
rect 136081 59258 136147 59261
rect 138246 59258 138306 59334
rect 136081 59256 138306 59258
rect 136081 59200 136086 59256
rect 136142 59200 138306 59256
rect 136081 59198 138306 59200
rect 138657 59258 138723 59261
rect 139350 59258 139410 59334
rect 138657 59256 139410 59258
rect 138657 59200 138662 59256
rect 138718 59200 139410 59256
rect 138657 59198 139410 59200
rect 104157 59195 104223 59198
rect 115841 59195 115907 59198
rect 119337 59195 119403 59198
rect 123661 59195 123727 59198
rect 134701 59195 134767 59198
rect 136081 59195 136147 59198
rect 138657 59195 138723 59198
rect 93853 59120 97274 59122
rect 93853 59064 93858 59120
rect 93914 59064 97274 59120
rect 93853 59062 97274 59064
rect 138841 59122 138907 59125
rect 141006 59122 141066 59606
rect 141693 59603 141759 59606
rect 141509 59530 141575 59533
rect 144012 59530 144072 60044
rect 144840 59938 144900 60044
rect 141509 59528 144072 59530
rect 141509 59472 141514 59528
rect 141570 59472 144072 59528
rect 141509 59470 144072 59472
rect 144318 59878 144900 59938
rect 141509 59467 141575 59470
rect 142889 59394 142955 59397
rect 144177 59394 144243 59397
rect 142889 59392 144243 59394
rect 142889 59336 142894 59392
rect 142950 59336 144182 59392
rect 144238 59336 144243 59392
rect 142889 59334 144243 59336
rect 142889 59331 142955 59334
rect 144177 59331 144243 59334
rect 142061 59258 142127 59261
rect 144318 59258 144378 59878
rect 144453 59802 144519 59805
rect 145668 59802 145728 60044
rect 144453 59800 145728 59802
rect 144453 59744 144458 59800
rect 144514 59744 145728 59800
rect 144453 59742 145728 59744
rect 145833 59802 145899 59805
rect 146496 59802 146556 60044
rect 145833 59800 146556 59802
rect 145833 59744 145838 59800
rect 145894 59744 146556 59800
rect 145833 59742 146556 59744
rect 144453 59739 144519 59742
rect 145833 59739 145899 59742
rect 144545 59666 144611 59669
rect 147324 59666 147384 60044
rect 144545 59664 147384 59666
rect 144545 59608 144550 59664
rect 144606 59608 147384 59664
rect 144545 59606 147384 59608
rect 144545 59603 144611 59606
rect 144729 59530 144795 59533
rect 145833 59530 145899 59533
rect 144729 59528 145899 59530
rect 144729 59472 144734 59528
rect 144790 59472 145838 59528
rect 145894 59472 145899 59528
rect 144729 59470 145899 59472
rect 144729 59467 144795 59470
rect 145833 59467 145899 59470
rect 146201 59394 146267 59397
rect 148152 59394 148212 60044
rect 149808 59938 149868 60044
rect 148688 59878 149868 59938
rect 148688 59805 148748 59878
rect 148685 59800 148751 59805
rect 148685 59744 148690 59800
rect 148746 59744 148751 59800
rect 148685 59739 148751 59744
rect 149973 59530 150039 59533
rect 150636 59530 150696 60044
rect 151464 59938 151524 60044
rect 149973 59528 150696 59530
rect 149973 59472 149978 59528
rect 150034 59472 150696 59528
rect 149973 59470 150696 59472
rect 150758 59878 151524 59938
rect 149973 59467 150039 59470
rect 150758 59394 150818 59878
rect 151905 59802 151971 59805
rect 152292 59802 152352 60044
rect 153120 59938 153180 60044
rect 151905 59800 152352 59802
rect 151905 59744 151910 59800
rect 151966 59744 152352 59800
rect 151905 59742 152352 59744
rect 152414 59878 153180 59938
rect 151905 59739 151971 59742
rect 151629 59666 151695 59669
rect 152414 59666 152474 59878
rect 153948 59802 154008 60044
rect 151629 59664 152474 59666
rect 151629 59608 151634 59664
rect 151690 59608 152474 59664
rect 151629 59606 152474 59608
rect 152598 59742 154008 59802
rect 151629 59603 151695 59606
rect 151721 59530 151787 59533
rect 152598 59530 152658 59742
rect 152825 59666 152891 59669
rect 154776 59666 154836 60044
rect 152825 59664 154836 59666
rect 152825 59608 152830 59664
rect 152886 59608 154836 59664
rect 152825 59606 154836 59608
rect 154941 59666 155007 59669
rect 155604 59666 155664 60044
rect 154941 59664 155664 59666
rect 154941 59608 154946 59664
rect 155002 59608 155664 59664
rect 154941 59606 155664 59608
rect 152825 59603 152891 59606
rect 154941 59603 155007 59606
rect 151721 59528 152658 59530
rect 151721 59472 151726 59528
rect 151782 59472 152658 59528
rect 151721 59470 152658 59472
rect 154297 59530 154363 59533
rect 156432 59530 156492 60044
rect 157260 59669 157320 60044
rect 157241 59664 157320 59669
rect 157241 59608 157246 59664
rect 157302 59608 157320 59664
rect 157241 59606 157320 59608
rect 157609 59666 157675 59669
rect 157996 59666 158056 60044
rect 158161 59802 158227 59805
rect 158824 59802 158884 60044
rect 158161 59800 158884 59802
rect 158161 59744 158166 59800
rect 158222 59744 158884 59800
rect 158161 59742 158884 59744
rect 158161 59739 158227 59742
rect 159652 59666 159712 60044
rect 157609 59664 158056 59666
rect 157609 59608 157614 59664
rect 157670 59608 158056 59664
rect 157609 59606 158056 59608
rect 158118 59606 159712 59666
rect 157241 59603 157307 59606
rect 157609 59603 157675 59606
rect 154297 59528 156492 59530
rect 154297 59472 154302 59528
rect 154358 59472 156492 59528
rect 154297 59470 156492 59472
rect 156965 59530 157031 59533
rect 156965 59528 157810 59530
rect 156965 59472 156970 59528
rect 157026 59472 157810 59528
rect 156965 59470 157810 59472
rect 151721 59467 151787 59470
rect 154297 59467 154363 59470
rect 156965 59467 157031 59470
rect 146201 59392 148212 59394
rect 146201 59336 146206 59392
rect 146262 59336 148212 59392
rect 146201 59334 148212 59336
rect 150022 59334 150818 59394
rect 153009 59394 153075 59397
rect 154941 59394 155007 59397
rect 153009 59392 155007 59394
rect 153009 59336 153014 59392
rect 153070 59336 154946 59392
rect 155002 59336 155007 59392
rect 153009 59334 155007 59336
rect 146201 59331 146267 59334
rect 142061 59256 144378 59258
rect 142061 59200 142066 59256
rect 142122 59200 144378 59256
rect 142061 59198 144378 59200
rect 148869 59258 148935 59261
rect 150022 59258 150082 59334
rect 153009 59331 153075 59334
rect 154941 59331 155007 59334
rect 155861 59394 155927 59397
rect 157609 59394 157675 59397
rect 155861 59392 157675 59394
rect 155861 59336 155866 59392
rect 155922 59336 157614 59392
rect 157670 59336 157675 59392
rect 155861 59334 157675 59336
rect 157750 59394 157810 59470
rect 158118 59394 158178 59606
rect 158345 59530 158411 59533
rect 160480 59530 160540 60044
rect 161308 59666 161368 60044
rect 158345 59528 160540 59530
rect 158345 59472 158350 59528
rect 158406 59472 160540 59528
rect 158345 59470 160540 59472
rect 160694 59606 161368 59666
rect 162136 59666 162196 60044
rect 162761 59666 162827 59669
rect 162136 59664 162827 59666
rect 162136 59608 162766 59664
rect 162822 59608 162827 59664
rect 162136 59606 162827 59608
rect 158345 59467 158411 59470
rect 157750 59334 158178 59394
rect 158621 59394 158687 59397
rect 160694 59394 160754 59606
rect 162761 59603 162827 59606
rect 161197 59530 161263 59533
rect 162964 59530 163024 60044
rect 163792 59802 163852 60044
rect 164049 59802 164115 59805
rect 163792 59800 164115 59802
rect 163792 59744 164054 59800
rect 164110 59744 164115 59800
rect 163792 59742 164115 59744
rect 164049 59739 164115 59742
rect 164620 59666 164680 60044
rect 161197 59528 163024 59530
rect 161197 59472 161202 59528
rect 161258 59472 163024 59528
rect 161197 59470 163024 59472
rect 163086 59606 164680 59666
rect 164785 59666 164851 59669
rect 165448 59666 165508 60044
rect 164785 59664 165508 59666
rect 164785 59608 164790 59664
rect 164846 59608 165508 59664
rect 164785 59606 165508 59608
rect 161197 59467 161263 59470
rect 158621 59392 160754 59394
rect 158621 59336 158626 59392
rect 158682 59336 160754 59392
rect 158621 59334 160754 59336
rect 162485 59394 162551 59397
rect 163086 59394 163146 59606
rect 164785 59603 164851 59606
rect 164141 59530 164207 59533
rect 166276 59530 166336 60044
rect 166441 59666 166507 59669
rect 167104 59666 167164 60044
rect 166441 59664 167164 59666
rect 166441 59608 166446 59664
rect 166502 59608 167164 59664
rect 166441 59606 167164 59608
rect 167269 59666 167335 59669
rect 167932 59666 167992 60044
rect 167269 59664 167992 59666
rect 167269 59608 167274 59664
rect 167330 59608 167992 59664
rect 167269 59606 167992 59608
rect 166441 59603 166507 59606
rect 167269 59603 167335 59606
rect 164141 59528 166336 59530
rect 164141 59472 164146 59528
rect 164202 59472 166336 59528
rect 164141 59470 166336 59472
rect 166809 59530 166875 59533
rect 168760 59530 168820 60044
rect 166809 59528 168820 59530
rect 166809 59472 166814 59528
rect 166870 59472 168820 59528
rect 166809 59470 168820 59472
rect 168925 59530 168991 59533
rect 169588 59530 169648 60044
rect 168925 59528 169648 59530
rect 168925 59472 168930 59528
rect 168986 59472 169648 59528
rect 168925 59470 169648 59472
rect 164141 59467 164207 59470
rect 166809 59467 166875 59470
rect 168925 59467 168991 59470
rect 164785 59394 164851 59397
rect 162485 59392 163146 59394
rect 162485 59336 162490 59392
rect 162546 59336 163146 59392
rect 162485 59334 163146 59336
rect 163270 59392 164851 59394
rect 163270 59336 164790 59392
rect 164846 59336 164851 59392
rect 163270 59334 164851 59336
rect 155861 59331 155927 59334
rect 157609 59331 157675 59334
rect 158621 59331 158687 59334
rect 162485 59331 162551 59334
rect 148869 59256 150082 59258
rect 148869 59200 148874 59256
rect 148930 59200 150082 59256
rect 148869 59198 150082 59200
rect 162669 59258 162735 59261
rect 163270 59258 163330 59334
rect 164785 59331 164851 59334
rect 165245 59394 165311 59397
rect 167269 59394 167335 59397
rect 165245 59392 167335 59394
rect 165245 59336 165250 59392
rect 165306 59336 167274 59392
rect 167330 59336 167335 59392
rect 165245 59334 167335 59336
rect 165245 59331 165311 59334
rect 167269 59331 167335 59334
rect 168281 59394 168347 59397
rect 170416 59394 170476 60044
rect 171244 59530 171304 60044
rect 168281 59392 170476 59394
rect 168281 59336 168286 59392
rect 168342 59336 170476 59392
rect 168281 59334 170476 59336
rect 170630 59470 171304 59530
rect 171409 59530 171475 59533
rect 172072 59530 172132 60044
rect 171409 59528 172132 59530
rect 171409 59472 171414 59528
rect 171470 59472 172132 59528
rect 171409 59470 172132 59472
rect 168281 59331 168347 59334
rect 162669 59256 163330 59258
rect 162669 59200 162674 59256
rect 162730 59200 163330 59256
rect 162669 59198 163330 59200
rect 169569 59258 169635 59261
rect 170630 59258 170690 59470
rect 171409 59467 171475 59470
rect 170765 59394 170831 59397
rect 172900 59394 172960 60044
rect 173728 59938 173788 60044
rect 170765 59392 172960 59394
rect 170765 59336 170770 59392
rect 170826 59336 172960 59392
rect 170765 59334 172960 59336
rect 173206 59878 173788 59938
rect 170765 59331 170831 59334
rect 169569 59256 170690 59258
rect 169569 59200 169574 59256
rect 169630 59200 170690 59256
rect 169569 59198 170690 59200
rect 142061 59195 142127 59198
rect 148869 59195 148935 59198
rect 162669 59195 162735 59198
rect 169569 59195 169635 59198
rect 138841 59120 141066 59122
rect 138841 59064 138846 59120
rect 138902 59064 141066 59120
rect 138841 59062 141066 59064
rect 170949 59122 171015 59125
rect 173206 59122 173266 59878
rect 173341 59802 173407 59805
rect 174464 59802 174524 60044
rect 173341 59800 174524 59802
rect 173341 59744 173346 59800
rect 173402 59744 174524 59800
rect 173341 59742 174524 59744
rect 173341 59739 173407 59742
rect 173525 59666 173591 59669
rect 175292 59666 175352 60044
rect 173525 59664 175352 59666
rect 173525 59608 173530 59664
rect 173586 59608 175352 59664
rect 173525 59606 175352 59608
rect 175457 59666 175523 59669
rect 176120 59666 176180 60044
rect 175457 59664 176180 59666
rect 175457 59608 175462 59664
rect 175518 59608 176180 59664
rect 175457 59606 176180 59608
rect 173525 59603 173591 59606
rect 175457 59603 175523 59606
rect 175089 59530 175155 59533
rect 176948 59530 177008 60044
rect 177113 59666 177179 59669
rect 177776 59666 177836 60044
rect 177113 59664 177836 59666
rect 177113 59608 177118 59664
rect 177174 59608 177836 59664
rect 177113 59606 177836 59608
rect 177941 59666 178007 59669
rect 178604 59666 178664 60044
rect 177941 59664 178664 59666
rect 177941 59608 177946 59664
rect 178002 59608 178664 59664
rect 177941 59606 178664 59608
rect 177113 59603 177179 59606
rect 177941 59603 178007 59606
rect 175089 59528 177008 59530
rect 175089 59472 175094 59528
rect 175150 59472 177008 59528
rect 175089 59470 177008 59472
rect 177665 59530 177731 59533
rect 179432 59530 179492 60044
rect 177665 59528 179492 59530
rect 177665 59472 177670 59528
rect 177726 59472 179492 59528
rect 177665 59470 179492 59472
rect 175089 59467 175155 59470
rect 177665 59467 177731 59470
rect 173709 59394 173775 59397
rect 175457 59394 175523 59397
rect 173709 59392 175523 59394
rect 173709 59336 173714 59392
rect 173770 59336 175462 59392
rect 175518 59336 175523 59392
rect 173709 59334 175523 59336
rect 173709 59331 173775 59334
rect 175457 59331 175523 59334
rect 176561 59394 176627 59397
rect 177941 59394 178007 59397
rect 180260 59394 180320 60044
rect 180425 59530 180491 59533
rect 181088 59530 181148 60044
rect 180425 59528 181148 59530
rect 180425 59472 180430 59528
rect 180486 59472 181148 59528
rect 180425 59470 181148 59472
rect 180425 59467 180491 59470
rect 176561 59392 178007 59394
rect 176561 59336 176566 59392
rect 176622 59336 177946 59392
rect 178002 59336 178007 59392
rect 176561 59334 178007 59336
rect 176561 59331 176627 59334
rect 177941 59331 178007 59334
rect 178726 59334 180320 59394
rect 180701 59396 180767 59397
rect 180701 59392 180748 59396
rect 180812 59394 180818 59396
rect 181069 59394 181135 59397
rect 181916 59394 181976 60044
rect 182744 59394 182804 60044
rect 183572 59394 183632 60044
rect 183737 59802 183803 59805
rect 184400 59802 184460 60044
rect 183737 59800 184460 59802
rect 183737 59744 183742 59800
rect 183798 59744 184460 59800
rect 183737 59742 184460 59744
rect 183737 59739 183803 59742
rect 185228 59666 185288 60044
rect 185393 59802 185459 59805
rect 186056 59802 186116 60044
rect 185393 59800 186116 59802
rect 185393 59744 185398 59800
rect 185454 59744 186116 59800
rect 185393 59742 186116 59744
rect 186221 59802 186287 59805
rect 186884 59802 186944 60044
rect 186221 59800 186944 59802
rect 186221 59744 186226 59800
rect 186282 59744 186944 59800
rect 186221 59742 186944 59744
rect 185393 59739 185459 59742
rect 186221 59739 186287 59742
rect 180701 59336 180706 59392
rect 177849 59258 177915 59261
rect 178726 59258 178786 59334
rect 180701 59332 180748 59336
rect 180812 59334 180894 59394
rect 181069 59392 181976 59394
rect 181069 59336 181074 59392
rect 181130 59336 181976 59392
rect 181069 59334 181976 59336
rect 182038 59334 182804 59394
rect 182958 59334 183632 59394
rect 183694 59606 185288 59666
rect 185945 59666 186011 59669
rect 187712 59666 187772 60044
rect 185945 59664 187772 59666
rect 185945 59608 185950 59664
rect 186006 59608 187772 59664
rect 185945 59606 187772 59608
rect 187877 59666 187943 59669
rect 188540 59666 188600 60044
rect 187877 59664 188600 59666
rect 187877 59608 187882 59664
rect 187938 59608 188600 59664
rect 187877 59606 188600 59608
rect 180812 59332 180818 59334
rect 180701 59331 180767 59332
rect 181069 59331 181135 59334
rect 177849 59256 178786 59258
rect 177849 59200 177854 59256
rect 177910 59200 178786 59256
rect 177849 59198 178786 59200
rect 179137 59258 179203 59261
rect 180793 59258 180859 59261
rect 182038 59258 182098 59334
rect 179137 59256 180859 59258
rect 179137 59200 179142 59256
rect 179198 59200 180798 59256
rect 180854 59200 180859 59256
rect 179137 59198 180859 59200
rect 177849 59195 177915 59198
rect 179137 59195 179203 59198
rect 180793 59195 180859 59198
rect 181088 59198 182098 59258
rect 170949 59120 173266 59122
rect 170949 59064 170954 59120
rect 171010 59064 173266 59120
rect 170949 59062 173266 59064
rect 93853 59059 93919 59062
rect 138841 59059 138907 59062
rect 170949 59059 171015 59062
rect 180742 59060 180748 59124
rect 180812 59122 180818 59124
rect 181088 59122 181148 59198
rect 180812 59062 181148 59122
rect 181989 59122 182055 59125
rect 182958 59122 183018 59334
rect 183185 59258 183251 59261
rect 183694 59258 183754 59606
rect 185945 59603 186011 59606
rect 187877 59603 187943 59606
rect 184841 59530 184907 59533
rect 186221 59530 186287 59533
rect 184841 59528 186287 59530
rect 184841 59472 184846 59528
rect 184902 59472 186226 59528
rect 186282 59472 186287 59528
rect 184841 59470 186287 59472
rect 184841 59467 184907 59470
rect 186221 59467 186287 59470
rect 187325 59530 187391 59533
rect 189368 59530 189428 60044
rect 187325 59528 189428 59530
rect 187325 59472 187330 59528
rect 187386 59472 189428 59528
rect 187325 59470 189428 59472
rect 187325 59467 187391 59470
rect 185393 59394 185459 59397
rect 183185 59256 183754 59258
rect 183185 59200 183190 59256
rect 183246 59200 183754 59256
rect 183185 59198 183754 59200
rect 183878 59392 185459 59394
rect 183878 59336 185398 59392
rect 185454 59336 185459 59392
rect 183878 59334 185459 59336
rect 183185 59195 183251 59198
rect 181989 59120 183018 59122
rect 181989 59064 181994 59120
rect 182050 59064 183018 59120
rect 181989 59062 183018 59064
rect 183369 59122 183435 59125
rect 183878 59122 183938 59334
rect 185393 59331 185459 59334
rect 186129 59394 186195 59397
rect 187877 59394 187943 59397
rect 190104 59394 190164 60044
rect 190269 59530 190335 59533
rect 190932 59530 190992 60044
rect 190269 59528 190992 59530
rect 190269 59472 190274 59528
rect 190330 59472 190992 59528
rect 190269 59470 190992 59472
rect 190269 59467 190335 59470
rect 186129 59392 187943 59394
rect 186129 59336 186134 59392
rect 186190 59336 187882 59392
rect 187938 59336 187943 59392
rect 186129 59334 187943 59336
rect 186129 59331 186195 59334
rect 187877 59331 187943 59334
rect 188662 59334 190164 59394
rect 190545 59394 190611 59397
rect 191760 59394 191820 60044
rect 192588 59394 192648 60044
rect 193416 59394 193476 60044
rect 194244 59530 194304 60044
rect 194409 59802 194475 59805
rect 195072 59802 195132 60044
rect 195900 59938 195960 60044
rect 195286 59878 195960 59938
rect 195286 59805 195346 59878
rect 194409 59800 195132 59802
rect 194409 59744 194414 59800
rect 194470 59744 195132 59800
rect 194409 59742 195132 59744
rect 195237 59800 195346 59805
rect 196728 59802 196788 60044
rect 197556 59938 197616 60044
rect 195237 59744 195242 59800
rect 195298 59744 195346 59800
rect 195237 59742 195346 59744
rect 195470 59742 196788 59802
rect 196942 59878 197616 59938
rect 194409 59739 194475 59742
rect 195237 59739 195303 59742
rect 194501 59666 194567 59669
rect 194501 59664 194610 59666
rect 194501 59608 194506 59664
rect 194562 59608 194610 59664
rect 194501 59603 194610 59608
rect 194409 59530 194475 59533
rect 194244 59528 194475 59530
rect 194244 59472 194414 59528
rect 194470 59472 194475 59528
rect 194244 59470 194475 59472
rect 194550 59530 194610 59603
rect 195470 59530 195530 59742
rect 195789 59666 195855 59669
rect 196942 59666 197002 59878
rect 195789 59664 197002 59666
rect 195789 59608 195794 59664
rect 195850 59608 197002 59664
rect 195789 59606 197002 59608
rect 197077 59666 197143 59669
rect 198384 59666 198444 60044
rect 197077 59664 198444 59666
rect 197077 59608 197082 59664
rect 197138 59608 198444 59664
rect 197077 59606 198444 59608
rect 195789 59603 195855 59606
rect 197077 59603 197143 59606
rect 194550 59470 195530 59530
rect 197077 59530 197143 59533
rect 199212 59530 199272 60044
rect 200040 59802 200100 60044
rect 197077 59528 199272 59530
rect 197077 59472 197082 59528
rect 197138 59472 199272 59528
rect 197077 59470 199272 59472
rect 199334 59742 200100 59802
rect 194409 59467 194475 59470
rect 197077 59467 197143 59470
rect 195237 59394 195303 59397
rect 190545 59392 191820 59394
rect 190545 59336 190550 59392
rect 190606 59336 191820 59392
rect 190545 59334 191820 59336
rect 191974 59334 192648 59394
rect 192710 59334 193476 59394
rect 193630 59392 195303 59394
rect 193630 59336 195242 59392
rect 195298 59336 195303 59392
rect 193630 59334 195303 59336
rect 187509 59258 187575 59261
rect 188662 59258 188722 59334
rect 190545 59331 190611 59334
rect 187509 59256 188722 59258
rect 187509 59200 187514 59256
rect 187570 59200 188722 59256
rect 187509 59198 188722 59200
rect 190361 59258 190427 59261
rect 191974 59258 192034 59334
rect 190361 59256 192034 59258
rect 190361 59200 190366 59256
rect 190422 59200 192034 59256
rect 190361 59198 192034 59200
rect 187509 59195 187575 59198
rect 190361 59195 190427 59198
rect 183369 59120 183938 59122
rect 183369 59064 183374 59120
rect 183430 59064 183938 59120
rect 183369 59062 183938 59064
rect 191741 59122 191807 59125
rect 192710 59122 192770 59334
rect 193029 59258 193095 59261
rect 193630 59258 193690 59334
rect 195237 59331 195303 59334
rect 195605 59394 195671 59397
rect 196985 59394 197051 59397
rect 195605 59392 197051 59394
rect 195605 59336 195610 59392
rect 195666 59336 196990 59392
rect 197046 59336 197051 59392
rect 195605 59334 197051 59336
rect 195605 59331 195671 59334
rect 196985 59331 197051 59334
rect 197261 59394 197327 59397
rect 199334 59394 199394 59742
rect 200868 59666 200928 60044
rect 197261 59392 199394 59394
rect 197261 59336 197266 59392
rect 197322 59336 199394 59392
rect 197261 59334 199394 59336
rect 199518 59606 200928 59666
rect 201033 59666 201099 59669
rect 201696 59666 201756 60044
rect 201033 59664 201756 59666
rect 201033 59608 201038 59664
rect 201094 59608 201756 59664
rect 201033 59606 201756 59608
rect 197261 59331 197327 59334
rect 193029 59256 193690 59258
rect 193029 59200 193034 59256
rect 193090 59200 193690 59256
rect 193029 59198 193690 59200
rect 198641 59258 198707 59261
rect 199518 59258 199578 59606
rect 201033 59603 201099 59606
rect 200021 59530 200087 59533
rect 200205 59530 200271 59533
rect 202524 59530 202584 60044
rect 203352 59938 203412 60044
rect 204180 59938 204240 60044
rect 200021 59528 200130 59530
rect 200021 59472 200026 59528
rect 200082 59472 200130 59528
rect 200021 59467 200130 59472
rect 200205 59528 202584 59530
rect 200205 59472 200210 59528
rect 200266 59472 202584 59528
rect 200205 59470 202584 59472
rect 202646 59878 203412 59938
rect 203566 59878 204240 59938
rect 200205 59467 200271 59470
rect 200070 59394 200130 59467
rect 201033 59394 201099 59397
rect 200070 59392 201099 59394
rect 200070 59336 201038 59392
rect 201094 59336 201099 59392
rect 200070 59334 201099 59336
rect 201033 59331 201099 59334
rect 201217 59394 201283 59397
rect 202646 59394 202706 59878
rect 202781 59802 202847 59805
rect 203566 59802 203626 59878
rect 205008 59802 205068 60044
rect 202781 59800 203626 59802
rect 202781 59744 202786 59800
rect 202842 59744 203626 59800
rect 202781 59742 203626 59744
rect 203750 59742 205068 59802
rect 202781 59739 202847 59742
rect 202781 59530 202847 59533
rect 203750 59530 203810 59742
rect 204161 59666 204227 59669
rect 205836 59666 205896 60044
rect 204161 59664 205896 59666
rect 204161 59608 204166 59664
rect 204222 59608 205896 59664
rect 204161 59606 205896 59608
rect 206093 59666 206159 59669
rect 206572 59666 206632 60044
rect 206093 59664 206632 59666
rect 206093 59608 206098 59664
rect 206154 59608 206632 59664
rect 206093 59606 206632 59608
rect 204161 59603 204227 59606
rect 206093 59603 206159 59606
rect 202781 59528 203810 59530
rect 202781 59472 202786 59528
rect 202842 59472 203810 59528
rect 202781 59470 203810 59472
rect 205449 59530 205515 59533
rect 207400 59530 207460 60044
rect 205449 59528 207460 59530
rect 205449 59472 205454 59528
rect 205510 59472 207460 59528
rect 205449 59470 207460 59472
rect 207565 59530 207631 59533
rect 208228 59530 208288 60044
rect 207565 59528 208288 59530
rect 207565 59472 207570 59528
rect 207626 59472 208288 59528
rect 207565 59470 208288 59472
rect 202781 59467 202847 59470
rect 205449 59467 205515 59470
rect 207565 59467 207631 59470
rect 201217 59392 202706 59394
rect 201217 59336 201222 59392
rect 201278 59336 202706 59392
rect 201217 59334 202706 59336
rect 203977 59394 204043 59397
rect 206093 59394 206159 59397
rect 203977 59392 206159 59394
rect 203977 59336 203982 59392
rect 204038 59336 206098 59392
rect 206154 59336 206159 59392
rect 203977 59334 206159 59336
rect 201217 59331 201283 59334
rect 203977 59331 204043 59334
rect 206093 59331 206159 59334
rect 206921 59394 206987 59397
rect 209056 59394 209116 60044
rect 209884 59938 209944 60044
rect 210712 59938 210772 60044
rect 206921 59392 209116 59394
rect 206921 59336 206926 59392
rect 206982 59336 209116 59392
rect 206921 59334 209116 59336
rect 209270 59878 209944 59938
rect 210006 59878 210772 59938
rect 206921 59331 206987 59334
rect 198641 59256 199578 59258
rect 198641 59200 198646 59256
rect 198702 59200 199578 59256
rect 198641 59198 199578 59200
rect 208025 59258 208091 59261
rect 209270 59258 209330 59878
rect 209405 59802 209471 59805
rect 210006 59802 210066 59878
rect 211540 59802 211600 60044
rect 209405 59800 210066 59802
rect 209405 59744 209410 59800
rect 209466 59744 210066 59800
rect 209405 59742 210066 59744
rect 210926 59742 211600 59802
rect 211705 59802 211771 59805
rect 212368 59802 212428 60044
rect 211705 59800 212428 59802
rect 211705 59744 211710 59800
rect 211766 59744 212428 59800
rect 211705 59742 212428 59744
rect 209405 59739 209471 59742
rect 209405 59530 209471 59533
rect 210926 59530 210986 59742
rect 211705 59739 211771 59742
rect 211061 59666 211127 59669
rect 213196 59666 213256 60044
rect 211061 59664 213256 59666
rect 211061 59608 211066 59664
rect 211122 59608 213256 59664
rect 211061 59606 213256 59608
rect 211061 59603 211127 59606
rect 209405 59528 210986 59530
rect 209405 59472 209410 59528
rect 209466 59472 210986 59528
rect 209405 59470 210986 59472
rect 212349 59530 212415 59533
rect 214024 59530 214084 60044
rect 212349 59528 214084 59530
rect 212349 59472 212354 59528
rect 212410 59472 214084 59528
rect 212349 59470 214084 59472
rect 209405 59467 209471 59470
rect 212349 59467 212415 59470
rect 211705 59394 211771 59397
rect 210926 59392 211771 59394
rect 210926 59336 211710 59392
rect 211766 59336 211771 59392
rect 210926 59334 211771 59336
rect 208025 59256 209330 59258
rect 208025 59200 208030 59256
rect 208086 59200 209330 59256
rect 208025 59198 209330 59200
rect 209589 59258 209655 59261
rect 210926 59258 210986 59334
rect 211705 59331 211771 59334
rect 212165 59394 212231 59397
rect 214852 59394 214912 60044
rect 215680 59530 215740 60044
rect 215845 59802 215911 59805
rect 216508 59802 216568 60044
rect 215845 59800 216568 59802
rect 215845 59744 215850 59800
rect 215906 59744 216568 59800
rect 215845 59742 216568 59744
rect 215845 59739 215911 59742
rect 217336 59666 217396 60044
rect 212165 59392 214912 59394
rect 212165 59336 212170 59392
rect 212226 59336 214912 59392
rect 212165 59334 214912 59336
rect 214974 59470 215740 59530
rect 215894 59606 217396 59666
rect 212165 59331 212231 59334
rect 209589 59256 210986 59258
rect 209589 59200 209594 59256
rect 209650 59200 210986 59256
rect 209589 59198 210986 59200
rect 213729 59258 213795 59261
rect 214974 59258 215034 59470
rect 215201 59394 215267 59397
rect 215894 59394 215954 59606
rect 216489 59530 216555 59533
rect 218164 59530 218224 60044
rect 216489 59528 218224 59530
rect 216489 59472 216494 59528
rect 216550 59472 218224 59528
rect 216489 59470 218224 59472
rect 216489 59467 216555 59470
rect 215201 59392 215954 59394
rect 215201 59336 215206 59392
rect 215262 59336 215954 59392
rect 215201 59334 215954 59336
rect 216305 59394 216371 59397
rect 218992 59394 219052 60044
rect 219157 59666 219223 59669
rect 219820 59666 219880 60044
rect 219157 59664 219880 59666
rect 219157 59608 219162 59664
rect 219218 59608 219880 59664
rect 219157 59606 219880 59608
rect 219985 59666 220051 59669
rect 220648 59666 220708 60044
rect 219985 59664 220708 59666
rect 219985 59608 219990 59664
rect 220046 59608 220708 59664
rect 219985 59606 220708 59608
rect 219157 59603 219223 59606
rect 219985 59603 220051 59606
rect 219341 59530 219407 59533
rect 221476 59530 221536 60044
rect 222304 59938 222364 60044
rect 219341 59528 221536 59530
rect 219341 59472 219346 59528
rect 219402 59472 221536 59528
rect 219341 59470 221536 59472
rect 221598 59878 222364 59938
rect 219341 59467 219407 59470
rect 219985 59394 220051 59397
rect 221598 59394 221658 59878
rect 223040 59666 223100 60044
rect 223205 59802 223271 59805
rect 223868 59802 223928 60044
rect 224696 59938 224756 60044
rect 223205 59800 223928 59802
rect 223205 59744 223210 59800
rect 223266 59744 223928 59800
rect 223205 59742 223928 59744
rect 223990 59878 224756 59938
rect 223205 59739 223271 59742
rect 216305 59392 219052 59394
rect 216305 59336 216310 59392
rect 216366 59336 219052 59392
rect 216305 59334 219052 59336
rect 219206 59392 220051 59394
rect 219206 59336 219990 59392
rect 220046 59336 220051 59392
rect 219206 59334 220051 59336
rect 215201 59331 215267 59334
rect 216305 59331 216371 59334
rect 213729 59256 215034 59258
rect 213729 59200 213734 59256
rect 213790 59200 215034 59256
rect 213729 59198 215034 59200
rect 217869 59258 217935 59261
rect 219206 59258 219266 59334
rect 219985 59331 220051 59334
rect 220862 59334 221658 59394
rect 221782 59606 223100 59666
rect 217869 59256 219266 59258
rect 217869 59200 217874 59256
rect 217930 59200 219266 59256
rect 217869 59198 219266 59200
rect 220445 59258 220511 59261
rect 220862 59258 220922 59334
rect 220445 59256 220922 59258
rect 220445 59200 220450 59256
rect 220506 59200 220922 59256
rect 220445 59198 220922 59200
rect 193029 59195 193095 59198
rect 198641 59195 198707 59198
rect 208025 59195 208091 59198
rect 209589 59195 209655 59198
rect 213729 59195 213795 59198
rect 217869 59195 217935 59198
rect 220445 59195 220511 59198
rect 191741 59120 192770 59122
rect 191741 59064 191746 59120
rect 191802 59064 192770 59120
rect 191741 59062 192770 59064
rect 220629 59122 220695 59125
rect 221782 59122 221842 59606
rect 222009 59530 222075 59533
rect 223990 59530 224050 59878
rect 225524 59666 225584 60044
rect 224726 59606 225584 59666
rect 224726 59530 224786 59606
rect 222009 59528 224050 59530
rect 222009 59472 222014 59528
rect 222070 59472 224050 59528
rect 222009 59470 224050 59472
rect 224358 59470 224786 59530
rect 224861 59530 224927 59533
rect 226352 59530 226412 60044
rect 224861 59528 226412 59530
rect 224861 59472 224866 59528
rect 224922 59472 226412 59528
rect 224861 59470 226412 59472
rect 226517 59530 226583 59533
rect 227180 59530 227240 60044
rect 226517 59528 227240 59530
rect 226517 59472 226522 59528
rect 226578 59472 227240 59528
rect 226517 59470 227240 59472
rect 222009 59467 222075 59470
rect 221917 59394 221983 59397
rect 223205 59394 223271 59397
rect 221917 59392 223271 59394
rect 221917 59336 221922 59392
rect 221978 59336 223210 59392
rect 223266 59336 223271 59392
rect 221917 59334 223271 59336
rect 221917 59331 221983 59334
rect 223205 59331 223271 59334
rect 223481 59394 223547 59397
rect 224358 59394 224418 59470
rect 224861 59467 224927 59470
rect 226517 59467 226583 59470
rect 223481 59392 224418 59394
rect 223481 59336 223486 59392
rect 223542 59336 224418 59392
rect 223481 59334 224418 59336
rect 224769 59394 224835 59397
rect 225965 59394 226031 59397
rect 224769 59392 226031 59394
rect 224769 59336 224774 59392
rect 224830 59336 225970 59392
rect 226026 59336 226031 59392
rect 224769 59334 226031 59336
rect 223481 59331 223547 59334
rect 224769 59331 224835 59334
rect 225965 59331 226031 59334
rect 226149 59394 226215 59397
rect 228008 59394 228068 60044
rect 228836 59394 228896 60044
rect 229664 59938 229724 60044
rect 230492 59938 230552 60044
rect 229664 59878 229754 59938
rect 229001 59802 229067 59805
rect 229461 59802 229527 59805
rect 229001 59800 229527 59802
rect 229001 59744 229006 59800
rect 229062 59744 229466 59800
rect 229522 59744 229527 59800
rect 229001 59742 229527 59744
rect 229001 59739 229067 59742
rect 229461 59739 229527 59742
rect 229694 59700 229754 59878
rect 229001 59666 229067 59669
rect 229664 59666 229754 59700
rect 229001 59664 229754 59666
rect 229001 59608 229006 59664
rect 229062 59640 229754 59664
rect 229878 59878 230552 59938
rect 229062 59608 229724 59640
rect 229001 59606 229724 59608
rect 229001 59603 229067 59606
rect 229001 59530 229067 59533
rect 229878 59530 229938 59878
rect 230657 59802 230723 59805
rect 231320 59802 231380 60044
rect 232148 59938 232208 60044
rect 232976 59938 233036 60044
rect 230657 59800 231380 59802
rect 230657 59744 230662 59800
rect 230718 59744 231380 59800
rect 230657 59742 231380 59744
rect 231534 59878 232208 59938
rect 232270 59878 233036 59938
rect 230657 59739 230723 59742
rect 229001 59528 229938 59530
rect 229001 59472 229006 59528
rect 229062 59472 229938 59528
rect 229001 59470 229938 59472
rect 229001 59467 229067 59470
rect 226149 59392 228068 59394
rect 226149 59336 226154 59392
rect 226210 59336 228068 59392
rect 226149 59334 228068 59336
rect 228222 59334 228896 59394
rect 229921 59394 229987 59397
rect 231534 59394 231594 59878
rect 232270 59394 232330 59878
rect 233804 59802 233864 60044
rect 229921 59392 231594 59394
rect 229921 59336 229926 59392
rect 229982 59336 231594 59392
rect 229921 59334 231594 59336
rect 231718 59334 232330 59394
rect 232454 59742 233864 59802
rect 226149 59331 226215 59334
rect 225965 59258 226031 59261
rect 228222 59258 228282 59334
rect 229921 59331 229987 59334
rect 225965 59256 228282 59258
rect 225965 59200 225970 59256
rect 226026 59200 228282 59256
rect 225965 59198 228282 59200
rect 229737 59258 229803 59261
rect 231718 59258 231778 59334
rect 229737 59256 231778 59258
rect 229737 59200 229742 59256
rect 229798 59200 231778 59256
rect 229737 59198 231778 59200
rect 225965 59195 226031 59198
rect 229737 59195 229803 59198
rect 220629 59120 221842 59122
rect 220629 59064 220634 59120
rect 220690 59064 221842 59120
rect 220629 59062 221842 59064
rect 231117 59122 231183 59125
rect 232454 59122 232514 59742
rect 232681 59666 232747 59669
rect 234632 59666 234692 60044
rect 234797 59802 234863 59805
rect 235460 59802 235520 60044
rect 234797 59800 235520 59802
rect 234797 59744 234802 59800
rect 234858 59744 235520 59800
rect 234797 59742 235520 59744
rect 235625 59802 235691 59805
rect 236288 59802 236348 60044
rect 235625 59800 236348 59802
rect 235625 59744 235630 59800
rect 235686 59744 236348 59800
rect 235625 59742 236348 59744
rect 234797 59739 234863 59742
rect 235625 59739 235691 59742
rect 232681 59664 234692 59666
rect 232681 59608 232686 59664
rect 232742 59608 234692 59664
rect 232681 59606 234692 59608
rect 234797 59666 234863 59669
rect 237116 59666 237176 60044
rect 234797 59664 237176 59666
rect 234797 59608 234802 59664
rect 234858 59608 237176 59664
rect 234797 59606 237176 59608
rect 232681 59603 232747 59606
rect 234797 59603 234863 59606
rect 234061 59530 234127 59533
rect 235625 59530 235691 59533
rect 234061 59528 235691 59530
rect 234061 59472 234066 59528
rect 234122 59472 235630 59528
rect 235686 59472 235691 59528
rect 234061 59470 235691 59472
rect 234061 59467 234127 59470
rect 235625 59467 235691 59470
rect 233877 59394 233943 59397
rect 234797 59394 234863 59397
rect 233877 59392 234863 59394
rect 233877 59336 233882 59392
rect 233938 59336 234802 59392
rect 234858 59336 234863 59392
rect 233877 59334 234863 59336
rect 233877 59331 233943 59334
rect 234797 59331 234863 59334
rect 235441 59394 235507 59397
rect 237944 59394 238004 60044
rect 238680 59666 238740 60044
rect 238845 59802 238911 59805
rect 239508 59802 239568 60044
rect 238845 59800 239568 59802
rect 238845 59744 238850 59800
rect 238906 59744 239568 59800
rect 238845 59742 239568 59744
rect 238845 59739 238911 59742
rect 235441 59392 238004 59394
rect 235441 59336 235446 59392
rect 235502 59336 238004 59392
rect 235441 59334 238004 59336
rect 238158 59606 238740 59666
rect 235441 59331 235507 59334
rect 235257 59258 235323 59261
rect 238158 59258 238218 59606
rect 238293 59530 238359 59533
rect 240336 59530 240396 60044
rect 240501 59802 240567 59805
rect 241164 59802 241224 60044
rect 240501 59800 241224 59802
rect 240501 59744 240506 59800
rect 240562 59744 241224 59800
rect 240501 59742 241224 59744
rect 240501 59739 240567 59742
rect 238293 59528 240396 59530
rect 238293 59472 238298 59528
rect 238354 59472 240396 59528
rect 238293 59470 240396 59472
rect 238293 59467 238359 59470
rect 239581 59394 239647 59397
rect 241992 59394 242052 60044
rect 242157 59802 242223 59805
rect 242820 59802 242880 60044
rect 242157 59800 242880 59802
rect 242157 59744 242162 59800
rect 242218 59744 242880 59800
rect 242157 59742 242880 59744
rect 242157 59739 242223 59742
rect 243648 59666 243708 60044
rect 239581 59392 242052 59394
rect 239581 59336 239586 59392
rect 239642 59336 242052 59392
rect 239581 59334 242052 59336
rect 242206 59606 243708 59666
rect 239581 59331 239647 59334
rect 235257 59256 238218 59258
rect 235257 59200 235262 59256
rect 235318 59200 238218 59256
rect 235257 59198 238218 59200
rect 240777 59258 240843 59261
rect 242206 59258 242266 59606
rect 242341 59530 242407 59533
rect 244476 59530 244536 60044
rect 245304 59666 245364 60044
rect 245469 59802 245535 59805
rect 246132 59802 246192 60044
rect 245469 59800 246192 59802
rect 245469 59744 245474 59800
rect 245530 59744 246192 59800
rect 245469 59742 246192 59744
rect 245469 59739 245535 59742
rect 242341 59528 244536 59530
rect 242341 59472 242346 59528
rect 242402 59472 244536 59528
rect 242341 59470 244536 59472
rect 244598 59606 245364 59666
rect 245469 59666 245535 59669
rect 246960 59666 247020 60044
rect 245469 59664 247020 59666
rect 245469 59608 245474 59664
rect 245530 59608 247020 59664
rect 245469 59606 247020 59608
rect 242341 59467 242407 59470
rect 244598 59394 244658 59606
rect 245469 59603 245535 59606
rect 244917 59530 244983 59533
rect 247788 59530 247848 60044
rect 244917 59528 247848 59530
rect 244917 59472 244922 59528
rect 244978 59472 247848 59528
rect 244917 59470 247848 59472
rect 247953 59530 248019 59533
rect 248616 59530 248676 60044
rect 248873 59666 248939 59669
rect 249444 59666 249504 60044
rect 248873 59664 249504 59666
rect 248873 59608 248878 59664
rect 248934 59608 249504 59664
rect 248873 59606 249504 59608
rect 249609 59666 249675 59669
rect 250272 59666 250332 60044
rect 250529 59802 250595 59805
rect 251100 59802 251160 60044
rect 251928 59938 251988 60044
rect 252756 59938 252816 60044
rect 253584 59938 253644 60044
rect 251406 59878 251988 59938
rect 252142 59878 252816 59938
rect 252878 59878 253644 59938
rect 250529 59800 251160 59802
rect 250529 59744 250534 59800
rect 250590 59744 251160 59800
rect 250529 59742 251160 59744
rect 251265 59802 251331 59805
rect 251406 59802 251466 59878
rect 252142 59802 252202 59878
rect 251265 59800 251466 59802
rect 251265 59744 251270 59800
rect 251326 59744 251466 59800
rect 251265 59742 251466 59744
rect 251590 59742 252202 59802
rect 252277 59802 252343 59805
rect 252878 59802 252938 59878
rect 252277 59800 252938 59802
rect 252277 59744 252282 59800
rect 252338 59744 252938 59800
rect 252277 59742 252938 59744
rect 250529 59739 250595 59742
rect 251265 59739 251331 59742
rect 249609 59664 250332 59666
rect 249609 59608 249614 59664
rect 249670 59608 250332 59664
rect 249609 59606 250332 59608
rect 250621 59666 250687 59669
rect 251590 59666 251650 59742
rect 252277 59739 252343 59742
rect 250621 59664 251650 59666
rect 250621 59608 250626 59664
rect 250682 59608 251650 59664
rect 250621 59606 251650 59608
rect 248873 59603 248939 59606
rect 249609 59603 249675 59606
rect 250621 59603 250687 59606
rect 247953 59528 248676 59530
rect 247953 59472 247958 59528
rect 248014 59472 248676 59528
rect 247953 59470 248676 59472
rect 250437 59530 250503 59533
rect 252001 59530 252067 59533
rect 250437 59528 252067 59530
rect 250437 59472 250442 59528
rect 250498 59472 252006 59528
rect 252062 59472 252067 59528
rect 250437 59470 252067 59472
rect 244917 59467 244983 59470
rect 247953 59467 248019 59470
rect 250437 59467 250503 59470
rect 252001 59467 252067 59470
rect 252277 59530 252343 59533
rect 254412 59530 254472 60044
rect 254577 59802 254643 59805
rect 255148 59802 255208 60044
rect 254577 59800 255208 59802
rect 254577 59744 254582 59800
rect 254638 59744 255208 59800
rect 254577 59742 255208 59744
rect 254577 59739 254643 59742
rect 255976 59666 256036 60044
rect 252277 59528 254472 59530
rect 252277 59472 252282 59528
rect 252338 59472 254472 59528
rect 252277 59470 254472 59472
rect 254718 59606 256036 59666
rect 252277 59467 252343 59470
rect 245469 59394 245535 59397
rect 240777 59256 242266 59258
rect 240777 59200 240782 59256
rect 240838 59200 242266 59256
rect 240777 59198 242266 59200
rect 242390 59334 244658 59394
rect 244782 59392 245535 59394
rect 244782 59336 245474 59392
rect 245530 59336 245535 59392
rect 244782 59334 245535 59336
rect 235257 59195 235323 59198
rect 240777 59195 240843 59198
rect 231117 59120 232514 59122
rect 231117 59064 231122 59120
rect 231178 59064 232514 59120
rect 231117 59062 232514 59064
rect 242157 59122 242223 59125
rect 242390 59122 242450 59334
rect 243537 59258 243603 59261
rect 244782 59258 244842 59334
rect 245469 59331 245535 59334
rect 247677 59394 247743 59397
rect 249609 59394 249675 59397
rect 254577 59394 254643 59397
rect 247677 59392 249675 59394
rect 247677 59336 247682 59392
rect 247738 59336 249614 59392
rect 249670 59336 249675 59392
rect 247677 59334 249675 59336
rect 247677 59331 247743 59334
rect 249609 59331 249675 59334
rect 252878 59392 254643 59394
rect 252878 59336 254582 59392
rect 254638 59336 254643 59392
rect 252878 59334 254643 59336
rect 243537 59256 244842 59258
rect 243537 59200 243542 59256
rect 243598 59200 244842 59256
rect 243537 59198 244842 59200
rect 252461 59258 252527 59261
rect 252878 59258 252938 59334
rect 254577 59331 254643 59334
rect 252461 59256 252938 59258
rect 252461 59200 252466 59256
rect 252522 59200 252938 59256
rect 252461 59198 252938 59200
rect 253841 59258 253907 59261
rect 254718 59258 254778 59606
rect 255129 59530 255195 59533
rect 256804 59530 256864 60044
rect 255129 59528 256864 59530
rect 255129 59472 255134 59528
rect 255190 59472 256864 59528
rect 255129 59470 256864 59472
rect 255129 59467 255195 59470
rect 254945 59394 255011 59397
rect 257632 59394 257692 60044
rect 257797 59666 257863 59669
rect 258460 59666 258520 60044
rect 257797 59664 258520 59666
rect 257797 59608 257802 59664
rect 257858 59608 258520 59664
rect 257797 59606 258520 59608
rect 258625 59666 258691 59669
rect 259288 59666 259348 60044
rect 258625 59664 259348 59666
rect 258625 59608 258630 59664
rect 258686 59608 259348 59664
rect 258625 59606 259348 59608
rect 257797 59603 257863 59606
rect 258625 59603 258691 59606
rect 257981 59530 258047 59533
rect 260116 59530 260176 60044
rect 260944 59666 261004 60044
rect 257981 59528 260176 59530
rect 257981 59472 257986 59528
rect 258042 59472 260176 59528
rect 257981 59470 260176 59472
rect 260238 59606 261004 59666
rect 261109 59666 261175 59669
rect 261772 59666 261832 60044
rect 261109 59664 261832 59666
rect 261109 59608 261114 59664
rect 261170 59608 261832 59664
rect 261109 59606 261832 59608
rect 257981 59467 258047 59470
rect 258625 59394 258691 59397
rect 260238 59394 260298 59606
rect 261109 59603 261175 59606
rect 260741 59530 260807 59533
rect 262600 59530 262660 60044
rect 260741 59528 262660 59530
rect 260741 59472 260746 59528
rect 260802 59472 262660 59528
rect 260741 59470 262660 59472
rect 263428 59530 263488 60044
rect 264256 59530 264316 60044
rect 265084 59666 265144 60044
rect 265709 59666 265775 59669
rect 265084 59664 265775 59666
rect 265084 59608 265714 59664
rect 265770 59608 265775 59664
rect 265084 59606 265775 59608
rect 265912 59666 265972 60044
rect 266740 59802 266800 60044
rect 267568 59938 267628 60044
rect 267568 59878 267658 59938
rect 267457 59802 267523 59805
rect 266740 59800 267523 59802
rect 266740 59744 267462 59800
rect 267518 59744 267523 59800
rect 266740 59742 267523 59744
rect 267457 59739 267523 59742
rect 267598 59666 267658 59878
rect 265912 59606 267474 59666
rect 265709 59603 265775 59606
rect 266997 59530 267063 59533
rect 263428 59470 263610 59530
rect 264256 59528 267063 59530
rect 264256 59472 267002 59528
rect 267058 59472 267063 59528
rect 264256 59470 267063 59472
rect 260741 59467 260807 59470
rect 254945 59392 257692 59394
rect 254945 59336 254950 59392
rect 255006 59336 257692 59392
rect 254945 59334 257692 59336
rect 257846 59392 258691 59394
rect 257846 59336 258630 59392
rect 258686 59336 258691 59392
rect 257846 59334 258691 59336
rect 254945 59331 255011 59334
rect 253841 59256 254778 59258
rect 253841 59200 253846 59256
rect 253902 59200 254778 59256
rect 253841 59198 254778 59200
rect 256509 59258 256575 59261
rect 257846 59258 257906 59334
rect 258625 59331 258691 59334
rect 259502 59334 260298 59394
rect 263550 59394 263610 59470
rect 266997 59467 267063 59470
rect 265525 59394 265591 59397
rect 263550 59392 265591 59394
rect 263550 59336 265530 59392
rect 265586 59336 265591 59392
rect 263550 59334 265591 59336
rect 256509 59256 257906 59258
rect 256509 59200 256514 59256
rect 256570 59200 257906 59256
rect 256509 59198 257906 59200
rect 259269 59258 259335 59261
rect 259502 59258 259562 59334
rect 265525 59331 265591 59334
rect 265709 59394 265775 59397
rect 267414 59394 267474 59606
rect 267568 59606 267658 59666
rect 268396 59666 268456 60044
rect 269224 59802 269284 60044
rect 269849 59802 269915 59805
rect 269224 59800 269915 59802
rect 269224 59744 269854 59800
rect 269910 59744 269915 59800
rect 269224 59742 269915 59744
rect 270052 59802 270112 60044
rect 270677 59802 270743 59805
rect 270052 59800 270743 59802
rect 270052 59744 270682 59800
rect 270738 59744 270743 59800
rect 270052 59742 270743 59744
rect 269849 59739 269915 59742
rect 270677 59739 270743 59742
rect 270677 59666 270743 59669
rect 268396 59664 270743 59666
rect 268396 59608 270682 59664
rect 270738 59608 270743 59664
rect 268396 59606 270743 59608
rect 267568 59530 267628 59606
rect 270677 59603 270743 59606
rect 269757 59530 269823 59533
rect 267568 59528 269823 59530
rect 267568 59472 269762 59528
rect 269818 59472 269823 59528
rect 267568 59470 269823 59472
rect 269757 59467 269823 59470
rect 268561 59394 268627 59397
rect 265709 59392 267290 59394
rect 265709 59336 265714 59392
rect 265770 59336 267290 59392
rect 265709 59334 267290 59336
rect 267414 59392 268627 59394
rect 267414 59336 268566 59392
rect 268622 59336 268627 59392
rect 267414 59334 268627 59336
rect 270880 59394 270940 60044
rect 271616 59530 271676 60044
rect 272241 59530 272307 59533
rect 271616 59528 272307 59530
rect 271616 59472 272246 59528
rect 272302 59472 272307 59528
rect 271616 59470 272307 59472
rect 272241 59467 272307 59470
rect 272444 59394 272504 60044
rect 273272 59530 273332 60044
rect 273897 59530 273963 59533
rect 273272 59528 273963 59530
rect 273272 59472 273902 59528
rect 273958 59472 273963 59528
rect 273272 59470 273963 59472
rect 273897 59467 273963 59470
rect 274100 59394 274160 60044
rect 274928 59530 274988 60044
rect 275756 59666 275816 60044
rect 276381 59666 276447 59669
rect 275756 59664 276447 59666
rect 275756 59608 276386 59664
rect 276442 59608 276447 59664
rect 275756 59606 276447 59608
rect 276584 59666 276644 60044
rect 277412 59802 277472 60044
rect 278037 59802 278103 59805
rect 277412 59800 278103 59802
rect 277412 59744 278042 59800
rect 278098 59744 278103 59800
rect 277412 59742 278103 59744
rect 278240 59802 278300 60044
rect 278865 59802 278931 59805
rect 278240 59800 278931 59802
rect 278240 59744 278870 59800
rect 278926 59744 278931 59800
rect 278240 59742 278931 59744
rect 279068 59802 279128 60044
rect 279896 59938 279956 60044
rect 279896 59878 280538 59938
rect 279068 59742 279802 59802
rect 278037 59739 278103 59742
rect 278865 59739 278931 59742
rect 279417 59666 279483 59669
rect 276584 59606 277410 59666
rect 276381 59603 276447 59606
rect 277209 59530 277275 59533
rect 274928 59528 277275 59530
rect 274928 59472 277214 59528
rect 277270 59472 277275 59528
rect 274928 59470 277275 59472
rect 277350 59530 277410 59606
rect 277534 59664 279483 59666
rect 277534 59608 279422 59664
rect 279478 59608 279483 59664
rect 277534 59606 279483 59608
rect 279742 59666 279802 59742
rect 280337 59666 280403 59669
rect 279742 59664 280403 59666
rect 279742 59608 280342 59664
rect 280398 59608 280403 59664
rect 279742 59606 280403 59608
rect 280478 59666 280538 59878
rect 280724 59802 280784 60044
rect 281552 59938 281612 60044
rect 281552 59878 281642 59938
rect 281349 59802 281415 59805
rect 280724 59800 281415 59802
rect 280724 59744 281354 59800
rect 281410 59744 281415 59800
rect 280724 59742 281415 59744
rect 281349 59739 281415 59742
rect 281582 59666 281642 59878
rect 282380 59802 282440 60044
rect 283005 59802 283071 59805
rect 282380 59800 283071 59802
rect 282380 59744 283010 59800
rect 283066 59744 283071 59800
rect 282380 59742 283071 59744
rect 283005 59739 283071 59742
rect 280478 59606 281458 59666
rect 277534 59530 277594 59606
rect 279417 59603 279483 59606
rect 280337 59603 280403 59606
rect 277350 59470 277594 59530
rect 278037 59530 278103 59533
rect 278865 59530 278931 59533
rect 280797 59530 280863 59533
rect 278037 59528 278698 59530
rect 278037 59472 278042 59528
rect 278098 59472 278698 59528
rect 278037 59470 278698 59472
rect 277209 59467 277275 59470
rect 278037 59467 278103 59470
rect 276381 59394 276447 59397
rect 277945 59394 278011 59397
rect 270880 59334 272258 59394
rect 272444 59334 273914 59394
rect 274100 59334 276306 59394
rect 265709 59331 265775 59334
rect 259269 59256 259562 59258
rect 259269 59200 259274 59256
rect 259330 59200 259562 59256
rect 259269 59198 259562 59200
rect 267230 59258 267290 59334
rect 268561 59331 268627 59334
rect 268377 59258 268443 59261
rect 267230 59256 268443 59258
rect 267230 59200 268382 59256
rect 268438 59200 268443 59256
rect 267230 59198 268443 59200
rect 272198 59258 272258 59334
rect 273713 59258 273779 59261
rect 272198 59256 273779 59258
rect 272198 59200 273718 59256
rect 273774 59200 273779 59256
rect 272198 59198 273779 59200
rect 273854 59258 273914 59334
rect 274633 59258 274699 59261
rect 273854 59256 274699 59258
rect 273854 59200 274638 59256
rect 274694 59200 274699 59256
rect 273854 59198 274699 59200
rect 276246 59258 276306 59334
rect 276381 59392 278011 59394
rect 276381 59336 276386 59392
rect 276442 59336 277950 59392
rect 278006 59336 278011 59392
rect 276381 59334 278011 59336
rect 278638 59394 278698 59470
rect 278865 59528 280863 59530
rect 278865 59472 278870 59528
rect 278926 59472 280802 59528
rect 280858 59472 280863 59528
rect 278865 59470 280863 59472
rect 278865 59467 278931 59470
rect 280797 59467 280863 59470
rect 280981 59394 281047 59397
rect 278638 59392 281047 59394
rect 278638 59336 280986 59392
rect 281042 59336 281047 59392
rect 278638 59334 281047 59336
rect 276381 59331 276447 59334
rect 277945 59331 278011 59334
rect 280981 59331 281047 59334
rect 276841 59258 276907 59261
rect 276246 59256 276907 59258
rect 276246 59200 276846 59256
rect 276902 59200 276907 59256
rect 276246 59198 276907 59200
rect 281398 59258 281458 59606
rect 281552 59606 281642 59666
rect 281552 59394 281612 59606
rect 281717 59530 281783 59533
rect 283005 59530 283071 59533
rect 281717 59528 283071 59530
rect 281717 59472 281722 59528
rect 281778 59472 283010 59528
rect 283066 59472 283071 59528
rect 281717 59470 283071 59472
rect 281717 59467 281783 59470
rect 283005 59467 283071 59470
rect 283208 59394 283268 60044
rect 284036 59530 284096 60044
rect 284864 59666 284924 60044
rect 285692 59802 285752 60044
rect 286317 59802 286383 59805
rect 285692 59800 286383 59802
rect 285692 59744 286322 59800
rect 286378 59744 286383 59800
rect 285692 59742 286383 59744
rect 286520 59802 286580 60044
rect 287145 59802 287211 59805
rect 286520 59800 287211 59802
rect 286520 59744 287150 59800
rect 287206 59744 287211 59800
rect 286520 59742 287211 59744
rect 287348 59802 287408 60044
rect 287881 59802 287947 59805
rect 287348 59800 287947 59802
rect 287348 59744 287886 59800
rect 287942 59744 287947 59800
rect 287348 59742 287947 59744
rect 286317 59739 286383 59742
rect 287145 59739 287211 59742
rect 287881 59739 287947 59742
rect 287697 59666 287763 59669
rect 284864 59664 287763 59666
rect 284864 59608 287702 59664
rect 287758 59608 287763 59664
rect 284864 59606 287763 59608
rect 287697 59603 287763 59606
rect 286317 59530 286383 59533
rect 284036 59528 286383 59530
rect 284036 59472 286322 59528
rect 286378 59472 286383 59528
rect 284036 59470 286383 59472
rect 288084 59530 288144 60044
rect 288912 59666 288972 60044
rect 289537 59666 289603 59669
rect 288912 59664 289603 59666
rect 288912 59608 289542 59664
rect 289598 59608 289603 59664
rect 288912 59606 289603 59608
rect 289740 59666 289800 60044
rect 290568 59802 290628 60044
rect 291396 59938 291456 60044
rect 292224 59938 292284 60044
rect 293052 59938 293112 60044
rect 291396 59878 291946 59938
rect 292224 59878 292866 59938
rect 293052 59878 293602 59938
rect 291745 59802 291811 59805
rect 291886 59804 291946 59878
rect 290568 59800 291811 59802
rect 290568 59744 291750 59800
rect 291806 59744 291811 59800
rect 290568 59742 291811 59744
rect 291745 59739 291811 59742
rect 291878 59740 291884 59804
rect 291948 59740 291954 59804
rect 292806 59802 292866 59878
rect 293401 59802 293467 59805
rect 292806 59800 293467 59802
rect 292806 59744 293406 59800
rect 293462 59744 293467 59800
rect 292806 59742 293467 59744
rect 293542 59802 293602 59878
rect 293677 59802 293743 59805
rect 293542 59800 293743 59802
rect 293542 59744 293682 59800
rect 293738 59744 293743 59800
rect 293542 59742 293743 59744
rect 293880 59802 293940 60044
rect 294413 59802 294479 59805
rect 293880 59800 294479 59802
rect 293880 59744 294418 59800
rect 294474 59744 294479 59800
rect 293880 59742 294479 59744
rect 293401 59739 293467 59742
rect 293677 59739 293743 59742
rect 294413 59739 294479 59742
rect 292021 59666 292087 59669
rect 289740 59664 292087 59666
rect 289740 59608 292026 59664
rect 292082 59608 292087 59664
rect 289740 59606 292087 59608
rect 289537 59603 289603 59606
rect 292021 59603 292087 59606
rect 290457 59530 290523 59533
rect 288084 59528 290523 59530
rect 288084 59472 290462 59528
rect 290518 59472 290523 59528
rect 288084 59470 290523 59472
rect 294708 59530 294768 60044
rect 295536 59666 295596 60044
rect 296364 59802 296424 60044
rect 296989 59802 297055 59805
rect 296364 59800 297055 59802
rect 296364 59744 296994 59800
rect 297050 59744 297055 59800
rect 296364 59742 297055 59744
rect 296989 59739 297055 59742
rect 296529 59666 296595 59669
rect 295536 59664 296595 59666
rect 295536 59608 296534 59664
rect 296590 59608 296595 59664
rect 295536 59606 296595 59608
rect 296529 59603 296595 59606
rect 296989 59530 297055 59533
rect 294708 59528 297055 59530
rect 294708 59472 296994 59528
rect 297050 59472 297055 59528
rect 294708 59470 297055 59472
rect 286317 59467 286383 59470
rect 290457 59467 290523 59470
rect 296989 59467 297055 59470
rect 287145 59394 287211 59397
rect 289077 59394 289143 59397
rect 281552 59334 283114 59394
rect 283208 59334 286426 59394
rect 282361 59258 282427 59261
rect 281398 59256 282427 59258
rect 281398 59200 282366 59256
rect 282422 59200 282427 59256
rect 281398 59198 282427 59200
rect 283054 59258 283114 59334
rect 284937 59258 285003 59261
rect 283054 59256 285003 59258
rect 283054 59200 284942 59256
rect 284998 59200 285003 59256
rect 283054 59198 285003 59200
rect 286366 59258 286426 59334
rect 287145 59392 289143 59394
rect 287145 59336 287150 59392
rect 287206 59336 289082 59392
rect 289138 59336 289143 59392
rect 287145 59334 289143 59336
rect 287145 59331 287211 59334
rect 289077 59331 289143 59334
rect 289537 59394 289603 59397
rect 291837 59394 291903 59397
rect 289537 59392 291903 59394
rect 289537 59336 289542 59392
rect 289598 59336 291842 59392
rect 291898 59336 291903 59392
rect 289537 59334 291903 59336
rect 289537 59331 289603 59334
rect 291837 59331 291903 59334
rect 294413 59394 294479 59397
rect 296161 59394 296227 59397
rect 294413 59392 296227 59394
rect 294413 59336 294418 59392
rect 294474 59336 296166 59392
rect 296222 59336 296227 59392
rect 294413 59334 296227 59336
rect 297192 59394 297252 60044
rect 298020 59530 298080 60044
rect 298848 59666 298908 60044
rect 299676 59802 299736 60044
rect 300301 59802 300367 59805
rect 299676 59800 300367 59802
rect 299676 59744 300306 59800
rect 300362 59744 300367 59800
rect 299676 59742 300367 59744
rect 300504 59802 300564 60044
rect 301129 59802 301195 59805
rect 300504 59800 301195 59802
rect 300504 59744 301134 59800
rect 301190 59744 301195 59800
rect 300504 59742 301195 59744
rect 301332 59802 301392 60044
rect 301957 59802 302023 59805
rect 301332 59800 302023 59802
rect 301332 59744 301962 59800
rect 302018 59744 302023 59800
rect 301332 59742 302023 59744
rect 300301 59739 300367 59742
rect 301129 59739 301195 59742
rect 301957 59739 302023 59742
rect 301497 59666 301563 59669
rect 298848 59664 301563 59666
rect 298848 59608 301502 59664
rect 301558 59608 301563 59664
rect 298848 59606 301563 59608
rect 301497 59603 301563 59606
rect 300117 59530 300183 59533
rect 298020 59528 300183 59530
rect 298020 59472 300122 59528
rect 300178 59472 300183 59528
rect 298020 59470 300183 59472
rect 300117 59467 300183 59470
rect 300301 59394 300367 59397
rect 297192 59392 300367 59394
rect 297192 59336 300306 59392
rect 300362 59336 300367 59392
rect 297192 59334 300367 59336
rect 294413 59331 294479 59334
rect 296161 59331 296227 59334
rect 300301 59331 300367 59334
rect 301129 59394 301195 59397
rect 302160 59394 302220 60044
rect 302988 59530 303048 60044
rect 303724 59666 303784 60044
rect 304349 59666 304415 59669
rect 303724 59664 304415 59666
rect 303724 59608 304354 59664
rect 304410 59608 304415 59664
rect 303724 59606 304415 59608
rect 304552 59666 304612 60044
rect 305380 59802 305440 60044
rect 305913 59802 305979 59805
rect 305380 59800 305979 59802
rect 305380 59744 305918 59800
rect 305974 59744 305979 59800
rect 305380 59742 305979 59744
rect 305913 59739 305979 59742
rect 306005 59666 306071 59669
rect 304552 59664 306071 59666
rect 304552 59608 306010 59664
rect 306066 59608 306071 59664
rect 304552 59606 306071 59608
rect 304349 59603 304415 59606
rect 306005 59603 306071 59606
rect 305637 59530 305703 59533
rect 302988 59470 303722 59530
rect 303662 59394 303722 59470
rect 304214 59528 305703 59530
rect 304214 59472 305642 59528
rect 305698 59472 305703 59528
rect 304214 59470 305703 59472
rect 304214 59394 304274 59470
rect 305637 59467 305703 59470
rect 301129 59392 302066 59394
rect 301129 59336 301134 59392
rect 301190 59336 302066 59392
rect 301129 59334 302066 59336
rect 302160 59334 303538 59394
rect 303662 59334 304274 59394
rect 304349 59394 304415 59397
rect 306208 59394 306268 60044
rect 306833 59394 306899 59397
rect 304349 59392 306114 59394
rect 304349 59336 304354 59392
rect 304410 59336 306114 59392
rect 304349 59334 306114 59336
rect 306208 59392 306899 59394
rect 306208 59336 306838 59392
rect 306894 59336 306899 59392
rect 306208 59334 306899 59336
rect 307036 59394 307096 60044
rect 307864 59530 307924 60044
rect 308489 59530 308555 59533
rect 307864 59528 308555 59530
rect 307864 59472 308494 59528
rect 308550 59472 308555 59528
rect 307864 59470 308555 59472
rect 308489 59467 308555 59470
rect 308692 59394 308752 60044
rect 309520 59666 309580 60044
rect 310145 59666 310211 59669
rect 309520 59664 310211 59666
rect 309520 59608 310150 59664
rect 310206 59608 310211 59664
rect 309520 59606 310211 59608
rect 310145 59603 310211 59606
rect 310348 59530 310408 60044
rect 311176 59666 311236 60044
rect 312004 59802 312064 60044
rect 312629 59802 312695 59805
rect 312004 59800 312695 59802
rect 312004 59744 312634 59800
rect 312690 59744 312695 59800
rect 312004 59742 312695 59744
rect 312629 59739 312695 59742
rect 312537 59666 312603 59669
rect 311176 59664 312603 59666
rect 311176 59608 312542 59664
rect 312598 59608 312603 59664
rect 311176 59606 312603 59608
rect 312537 59603 312603 59606
rect 312537 59530 312603 59533
rect 310348 59528 312603 59530
rect 310348 59472 312542 59528
rect 312598 59472 312603 59528
rect 310348 59470 312603 59472
rect 312832 59530 312892 60044
rect 313660 59802 313720 60044
rect 314285 59802 314351 59805
rect 313660 59800 314351 59802
rect 313660 59744 314290 59800
rect 314346 59744 314351 59800
rect 313660 59742 314351 59744
rect 314285 59739 314351 59742
rect 314285 59530 314351 59533
rect 312832 59528 314351 59530
rect 312832 59472 314290 59528
rect 314346 59472 314351 59528
rect 312832 59470 314351 59472
rect 312537 59467 312603 59470
rect 314285 59467 314351 59470
rect 311341 59394 311407 59397
rect 307036 59334 308506 59394
rect 308692 59392 311407 59394
rect 308692 59336 311346 59392
rect 311402 59336 311407 59392
rect 308692 59334 311407 59336
rect 301129 59331 301195 59334
rect 286501 59258 286567 59261
rect 286366 59256 286567 59258
rect 286366 59200 286506 59256
rect 286562 59200 286567 59256
rect 286366 59198 286567 59200
rect 302006 59258 302066 59334
rect 303061 59258 303127 59261
rect 302006 59256 303127 59258
rect 302006 59200 303066 59256
rect 303122 59200 303127 59256
rect 302006 59198 303127 59200
rect 303478 59258 303538 59334
rect 304349 59331 304415 59334
rect 304441 59258 304507 59261
rect 303478 59256 304507 59258
rect 303478 59200 304446 59256
rect 304502 59200 304507 59256
rect 303478 59198 304507 59200
rect 306054 59258 306114 59334
rect 306833 59331 306899 59334
rect 307017 59258 307083 59261
rect 306054 59256 307083 59258
rect 306054 59200 307022 59256
rect 307078 59200 307083 59256
rect 306054 59198 307083 59200
rect 308446 59258 308506 59334
rect 311341 59331 311407 59334
rect 312629 59394 312695 59397
rect 314488 59394 314548 60044
rect 315316 59530 315376 60044
rect 316144 59802 316204 60044
rect 316972 59805 317032 60044
rect 316769 59802 316835 59805
rect 316144 59800 316835 59802
rect 316144 59744 316774 59800
rect 316830 59744 316835 59800
rect 316144 59742 316835 59744
rect 316769 59739 316835 59742
rect 316953 59800 317032 59805
rect 316953 59744 316958 59800
rect 317014 59744 317032 59800
rect 316953 59742 317032 59744
rect 316953 59739 317019 59742
rect 317413 59666 317479 59669
rect 315990 59664 317479 59666
rect 315990 59608 317418 59664
rect 317474 59608 317479 59664
rect 315990 59606 317479 59608
rect 315990 59530 316050 59606
rect 317413 59603 317479 59606
rect 315316 59470 316050 59530
rect 316769 59394 316835 59397
rect 317800 59394 317860 60044
rect 318628 59530 318688 60044
rect 319456 59666 319516 60044
rect 320192 59802 320252 60044
rect 320817 59802 320883 59805
rect 320192 59800 320883 59802
rect 320192 59744 320822 59800
rect 320878 59744 320883 59800
rect 320192 59742 320883 59744
rect 320817 59739 320883 59742
rect 319456 59606 320834 59666
rect 320357 59530 320423 59533
rect 318628 59528 320423 59530
rect 318628 59472 320362 59528
rect 320418 59472 320423 59528
rect 318628 59470 320423 59472
rect 320357 59467 320423 59470
rect 320541 59394 320607 59397
rect 312629 59392 314394 59394
rect 312629 59336 312634 59392
rect 312690 59336 314394 59392
rect 312629 59334 314394 59336
rect 314488 59334 316050 59394
rect 312629 59331 312695 59334
rect 309777 59258 309843 59261
rect 308446 59256 309843 59258
rect 308446 59200 309782 59256
rect 309838 59200 309843 59256
rect 308446 59198 309843 59200
rect 314334 59258 314394 59334
rect 315297 59258 315363 59261
rect 314334 59256 315363 59258
rect 314334 59200 315302 59256
rect 315358 59200 315363 59256
rect 314334 59198 315363 59200
rect 315990 59258 316050 59334
rect 316769 59392 317706 59394
rect 316769 59336 316774 59392
rect 316830 59336 317706 59392
rect 316769 59334 317706 59336
rect 317800 59392 320607 59394
rect 317800 59336 320546 59392
rect 320602 59336 320607 59392
rect 317800 59334 320607 59336
rect 320774 59394 320834 59606
rect 321020 59530 321080 60044
rect 321848 59666 321908 60044
rect 322473 59666 322539 59669
rect 321848 59664 322539 59666
rect 321848 59608 322478 59664
rect 322534 59608 322539 59664
rect 321848 59606 322539 59608
rect 322676 59666 322736 60044
rect 323504 59802 323564 60044
rect 324129 59802 324195 59805
rect 323504 59800 324195 59802
rect 323504 59744 324134 59800
rect 324190 59744 324195 59800
rect 323504 59742 324195 59744
rect 324332 59802 324392 60044
rect 324957 59802 325023 59805
rect 324332 59800 325023 59802
rect 324332 59744 324962 59800
rect 325018 59744 325023 59800
rect 324332 59742 325023 59744
rect 324129 59739 324195 59742
rect 324957 59739 325023 59742
rect 324773 59666 324839 59669
rect 322676 59664 324839 59666
rect 322676 59608 324778 59664
rect 324834 59608 324839 59664
rect 322676 59606 324839 59608
rect 322473 59603 322539 59606
rect 324773 59603 324839 59606
rect 323301 59530 323367 59533
rect 321020 59528 323367 59530
rect 321020 59472 323306 59528
rect 323362 59472 323367 59528
rect 321020 59470 323367 59472
rect 323301 59467 323367 59470
rect 321645 59394 321711 59397
rect 320774 59392 321711 59394
rect 320774 59336 321650 59392
rect 321706 59336 321711 59392
rect 320774 59334 321711 59336
rect 316769 59331 316835 59334
rect 316861 59258 316927 59261
rect 315990 59256 316927 59258
rect 315990 59200 316866 59256
rect 316922 59200 316927 59256
rect 315990 59198 316927 59200
rect 317646 59258 317706 59334
rect 320541 59331 320607 59334
rect 321645 59331 321711 59334
rect 322473 59394 322539 59397
rect 324129 59394 324195 59397
rect 325160 59394 325220 60044
rect 325785 59394 325851 59397
rect 322473 59392 323410 59394
rect 322473 59336 322478 59392
rect 322534 59336 323410 59392
rect 322473 59334 323410 59336
rect 322473 59331 322539 59334
rect 318885 59258 318951 59261
rect 317646 59256 318951 59258
rect 317646 59200 318890 59256
rect 318946 59200 318951 59256
rect 317646 59198 318951 59200
rect 323350 59258 323410 59334
rect 324129 59392 325066 59394
rect 324129 59336 324134 59392
rect 324190 59336 325066 59392
rect 324129 59334 325066 59336
rect 325160 59392 325851 59394
rect 325160 59336 325790 59392
rect 325846 59336 325851 59392
rect 325160 59334 325851 59336
rect 325988 59394 326048 60044
rect 326816 59394 326876 60044
rect 327644 59394 327704 60044
rect 328472 59530 328532 60044
rect 329097 59530 329163 59533
rect 328472 59528 329163 59530
rect 328472 59472 329102 59528
rect 329158 59472 329163 59528
rect 328472 59470 329163 59472
rect 329300 59530 329360 60044
rect 330128 59666 330188 60044
rect 330293 59802 330359 59805
rect 330956 59802 331016 60044
rect 330293 59800 331016 59802
rect 330293 59744 330298 59800
rect 330354 59744 331016 59800
rect 330293 59742 331016 59744
rect 330293 59739 330359 59742
rect 330128 59606 331690 59666
rect 331489 59530 331555 59533
rect 329300 59528 331555 59530
rect 329300 59472 331494 59528
rect 331550 59472 331555 59528
rect 329300 59470 331555 59472
rect 329097 59467 329163 59470
rect 331489 59467 331555 59470
rect 329925 59394 329991 59397
rect 325988 59334 326722 59394
rect 326816 59334 327458 59394
rect 327644 59392 329991 59394
rect 327644 59336 329930 59392
rect 329986 59336 329991 59392
rect 327644 59334 329991 59336
rect 331630 59394 331690 59606
rect 331784 59530 331844 60044
rect 332612 59666 332672 60044
rect 333237 59666 333303 59669
rect 332612 59664 333303 59666
rect 332612 59608 333242 59664
rect 333298 59608 333303 59664
rect 332612 59606 333303 59608
rect 333440 59666 333500 60044
rect 334268 59802 334328 60044
rect 334893 59802 334959 59805
rect 334268 59800 334959 59802
rect 334268 59744 334898 59800
rect 334954 59744 334959 59800
rect 334268 59742 334959 59744
rect 334893 59739 334959 59742
rect 333440 59606 335002 59666
rect 333237 59603 333303 59606
rect 334065 59530 334131 59533
rect 331784 59528 334131 59530
rect 331784 59472 334070 59528
rect 334126 59472 334131 59528
rect 331784 59470 334131 59472
rect 334065 59467 334131 59470
rect 332685 59394 332751 59397
rect 331630 59392 332751 59394
rect 331630 59336 332690 59392
rect 332746 59336 332751 59392
rect 331630 59334 332751 59336
rect 324129 59331 324195 59334
rect 324589 59258 324655 59261
rect 323350 59256 324655 59258
rect 323350 59200 324594 59256
rect 324650 59200 324655 59256
rect 323350 59198 324655 59200
rect 325006 59258 325066 59334
rect 325785 59331 325851 59334
rect 325693 59258 325759 59261
rect 325006 59256 325759 59258
rect 325006 59200 325698 59256
rect 325754 59200 325759 59256
rect 325006 59198 325759 59200
rect 243537 59195 243603 59198
rect 252461 59195 252527 59198
rect 253841 59195 253907 59198
rect 256509 59195 256575 59198
rect 259269 59195 259335 59198
rect 268377 59195 268443 59198
rect 273713 59195 273779 59198
rect 274633 59195 274699 59198
rect 276841 59195 276907 59198
rect 282361 59195 282427 59198
rect 284937 59195 285003 59198
rect 286501 59195 286567 59198
rect 303061 59195 303127 59198
rect 304441 59195 304507 59198
rect 307017 59195 307083 59198
rect 309777 59195 309843 59198
rect 315297 59195 315363 59198
rect 316861 59195 316927 59198
rect 318885 59195 318951 59198
rect 324589 59195 324655 59198
rect 325693 59195 325759 59198
rect 242157 59120 242450 59122
rect 242157 59064 242162 59120
rect 242218 59064 242450 59120
rect 242157 59062 242450 59064
rect 305913 59122 305979 59125
rect 308581 59122 308647 59125
rect 305913 59120 308647 59122
rect 305913 59064 305918 59120
rect 305974 59064 308586 59120
rect 308642 59064 308647 59120
rect 305913 59062 308647 59064
rect 326662 59122 326722 59334
rect 327398 59258 327458 59334
rect 329925 59331 329991 59334
rect 332685 59331 332751 59334
rect 333237 59394 333303 59397
rect 333237 59392 334818 59394
rect 333237 59336 333242 59392
rect 333298 59336 334818 59392
rect 333237 59334 334818 59336
rect 333237 59331 333303 59334
rect 328821 59258 328887 59261
rect 327398 59256 328887 59258
rect 327398 59200 328826 59256
rect 328882 59200 328887 59256
rect 327398 59198 328887 59200
rect 328821 59195 328887 59198
rect 328637 59122 328703 59125
rect 326662 59120 328703 59122
rect 326662 59064 328642 59120
rect 328698 59064 328703 59120
rect 326662 59062 328703 59064
rect 334758 59122 334818 59334
rect 334942 59258 335002 59606
rect 335096 59394 335156 60044
rect 335353 59394 335419 59397
rect 335096 59392 335419 59394
rect 335096 59336 335358 59392
rect 335414 59336 335419 59392
rect 335096 59334 335419 59336
rect 335924 59394 335984 60044
rect 336660 59530 336720 60044
rect 337488 59666 337548 60044
rect 338316 59802 338376 60044
rect 339144 59938 339204 60044
rect 339144 59878 339234 59938
rect 339033 59802 339099 59805
rect 338316 59800 339099 59802
rect 338316 59744 339038 59800
rect 339094 59744 339099 59800
rect 338316 59742 339099 59744
rect 339033 59739 339099 59742
rect 339174 59666 339234 59878
rect 337488 59606 339050 59666
rect 338113 59530 338179 59533
rect 336660 59528 338179 59530
rect 336660 59472 338118 59528
rect 338174 59472 338179 59528
rect 336660 59470 338179 59472
rect 338113 59467 338179 59470
rect 338205 59394 338271 59397
rect 335924 59392 338271 59394
rect 335924 59336 338210 59392
rect 338266 59336 338271 59392
rect 335924 59334 338271 59336
rect 338990 59394 339050 59606
rect 339144 59606 339234 59666
rect 339972 59666 340032 60044
rect 340800 59802 340860 60044
rect 341628 59938 341688 60044
rect 341628 59878 342362 59938
rect 341517 59802 341583 59805
rect 340800 59800 341583 59802
rect 340800 59744 341522 59800
rect 341578 59744 341583 59800
rect 340800 59742 341583 59744
rect 341517 59739 341583 59742
rect 339972 59606 341442 59666
rect 339144 59530 339204 59606
rect 340965 59530 341031 59533
rect 339144 59528 341031 59530
rect 339144 59472 340970 59528
rect 341026 59472 341031 59528
rect 339144 59470 341031 59472
rect 340965 59467 341031 59470
rect 339585 59394 339651 59397
rect 338990 59392 339651 59394
rect 338990 59336 339590 59392
rect 339646 59336 339651 59392
rect 338990 59334 339651 59336
rect 341382 59394 341442 59606
rect 342302 59530 342362 59878
rect 342456 59802 342516 60044
rect 343081 59802 343147 59805
rect 342456 59800 343147 59802
rect 342456 59744 343086 59800
rect 343142 59744 343147 59800
rect 342456 59742 343147 59744
rect 343081 59739 343147 59742
rect 343284 59666 343344 60044
rect 343284 59606 344018 59666
rect 343633 59530 343699 59533
rect 342302 59528 343699 59530
rect 342302 59472 343638 59528
rect 343694 59472 343699 59528
rect 342302 59470 343699 59472
rect 343633 59467 343699 59470
rect 342345 59394 342411 59397
rect 341382 59392 342411 59394
rect 341382 59336 342350 59392
rect 342406 59336 342411 59392
rect 341382 59334 342411 59336
rect 343958 59394 344018 59606
rect 344112 59530 344172 60044
rect 344737 59530 344803 59533
rect 344112 59528 344803 59530
rect 344112 59472 344742 59528
rect 344798 59472 344803 59528
rect 344112 59470 344803 59472
rect 344940 59530 345000 60044
rect 344940 59470 345674 59530
rect 344737 59467 344803 59470
rect 345289 59394 345355 59397
rect 343958 59392 345355 59394
rect 343958 59336 345294 59392
rect 345350 59336 345355 59392
rect 343958 59334 345355 59336
rect 335353 59331 335419 59334
rect 338205 59331 338271 59334
rect 339585 59331 339651 59334
rect 342345 59331 342411 59334
rect 345289 59331 345355 59334
rect 335537 59258 335603 59261
rect 334942 59256 335603 59258
rect 334942 59200 335542 59256
rect 335598 59200 335603 59256
rect 334942 59198 335603 59200
rect 345614 59258 345674 59470
rect 345768 59394 345828 60044
rect 346596 59666 346656 60044
rect 347424 59802 347484 60044
rect 347957 59802 348023 59805
rect 347424 59800 348023 59802
rect 347424 59744 347962 59800
rect 348018 59744 348023 59800
rect 347424 59742 348023 59744
rect 347957 59739 348023 59742
rect 348049 59666 348115 59669
rect 346596 59664 348115 59666
rect 346596 59608 348054 59664
rect 348110 59608 348115 59664
rect 346596 59606 348115 59608
rect 348252 59666 348312 60044
rect 348417 59802 348483 59805
rect 349080 59802 349140 60044
rect 348417 59800 349140 59802
rect 348417 59744 348422 59800
rect 348478 59744 349140 59800
rect 348417 59742 349140 59744
rect 348417 59739 348483 59742
rect 348252 59606 349722 59666
rect 348049 59603 348115 59606
rect 347957 59530 348023 59533
rect 349245 59530 349311 59533
rect 347957 59528 349311 59530
rect 347957 59472 347962 59528
rect 348018 59472 349250 59528
rect 349306 59472 349311 59528
rect 347957 59470 349311 59472
rect 347957 59467 348023 59470
rect 349245 59467 349311 59470
rect 347865 59394 347931 59397
rect 345768 59392 347931 59394
rect 345768 59336 347870 59392
rect 347926 59336 347931 59392
rect 345768 59334 347931 59336
rect 347865 59331 347931 59334
rect 348049 59394 348115 59397
rect 349429 59394 349495 59397
rect 348049 59392 349495 59394
rect 348049 59336 348054 59392
rect 348110 59336 349434 59392
rect 349490 59336 349495 59392
rect 348049 59334 349495 59336
rect 348049 59331 348115 59334
rect 349429 59331 349495 59334
rect 346393 59258 346459 59261
rect 345614 59256 346459 59258
rect 345614 59200 346398 59256
rect 346454 59200 346459 59256
rect 345614 59198 346459 59200
rect 349662 59258 349722 59606
rect 349908 59394 349968 60044
rect 350736 59530 350796 60044
rect 351361 59530 351427 59533
rect 350736 59528 351427 59530
rect 350736 59472 351366 59528
rect 351422 59472 351427 59528
rect 350736 59470 351427 59472
rect 351361 59467 351427 59470
rect 351564 59394 351624 60044
rect 352300 59394 352360 60044
rect 353128 59530 353188 60044
rect 353956 59802 354016 60044
rect 354784 59836 354844 60044
rect 355612 59938 355672 60044
rect 355612 59878 356346 59938
rect 354784 59802 354874 59836
rect 355225 59802 355291 59805
rect 353956 59742 354690 59802
rect 354784 59800 355291 59802
rect 354784 59776 355230 59800
rect 354814 59744 355230 59776
rect 355286 59744 355291 59800
rect 354814 59742 355291 59744
rect 354630 59666 354690 59742
rect 355225 59739 355291 59742
rect 354630 59606 355242 59666
rect 354949 59530 355015 59533
rect 353128 59528 355015 59530
rect 353128 59472 354954 59528
rect 355010 59472 355015 59528
rect 353128 59470 355015 59472
rect 355182 59530 355242 59606
rect 356053 59530 356119 59533
rect 355182 59528 356119 59530
rect 355182 59472 356058 59528
rect 356114 59472 356119 59528
rect 355182 59470 356119 59472
rect 356286 59530 356346 59878
rect 356440 59666 356500 60044
rect 357065 59666 357131 59669
rect 356440 59664 357131 59666
rect 356440 59608 357070 59664
rect 357126 59608 357131 59664
rect 356440 59606 357131 59608
rect 357268 59666 357328 60044
rect 358096 59802 358156 60044
rect 358924 59938 358984 60044
rect 358924 59878 359658 59938
rect 359598 59805 359658 59878
rect 358096 59742 359290 59802
rect 358905 59666 358971 59669
rect 357268 59664 358971 59666
rect 357268 59608 358910 59664
rect 358966 59608 358971 59664
rect 357268 59606 358971 59608
rect 357065 59603 357131 59606
rect 358905 59603 358971 59606
rect 357617 59530 357683 59533
rect 356286 59528 357683 59530
rect 356286 59472 357622 59528
rect 357678 59472 357683 59528
rect 356286 59470 357683 59472
rect 359230 59530 359290 59742
rect 359549 59800 359658 59805
rect 359549 59744 359554 59800
rect 359610 59744 359658 59800
rect 359549 59742 359658 59744
rect 359549 59739 359615 59742
rect 359752 59530 359812 60044
rect 359230 59470 359658 59530
rect 359752 59470 360394 59530
rect 354949 59467 355015 59470
rect 356053 59467 356119 59470
rect 357617 59467 357683 59470
rect 354581 59394 354647 59397
rect 349908 59334 351378 59394
rect 351564 59334 352114 59394
rect 352300 59392 354647 59394
rect 352300 59336 354586 59392
rect 354642 59336 354647 59392
rect 352300 59334 354647 59336
rect 350533 59258 350599 59261
rect 349662 59256 350599 59258
rect 349662 59200 350538 59256
rect 350594 59200 350599 59256
rect 349662 59198 350599 59200
rect 351318 59258 351378 59334
rect 351913 59258 351979 59261
rect 351318 59256 351979 59258
rect 351318 59200 351918 59256
rect 351974 59200 351979 59256
rect 351318 59198 351979 59200
rect 352054 59258 352114 59334
rect 354581 59331 354647 59334
rect 355225 59394 355291 59397
rect 357065 59394 357131 59397
rect 358813 59394 358879 59397
rect 355225 59392 356898 59394
rect 355225 59336 355230 59392
rect 355286 59336 356898 59392
rect 355225 59334 356898 59336
rect 355225 59331 355291 59334
rect 353385 59258 353451 59261
rect 352054 59256 353451 59258
rect 352054 59200 353390 59256
rect 353446 59200 353451 59256
rect 352054 59198 353451 59200
rect 356838 59258 356898 59334
rect 357065 59392 358879 59394
rect 357065 59336 357070 59392
rect 357126 59336 358818 59392
rect 358874 59336 358879 59392
rect 357065 59334 358879 59336
rect 359598 59394 359658 59470
rect 360193 59394 360259 59397
rect 359598 59392 360259 59394
rect 359598 59336 360198 59392
rect 360254 59336 360259 59392
rect 359598 59334 360259 59336
rect 357065 59331 357131 59334
rect 358813 59331 358879 59334
rect 360193 59331 360259 59334
rect 357801 59258 357867 59261
rect 356838 59256 357867 59258
rect 356838 59200 357806 59256
rect 357862 59200 357867 59256
rect 356838 59198 357867 59200
rect 360334 59258 360394 59470
rect 360580 59394 360640 60044
rect 361408 59530 361468 60044
rect 362236 59666 362296 60044
rect 363064 59802 363124 60044
rect 363689 59802 363755 59805
rect 363064 59800 363755 59802
rect 363064 59744 363694 59800
rect 363750 59744 363755 59800
rect 363064 59742 363755 59744
rect 363892 59802 363952 60044
rect 364720 59938 364780 60044
rect 364720 59878 365362 59938
rect 365161 59802 365227 59805
rect 363892 59800 365227 59802
rect 363892 59744 365166 59800
rect 365222 59744 365227 59800
rect 363892 59742 365227 59744
rect 363689 59739 363755 59742
rect 365161 59739 365227 59742
rect 364977 59666 365043 59669
rect 362236 59664 365043 59666
rect 362236 59608 364982 59664
rect 365038 59608 365043 59664
rect 362236 59606 365043 59608
rect 364977 59603 365043 59606
rect 363781 59530 363847 59533
rect 361408 59528 363847 59530
rect 361408 59472 363786 59528
rect 363842 59472 363847 59528
rect 361408 59470 363847 59472
rect 363781 59467 363847 59470
rect 363597 59394 363663 59397
rect 360580 59392 363663 59394
rect 360580 59336 363602 59392
rect 363658 59336 363663 59392
rect 360580 59334 363663 59336
rect 363597 59331 363663 59334
rect 361573 59258 361639 59261
rect 360334 59256 361639 59258
rect 360334 59200 361578 59256
rect 361634 59200 361639 59256
rect 360334 59198 361639 59200
rect 335537 59195 335603 59198
rect 346393 59195 346459 59198
rect 350533 59195 350599 59198
rect 351913 59195 351979 59198
rect 353385 59195 353451 59198
rect 357801 59195 357867 59198
rect 361573 59195 361639 59198
rect 335445 59122 335511 59125
rect 334758 59120 335511 59122
rect 334758 59064 335450 59120
rect 335506 59064 335511 59120
rect 334758 59062 335511 59064
rect 365302 59122 365362 59878
rect 365548 59394 365608 60044
rect 366376 59938 366436 60044
rect 366376 59878 367018 59938
rect 366958 59805 367018 59878
rect 366958 59800 367067 59805
rect 366958 59744 367006 59800
rect 367062 59744 367067 59800
rect 366958 59742 367067 59744
rect 367001 59739 367067 59742
rect 367204 59394 367264 60044
rect 368032 59394 368092 60044
rect 368768 59802 368828 60044
rect 369393 59802 369459 59805
rect 368768 59800 369459 59802
rect 368768 59744 369398 59800
rect 369454 59744 369459 59800
rect 368768 59742 369459 59744
rect 369393 59739 369459 59742
rect 369596 59530 369656 60044
rect 370424 59802 370484 60044
rect 371049 59802 371115 59805
rect 370424 59800 371115 59802
rect 370424 59744 371054 59800
rect 371110 59744 371115 59800
rect 370424 59742 371115 59744
rect 371049 59739 371115 59742
rect 371049 59666 371115 59669
rect 369810 59664 371115 59666
rect 369810 59608 371054 59664
rect 371110 59608 371115 59664
rect 369810 59606 371115 59608
rect 369810 59530 369870 59606
rect 371049 59603 371115 59606
rect 369596 59470 369870 59530
rect 369945 59530 370011 59533
rect 370681 59530 370747 59533
rect 369945 59528 370747 59530
rect 369945 59472 369950 59528
rect 370006 59472 370686 59528
rect 370742 59472 370747 59528
rect 369945 59470 370747 59472
rect 369945 59467 370011 59470
rect 370681 59467 370747 59470
rect 369945 59394 370011 59397
rect 370497 59394 370563 59397
rect 365548 59334 367018 59394
rect 367204 59334 367938 59394
rect 368032 59392 370011 59394
rect 368032 59336 369950 59392
rect 370006 59336 370011 59392
rect 368032 59334 370011 59336
rect 366958 59258 367018 59334
rect 367737 59258 367803 59261
rect 366958 59256 367803 59258
rect 366958 59200 367742 59256
rect 367798 59200 367803 59256
rect 366958 59198 367803 59200
rect 367878 59258 367938 59334
rect 369945 59331 370011 59334
rect 370086 59392 370563 59394
rect 370086 59336 370502 59392
rect 370558 59336 370563 59392
rect 370086 59334 370563 59336
rect 371252 59394 371312 60044
rect 372080 59530 372140 60044
rect 372705 59530 372771 59533
rect 372080 59528 372771 59530
rect 372080 59472 372710 59528
rect 372766 59472 372771 59528
rect 372080 59470 372771 59472
rect 372705 59467 372771 59470
rect 372908 59394 372968 60044
rect 373736 59530 373796 60044
rect 374564 59666 374624 60044
rect 375392 59802 375452 60044
rect 376017 59802 376083 59805
rect 375392 59800 376083 59802
rect 375392 59744 376022 59800
rect 376078 59744 376083 59800
rect 375392 59742 376083 59744
rect 376017 59739 376083 59742
rect 376017 59666 376083 59669
rect 374564 59664 376083 59666
rect 374564 59608 376022 59664
rect 376078 59608 376083 59664
rect 374564 59606 376083 59608
rect 376017 59603 376083 59606
rect 376017 59530 376083 59533
rect 373736 59528 376083 59530
rect 373736 59472 376022 59528
rect 376078 59472 376083 59528
rect 373736 59470 376083 59472
rect 376017 59467 376083 59470
rect 376220 59394 376280 60044
rect 377048 59530 377108 60044
rect 377876 59666 377936 60044
rect 378501 59666 378567 59669
rect 377876 59664 378567 59666
rect 377876 59608 378506 59664
rect 378562 59608 378567 59664
rect 377876 59606 378567 59608
rect 378704 59666 378764 60044
rect 379532 59802 379592 60044
rect 380065 59802 380131 59805
rect 379532 59800 380131 59802
rect 379532 59744 380070 59800
rect 380126 59744 380131 59800
rect 379532 59742 380131 59744
rect 380360 59802 380420 60044
rect 380985 59802 381051 59805
rect 380360 59800 381051 59802
rect 380360 59744 380990 59800
rect 381046 59744 381051 59800
rect 380360 59742 381051 59744
rect 380065 59739 380131 59742
rect 380985 59739 381051 59742
rect 380985 59666 381051 59669
rect 378704 59664 381051 59666
rect 378704 59608 380990 59664
rect 381046 59608 381051 59664
rect 378704 59606 381051 59608
rect 378501 59603 378567 59606
rect 380985 59603 381051 59606
rect 379421 59530 379487 59533
rect 377048 59528 379487 59530
rect 377048 59472 379426 59528
rect 379482 59472 379487 59528
rect 377048 59470 379487 59472
rect 379421 59467 379487 59470
rect 378501 59394 378567 59397
rect 380801 59394 380867 59397
rect 371252 59334 372722 59394
rect 372908 59334 376034 59394
rect 376220 59334 378426 59394
rect 370086 59258 370146 59334
rect 370497 59331 370563 59334
rect 367878 59198 370146 59258
rect 372662 59258 372722 59334
rect 374637 59258 374703 59261
rect 372662 59256 374703 59258
rect 372662 59200 374642 59256
rect 374698 59200 374703 59256
rect 372662 59198 374703 59200
rect 375974 59258 376034 59334
rect 376201 59258 376267 59261
rect 375974 59256 376267 59258
rect 375974 59200 376206 59256
rect 376262 59200 376267 59256
rect 375974 59198 376267 59200
rect 378366 59258 378426 59334
rect 378501 59392 380867 59394
rect 378501 59336 378506 59392
rect 378562 59336 380806 59392
rect 380862 59336 380867 59392
rect 378501 59334 380867 59336
rect 381188 59394 381248 60044
rect 382016 59530 382076 60044
rect 382844 59666 382904 60044
rect 383193 59666 383259 59669
rect 382844 59664 383259 59666
rect 382844 59608 383198 59664
rect 383254 59608 383259 59664
rect 382844 59606 383259 59608
rect 383193 59603 383259 59606
rect 383469 59530 383535 59533
rect 382016 59528 383535 59530
rect 382016 59472 383474 59528
rect 383530 59472 383535 59528
rect 382016 59470 383535 59472
rect 383672 59530 383732 60044
rect 384500 59530 384560 60044
rect 385236 59666 385296 60044
rect 385861 59666 385927 59669
rect 385236 59664 385927 59666
rect 385236 59608 385866 59664
rect 385922 59608 385927 59664
rect 385236 59606 385927 59608
rect 386064 59666 386124 60044
rect 386892 59802 386952 60044
rect 387517 59802 387583 59805
rect 386892 59800 387583 59802
rect 386892 59744 387522 59800
rect 387578 59744 387583 59800
rect 386892 59742 387583 59744
rect 387517 59739 387583 59742
rect 386064 59606 387626 59666
rect 385861 59603 385927 59606
rect 387241 59530 387307 59533
rect 383672 59470 384314 59530
rect 384500 59528 387307 59530
rect 384500 59472 387246 59528
rect 387302 59472 387307 59528
rect 384500 59470 387307 59472
rect 383469 59467 383535 59470
rect 383193 59394 383259 59397
rect 384113 59394 384179 59397
rect 381188 59334 382658 59394
rect 378501 59331 378567 59334
rect 380801 59331 380867 59334
rect 378777 59258 378843 59261
rect 378366 59256 378843 59258
rect 378366 59200 378782 59256
rect 378838 59200 378843 59256
rect 378366 59198 378843 59200
rect 382598 59258 382658 59334
rect 383193 59392 384179 59394
rect 383193 59336 383198 59392
rect 383254 59336 384118 59392
rect 384174 59336 384179 59392
rect 383193 59334 384179 59336
rect 384254 59394 384314 59470
rect 387241 59467 387307 59470
rect 385861 59394 385927 59397
rect 387566 59394 387626 59606
rect 387720 59530 387780 60044
rect 388548 59666 388608 60044
rect 389376 59802 389436 60044
rect 390001 59802 390067 59805
rect 389376 59800 390067 59802
rect 389376 59744 390006 59800
rect 390062 59744 390067 59800
rect 389376 59742 390067 59744
rect 390204 59802 390264 60044
rect 390829 59802 390895 59805
rect 390204 59800 390895 59802
rect 390204 59744 390834 59800
rect 390890 59744 390895 59800
rect 390204 59742 390895 59744
rect 391032 59802 391092 60044
rect 391657 59802 391723 59805
rect 391032 59800 391723 59802
rect 391032 59744 391662 59800
rect 391718 59744 391723 59800
rect 391032 59742 391723 59744
rect 390001 59739 390067 59742
rect 390829 59739 390895 59742
rect 391657 59739 391723 59742
rect 391197 59666 391263 59669
rect 388548 59664 391263 59666
rect 388548 59608 391202 59664
rect 391258 59608 391263 59664
rect 388548 59606 391263 59608
rect 391197 59603 391263 59606
rect 390001 59530 390067 59533
rect 387720 59528 390067 59530
rect 387720 59472 390006 59528
rect 390062 59472 390067 59528
rect 387720 59470 390067 59472
rect 391860 59530 391920 60044
rect 392688 59666 392748 60044
rect 393313 59666 393379 59669
rect 392688 59664 393379 59666
rect 392688 59608 393318 59664
rect 393374 59608 393379 59664
rect 392688 59606 393379 59608
rect 393313 59603 393379 59606
rect 393313 59530 393379 59533
rect 391860 59528 393379 59530
rect 391860 59472 393318 59528
rect 393374 59472 393379 59528
rect 391860 59470 393379 59472
rect 390001 59467 390067 59470
rect 393313 59467 393379 59470
rect 388621 59394 388687 59397
rect 384254 59334 385786 59394
rect 383193 59331 383259 59334
rect 384113 59331 384179 59334
rect 384297 59258 384363 59261
rect 382598 59256 384363 59258
rect 382598 59200 384302 59256
rect 384358 59200 384363 59256
rect 382598 59198 384363 59200
rect 385726 59258 385786 59334
rect 385861 59392 387442 59394
rect 385861 59336 385866 59392
rect 385922 59336 387442 59392
rect 385861 59334 387442 59336
rect 387566 59392 388687 59394
rect 387566 59336 388626 59392
rect 388682 59336 388687 59392
rect 387566 59334 388687 59336
rect 385861 59331 385927 59334
rect 387057 59258 387123 59261
rect 385726 59256 387123 59258
rect 385726 59200 387062 59256
rect 387118 59200 387123 59256
rect 385726 59198 387123 59200
rect 387382 59258 387442 59334
rect 388621 59331 388687 59334
rect 390829 59394 390895 59397
rect 392761 59394 392827 59397
rect 390829 59392 392827 59394
rect 390829 59336 390834 59392
rect 390890 59336 392766 59392
rect 392822 59336 392827 59392
rect 390829 59334 392827 59336
rect 393516 59394 393576 60044
rect 393681 59530 393747 59533
rect 394141 59530 394207 59533
rect 393681 59528 394207 59530
rect 393681 59472 393686 59528
rect 393742 59472 394146 59528
rect 394202 59472 394207 59528
rect 393681 59470 394207 59472
rect 394344 59530 394404 60044
rect 395172 59666 395232 60044
rect 395797 59666 395863 59669
rect 395172 59664 395863 59666
rect 395172 59608 395802 59664
rect 395858 59608 395863 59664
rect 395172 59606 395863 59608
rect 396000 59666 396060 60044
rect 396828 59802 396888 60044
rect 397453 59802 397519 59805
rect 396828 59800 397519 59802
rect 396828 59744 397458 59800
rect 397514 59744 397519 59800
rect 396828 59742 397519 59744
rect 397453 59739 397519 59742
rect 397453 59666 397519 59669
rect 396000 59664 397519 59666
rect 396000 59608 397458 59664
rect 397514 59608 397519 59664
rect 396000 59606 397519 59608
rect 395797 59603 395863 59606
rect 397453 59603 397519 59606
rect 396717 59530 396783 59533
rect 394344 59528 396783 59530
rect 394344 59472 396722 59528
rect 396778 59472 396783 59528
rect 394344 59470 396783 59472
rect 397656 59530 397716 60044
rect 397821 59666 397887 59669
rect 398281 59666 398347 59669
rect 397821 59664 398347 59666
rect 397821 59608 397826 59664
rect 397882 59608 398286 59664
rect 398342 59608 398347 59664
rect 397821 59606 398347 59608
rect 397821 59603 397887 59606
rect 398281 59603 398347 59606
rect 398097 59530 398163 59533
rect 397656 59528 398163 59530
rect 397656 59472 398102 59528
rect 398158 59472 398163 59528
rect 397656 59470 398163 59472
rect 398484 59530 398544 60044
rect 399312 59666 399372 60044
rect 399937 59666 400003 59669
rect 399312 59664 400003 59666
rect 399312 59608 399942 59664
rect 399998 59608 400003 59664
rect 399312 59606 400003 59608
rect 400140 59666 400200 60044
rect 400765 59666 400831 59669
rect 400140 59664 400831 59666
rect 400140 59608 400770 59664
rect 400826 59608 400831 59664
rect 400140 59606 400831 59608
rect 400968 59666 401028 60044
rect 401704 59802 401764 60044
rect 402329 59802 402395 59805
rect 401704 59800 402395 59802
rect 401704 59744 402334 59800
rect 402390 59744 402395 59800
rect 401704 59742 402395 59744
rect 402329 59739 402395 59742
rect 400968 59606 401978 59666
rect 399937 59603 400003 59606
rect 400765 59603 400831 59606
rect 400857 59530 400923 59533
rect 398484 59528 400923 59530
rect 398484 59472 400862 59528
rect 400918 59472 400923 59528
rect 398484 59470 400923 59472
rect 393681 59467 393747 59470
rect 394141 59467 394207 59470
rect 396717 59467 396783 59470
rect 398097 59467 398163 59470
rect 400857 59467 400923 59470
rect 395797 59394 395863 59397
rect 398005 59394 398071 59397
rect 393516 59334 395722 59394
rect 390829 59331 390895 59334
rect 392761 59331 392827 59334
rect 388437 59258 388503 59261
rect 387382 59256 388503 59258
rect 387382 59200 388442 59256
rect 388498 59200 388503 59256
rect 387382 59198 388503 59200
rect 395662 59258 395722 59334
rect 395797 59392 398071 59394
rect 395797 59336 395802 59392
rect 395858 59336 398010 59392
rect 398066 59336 398071 59392
rect 395797 59334 398071 59336
rect 395797 59331 395863 59334
rect 398005 59331 398071 59334
rect 399937 59394 400003 59397
rect 400765 59394 400831 59397
rect 401593 59394 401659 59397
rect 399937 59392 400690 59394
rect 399937 59336 399942 59392
rect 399998 59336 400690 59392
rect 399937 59334 400690 59336
rect 399937 59331 400003 59334
rect 396901 59258 396967 59261
rect 395662 59256 396967 59258
rect 395662 59200 396906 59256
rect 396962 59200 396967 59256
rect 395662 59198 396967 59200
rect 400630 59258 400690 59334
rect 400765 59392 401659 59394
rect 400765 59336 400770 59392
rect 400826 59336 401598 59392
rect 401654 59336 401659 59392
rect 400765 59334 401659 59336
rect 401918 59394 401978 59606
rect 402532 59530 402592 60044
rect 402532 59470 403266 59530
rect 403065 59394 403131 59397
rect 401918 59392 403131 59394
rect 401918 59336 403070 59392
rect 403126 59336 403131 59392
rect 401918 59334 403131 59336
rect 400765 59331 400831 59334
rect 401593 59331 401659 59334
rect 403065 59331 403131 59334
rect 402237 59258 402303 59261
rect 400630 59256 402303 59258
rect 400630 59200 402242 59256
rect 402298 59200 402303 59256
rect 400630 59198 402303 59200
rect 403206 59258 403266 59470
rect 403360 59394 403420 60044
rect 404188 59530 404248 60044
rect 405016 59666 405076 60044
rect 405844 59802 405904 60044
rect 406469 59802 406535 59805
rect 405844 59800 406535 59802
rect 405844 59744 406474 59800
rect 406530 59744 406535 59800
rect 405844 59742 406535 59744
rect 406469 59739 406535 59742
rect 405016 59606 406578 59666
rect 405917 59530 405983 59533
rect 404188 59528 405983 59530
rect 404188 59472 405922 59528
rect 405978 59472 405983 59528
rect 404188 59470 405983 59472
rect 405917 59467 405983 59470
rect 406101 59394 406167 59397
rect 403360 59392 406167 59394
rect 403360 59336 406106 59392
rect 406162 59336 406167 59392
rect 403360 59334 406167 59336
rect 406101 59331 406167 59334
rect 404353 59258 404419 59261
rect 403206 59256 404419 59258
rect 403206 59200 404358 59256
rect 404414 59200 404419 59256
rect 403206 59198 404419 59200
rect 406518 59258 406578 59606
rect 406672 59394 406732 60044
rect 407500 59530 407560 60044
rect 408125 59530 408191 59533
rect 407500 59528 408191 59530
rect 407500 59472 408130 59528
rect 408186 59472 408191 59528
rect 407500 59470 408191 59472
rect 408328 59530 408388 60044
rect 409156 59666 409216 60044
rect 409984 59802 410044 60044
rect 410609 59802 410675 59805
rect 409984 59800 410675 59802
rect 409984 59744 410614 59800
rect 410670 59744 410675 59800
rect 409984 59742 410675 59744
rect 410609 59739 410675 59742
rect 409156 59606 410626 59666
rect 409965 59530 410031 59533
rect 408328 59528 410031 59530
rect 408328 59472 409970 59528
rect 410026 59472 410031 59528
rect 408328 59470 410031 59472
rect 408125 59467 408191 59470
rect 409965 59467 410031 59470
rect 408677 59394 408743 59397
rect 406672 59392 408743 59394
rect 406672 59336 408682 59392
rect 408738 59336 408743 59392
rect 406672 59334 408743 59336
rect 410566 59394 410626 59606
rect 410812 59530 410872 60044
rect 411640 59666 411700 60044
rect 412081 59666 412147 59669
rect 411640 59664 412147 59666
rect 411640 59608 412086 59664
rect 412142 59608 412147 59664
rect 411640 59606 412147 59608
rect 412468 59666 412528 60044
rect 413093 59666 413159 59669
rect 412468 59664 413159 59666
rect 412468 59608 413098 59664
rect 413154 59608 413159 59664
rect 412468 59606 413159 59608
rect 412081 59603 412147 59606
rect 413093 59603 413159 59606
rect 412725 59530 412791 59533
rect 410812 59470 411546 59530
rect 411345 59394 411411 59397
rect 410566 59392 411411 59394
rect 410566 59336 411350 59392
rect 411406 59336 411411 59392
rect 410566 59334 411411 59336
rect 411486 59394 411546 59470
rect 411854 59528 412791 59530
rect 411854 59472 412730 59528
rect 412786 59472 412791 59528
rect 411854 59470 412791 59472
rect 411854 59394 411914 59470
rect 412725 59467 412791 59470
rect 412909 59530 412975 59533
rect 413296 59530 413356 60044
rect 412909 59528 413356 59530
rect 412909 59472 412914 59528
rect 412970 59472 413356 59528
rect 412909 59470 413356 59472
rect 412909 59467 412975 59470
rect 411486 59334 411914 59394
rect 412081 59394 412147 59397
rect 413921 59394 413987 59397
rect 412081 59392 413987 59394
rect 412081 59336 412086 59392
rect 412142 59336 413926 59392
rect 413982 59336 413987 59392
rect 412081 59334 413987 59336
rect 414124 59394 414184 60044
rect 414952 59530 415012 60044
rect 415780 59666 415840 60044
rect 416608 59938 416668 60044
rect 417344 59938 417404 60044
rect 416608 59878 416698 59938
rect 416405 59666 416471 59669
rect 415780 59664 416471 59666
rect 415780 59608 416410 59664
rect 416466 59608 416471 59664
rect 415780 59606 416471 59608
rect 416638 59666 416698 59878
rect 417006 59878 417404 59938
rect 416865 59802 416931 59805
rect 417006 59802 417066 59878
rect 416865 59800 417066 59802
rect 416865 59744 416870 59800
rect 416926 59744 417066 59800
rect 416865 59742 417066 59744
rect 416865 59739 416931 59742
rect 416638 59606 417250 59666
rect 416405 59603 416471 59606
rect 416773 59530 416839 59533
rect 414952 59528 416839 59530
rect 414952 59472 416778 59528
rect 416834 59472 416839 59528
rect 414952 59470 416839 59472
rect 416773 59467 416839 59470
rect 416957 59394 417023 59397
rect 414124 59392 417023 59394
rect 414124 59336 416962 59392
rect 417018 59336 417023 59392
rect 414124 59334 417023 59336
rect 417190 59394 417250 59606
rect 418172 59530 418232 60044
rect 419000 59938 419060 60044
rect 419828 59938 419888 60044
rect 419000 59878 419458 59938
rect 419398 59666 419458 59878
rect 419582 59878 419888 59938
rect 420656 59938 420716 60044
rect 420656 59878 421298 59938
rect 419582 59805 419642 59878
rect 419533 59800 419642 59805
rect 419533 59744 419538 59800
rect 419594 59744 419642 59800
rect 419533 59742 419642 59744
rect 419533 59739 419599 59742
rect 420913 59666 420979 59669
rect 419398 59664 420979 59666
rect 419398 59608 420918 59664
rect 420974 59608 420979 59664
rect 419398 59606 420979 59608
rect 420913 59603 420979 59606
rect 418172 59470 418906 59530
rect 418153 59394 418219 59397
rect 417190 59392 418219 59394
rect 417190 59336 418158 59392
rect 418214 59336 418219 59392
rect 417190 59334 418219 59336
rect 408677 59331 408743 59334
rect 411345 59331 411411 59334
rect 412081 59331 412147 59334
rect 413921 59331 413987 59334
rect 416957 59331 417023 59334
rect 418153 59331 418219 59334
rect 407297 59258 407363 59261
rect 406518 59256 407363 59258
rect 406518 59200 407302 59256
rect 407358 59200 407363 59256
rect 406518 59198 407363 59200
rect 418846 59258 418906 59470
rect 421238 59394 421298 59878
rect 421484 59530 421544 60044
rect 422312 59666 422372 60044
rect 422312 59606 422954 59666
rect 421484 59470 422770 59530
rect 422385 59394 422451 59397
rect 421238 59392 422451 59394
rect 421238 59336 422390 59392
rect 422446 59336 422451 59392
rect 421238 59334 422451 59336
rect 422385 59331 422451 59334
rect 421097 59258 421163 59261
rect 418846 59256 421163 59258
rect 418846 59200 421102 59256
rect 421158 59200 421163 59256
rect 418846 59198 421163 59200
rect 422710 59258 422770 59470
rect 422894 59394 422954 59606
rect 423140 59530 423200 60044
rect 423968 59666 424028 60044
rect 424796 59802 424856 60044
rect 425624 59938 425684 60044
rect 426452 59938 426512 60044
rect 425624 59878 426082 59938
rect 426452 59878 427002 59938
rect 425513 59802 425579 59805
rect 424796 59800 425579 59802
rect 424796 59744 425518 59800
rect 425574 59744 425579 59800
rect 424796 59742 425579 59744
rect 425513 59739 425579 59742
rect 423968 59606 425530 59666
rect 425329 59530 425395 59533
rect 423140 59528 425395 59530
rect 423140 59472 425334 59528
rect 425390 59472 425395 59528
rect 423140 59470 425395 59472
rect 425329 59467 425395 59470
rect 425145 59394 425211 59397
rect 422894 59392 425211 59394
rect 422894 59336 425150 59392
rect 425206 59336 425211 59392
rect 422894 59334 425211 59336
rect 425470 59394 425530 59606
rect 426022 59530 426082 59878
rect 426942 59802 427002 59878
rect 427077 59802 427143 59805
rect 426942 59800 427143 59802
rect 426942 59744 427082 59800
rect 427138 59744 427143 59800
rect 426942 59742 427143 59744
rect 427077 59739 427143 59742
rect 426022 59470 427186 59530
rect 425470 59334 426082 59394
rect 425145 59331 425211 59334
rect 423765 59258 423831 59261
rect 422710 59256 423831 59258
rect 422710 59200 423770 59256
rect 423826 59200 423831 59256
rect 422710 59198 423831 59200
rect 426022 59258 426082 59334
rect 426433 59258 426499 59261
rect 426022 59256 426499 59258
rect 426022 59200 426438 59256
rect 426494 59200 426499 59256
rect 426022 59198 426499 59200
rect 427126 59258 427186 59470
rect 427280 59394 427340 60044
rect 428108 59530 428168 60044
rect 428733 59530 428799 59533
rect 428108 59528 428799 59530
rect 428108 59472 428738 59528
rect 428794 59472 428799 59528
rect 428108 59470 428799 59472
rect 428936 59530 428996 60044
rect 429764 59666 429824 60044
rect 430592 59802 430652 60044
rect 431217 59802 431283 59805
rect 430592 59800 431283 59802
rect 430592 59744 431222 59800
rect 431278 59744 431283 59800
rect 430592 59742 431283 59744
rect 431217 59739 431283 59742
rect 429764 59606 430866 59666
rect 430573 59530 430639 59533
rect 428936 59528 430639 59530
rect 428936 59472 430578 59528
rect 430634 59472 430639 59528
rect 428936 59470 430639 59472
rect 428733 59467 428799 59470
rect 430573 59467 430639 59470
rect 429377 59394 429443 59397
rect 427280 59392 429443 59394
rect 427280 59336 429382 59392
rect 429438 59336 429443 59392
rect 427280 59334 429443 59336
rect 430806 59394 430866 59606
rect 431420 59530 431480 60044
rect 432045 59530 432111 59533
rect 431420 59528 432111 59530
rect 431420 59472 432050 59528
rect 432106 59472 432111 59528
rect 431420 59470 432111 59472
rect 432045 59467 432111 59470
rect 432045 59394 432111 59397
rect 430806 59392 432111 59394
rect 430806 59336 432050 59392
rect 432106 59336 432111 59392
rect 430806 59334 432111 59336
rect 432248 59394 432308 60044
rect 433076 59530 433136 60044
rect 433812 59666 433872 60044
rect 434640 59802 434700 60044
rect 435468 59938 435528 60044
rect 436296 59938 436356 60044
rect 435468 59878 436202 59938
rect 436296 59878 436938 59938
rect 435449 59802 435515 59805
rect 434640 59800 435515 59802
rect 434640 59744 435454 59800
rect 435510 59744 435515 59800
rect 434640 59742 435515 59744
rect 435449 59739 435515 59742
rect 436142 59666 436202 59878
rect 436878 59805 436938 59878
rect 436878 59800 436987 59805
rect 436878 59744 436926 59800
rect 436982 59744 436987 59800
rect 436878 59742 436987 59744
rect 436921 59739 436987 59742
rect 433812 59606 435282 59666
rect 436142 59606 436938 59666
rect 434713 59530 434779 59533
rect 433076 59528 434779 59530
rect 433076 59472 434718 59528
rect 434774 59472 434779 59528
rect 433076 59470 434779 59472
rect 434713 59467 434779 59470
rect 434897 59394 434963 59397
rect 432248 59392 434963 59394
rect 432248 59336 434902 59392
rect 434958 59336 434963 59392
rect 432248 59334 434963 59336
rect 429377 59331 429443 59334
rect 432045 59331 432111 59334
rect 434897 59331 434963 59334
rect 427905 59258 427971 59261
rect 427126 59256 427971 59258
rect 427126 59200 427910 59256
rect 427966 59200 427971 59256
rect 427126 59198 427971 59200
rect 435222 59258 435282 59606
rect 435633 59530 435699 59533
rect 436369 59530 436435 59533
rect 435633 59528 436435 59530
rect 435633 59472 435638 59528
rect 435694 59472 436374 59528
rect 436430 59472 436435 59528
rect 435633 59470 436435 59472
rect 435633 59467 435699 59470
rect 436369 59467 436435 59470
rect 436878 59394 436938 59606
rect 437124 59530 437184 60044
rect 437952 59666 438012 60044
rect 438577 59666 438643 59669
rect 437952 59664 438643 59666
rect 437952 59608 438582 59664
rect 438638 59608 438643 59664
rect 437952 59606 438643 59608
rect 438780 59666 438840 60044
rect 439608 59802 439668 60044
rect 440233 59802 440299 59805
rect 439608 59800 440299 59802
rect 439608 59744 440238 59800
rect 440294 59744 440299 59800
rect 439608 59742 440299 59744
rect 440436 59802 440496 60044
rect 441264 59938 441324 60044
rect 441264 59878 441354 59938
rect 441153 59802 441219 59805
rect 440436 59800 441219 59802
rect 440436 59744 441158 59800
rect 441214 59744 441219 59800
rect 440436 59742 441219 59744
rect 440233 59739 440299 59742
rect 441153 59739 441219 59742
rect 440417 59666 440483 59669
rect 441294 59666 441354 59878
rect 441429 59802 441495 59805
rect 441889 59802 441955 59805
rect 441429 59800 441955 59802
rect 441429 59744 441434 59800
rect 441490 59744 441894 59800
rect 441950 59744 441955 59800
rect 441429 59742 441955 59744
rect 441429 59739 441495 59742
rect 441889 59739 441955 59742
rect 438780 59664 440483 59666
rect 438780 59608 440422 59664
rect 440478 59608 440483 59664
rect 438780 59606 440483 59608
rect 438577 59603 438643 59606
rect 440417 59603 440483 59606
rect 441264 59606 441354 59666
rect 439037 59530 439103 59533
rect 437124 59528 439103 59530
rect 437124 59472 439042 59528
rect 439098 59472 439103 59528
rect 437124 59470 439103 59472
rect 439037 59467 439103 59470
rect 437473 59394 437539 59397
rect 436878 59392 437539 59394
rect 436878 59336 437478 59392
rect 437534 59336 437539 59392
rect 436878 59334 437539 59336
rect 437473 59331 437539 59334
rect 438577 59394 438643 59397
rect 440233 59394 440299 59397
rect 441264 59394 441324 59606
rect 442092 59394 442152 60044
rect 442920 59530 442980 60044
rect 443748 59666 443808 60044
rect 444576 59802 444636 60044
rect 445404 59938 445464 60044
rect 446232 59938 446292 60044
rect 445404 59878 446138 59938
rect 446232 59878 446874 59938
rect 445937 59802 446003 59805
rect 444576 59800 446003 59802
rect 444576 59744 445942 59800
rect 445998 59744 446003 59800
rect 444576 59742 446003 59744
rect 445937 59739 446003 59742
rect 445845 59666 445911 59669
rect 443748 59664 445911 59666
rect 443748 59608 445850 59664
rect 445906 59608 445911 59664
rect 443748 59606 445911 59608
rect 446078 59666 446138 59878
rect 446814 59805 446874 59878
rect 446814 59800 446923 59805
rect 446814 59744 446862 59800
rect 446918 59744 446923 59800
rect 446814 59742 446923 59744
rect 446857 59739 446923 59742
rect 446857 59666 446923 59669
rect 446078 59664 446923 59666
rect 446078 59608 446862 59664
rect 446918 59608 446923 59664
rect 446078 59606 446923 59608
rect 445845 59603 445911 59606
rect 446857 59603 446923 59606
rect 444373 59530 444439 59533
rect 442920 59528 444439 59530
rect 442920 59472 444378 59528
rect 444434 59472 444439 59528
rect 442920 59470 444439 59472
rect 447060 59530 447120 60044
rect 447888 59666 447948 60044
rect 448716 59802 448776 60044
rect 449544 59938 449604 60044
rect 449544 59878 449818 59938
rect 449758 59805 449818 59878
rect 449341 59802 449407 59805
rect 448716 59800 449407 59802
rect 448716 59744 449346 59800
rect 449402 59744 449407 59800
rect 448716 59742 449407 59744
rect 449341 59739 449407 59742
rect 449709 59800 449818 59805
rect 449709 59744 449714 59800
rect 449770 59744 449818 59800
rect 449709 59742 449818 59744
rect 449709 59739 449775 59742
rect 449249 59666 449315 59669
rect 447888 59664 449315 59666
rect 447888 59608 449254 59664
rect 449310 59608 449315 59664
rect 447888 59606 449315 59608
rect 449249 59603 449315 59606
rect 448605 59530 448671 59533
rect 447060 59528 448671 59530
rect 447060 59472 448610 59528
rect 448666 59472 448671 59528
rect 447060 59470 448671 59472
rect 444373 59467 444439 59470
rect 448605 59467 448671 59470
rect 444465 59394 444531 59397
rect 438577 59392 439514 59394
rect 438577 59336 438582 59392
rect 438638 59336 439514 59392
rect 438577 59334 439514 59336
rect 438577 59331 438643 59334
rect 436185 59258 436251 59261
rect 435222 59256 436251 59258
rect 435222 59200 436190 59256
rect 436246 59200 436251 59256
rect 435222 59198 436251 59200
rect 439454 59258 439514 59334
rect 440233 59392 441170 59394
rect 440233 59336 440238 59392
rect 440294 59336 441170 59392
rect 440233 59334 441170 59336
rect 441264 59334 441906 59394
rect 442092 59392 444531 59394
rect 442092 59336 444470 59392
rect 444526 59336 444531 59392
rect 442092 59334 444531 59336
rect 440233 59331 440299 59334
rect 440233 59258 440299 59261
rect 439454 59256 440299 59258
rect 439454 59200 440238 59256
rect 440294 59200 440299 59256
rect 439454 59198 440299 59200
rect 441110 59258 441170 59334
rect 441705 59258 441771 59261
rect 441110 59256 441771 59258
rect 441110 59200 441710 59256
rect 441766 59200 441771 59256
rect 441110 59198 441771 59200
rect 441846 59258 441906 59334
rect 444465 59331 444531 59334
rect 445937 59394 446003 59397
rect 447409 59394 447475 59397
rect 445937 59392 447475 59394
rect 445937 59336 445942 59392
rect 445998 59336 447414 59392
rect 447470 59336 447475 59392
rect 445937 59334 447475 59336
rect 445937 59331 446003 59334
rect 447409 59331 447475 59334
rect 449341 59394 449407 59397
rect 450280 59394 450340 60044
rect 451108 59530 451168 60044
rect 451108 59470 451842 59530
rect 449341 59392 450186 59394
rect 449341 59336 449346 59392
rect 449402 59336 450186 59392
rect 449341 59334 450186 59336
rect 450280 59334 451658 59394
rect 449341 59331 449407 59334
rect 443361 59258 443427 59261
rect 441846 59256 443427 59258
rect 441846 59200 443366 59256
rect 443422 59200 443427 59256
rect 441846 59198 443427 59200
rect 450126 59258 450186 59334
rect 451273 59258 451339 59261
rect 450126 59256 451339 59258
rect 450126 59200 451278 59256
rect 451334 59200 451339 59256
rect 450126 59198 451339 59200
rect 367737 59195 367803 59198
rect 374637 59195 374703 59198
rect 376201 59195 376267 59198
rect 378777 59195 378843 59198
rect 384297 59195 384363 59198
rect 387057 59195 387123 59198
rect 388437 59195 388503 59198
rect 396901 59195 396967 59198
rect 402237 59195 402303 59198
rect 404353 59195 404419 59198
rect 407297 59195 407363 59198
rect 421097 59195 421163 59198
rect 423765 59195 423831 59198
rect 426433 59195 426499 59198
rect 427905 59195 427971 59198
rect 436185 59195 436251 59198
rect 440233 59195 440299 59198
rect 441705 59195 441771 59198
rect 443361 59195 443427 59198
rect 451273 59195 451339 59198
rect 367737 59122 367803 59125
rect 365302 59120 367803 59122
rect 365302 59064 367742 59120
rect 367798 59064 367803 59120
rect 365302 59062 367803 59064
rect 451598 59122 451658 59334
rect 451782 59258 451842 59470
rect 451936 59394 451996 60044
rect 452764 59666 452824 60044
rect 453389 59666 453455 59669
rect 452764 59664 453455 59666
rect 452764 59608 453394 59664
rect 453450 59608 453455 59664
rect 452764 59606 453455 59608
rect 453389 59603 453455 59606
rect 453592 59394 453652 60044
rect 454420 59530 454480 60044
rect 455045 59530 455111 59533
rect 454420 59528 455111 59530
rect 454420 59472 455050 59528
rect 455106 59472 455111 59528
rect 454420 59470 455111 59472
rect 455248 59530 455308 60044
rect 456076 59666 456136 60044
rect 456904 59802 456964 60044
rect 457529 59802 457595 59805
rect 456904 59800 457595 59802
rect 456904 59744 457534 59800
rect 457590 59744 457595 59800
rect 456904 59742 457595 59744
rect 457529 59739 457595 59742
rect 456076 59606 457546 59666
rect 456793 59530 456859 59533
rect 455248 59528 456859 59530
rect 455248 59472 456798 59528
rect 456854 59472 456859 59528
rect 455248 59470 456859 59472
rect 455045 59467 455111 59470
rect 456793 59467 456859 59470
rect 455505 59394 455571 59397
rect 451936 59334 453498 59394
rect 453592 59392 455571 59394
rect 453592 59336 455510 59392
rect 455566 59336 455571 59392
rect 453592 59334 455571 59336
rect 452745 59258 452811 59261
rect 451782 59256 452811 59258
rect 451782 59200 452750 59256
rect 452806 59200 452811 59256
rect 451782 59198 452811 59200
rect 453438 59258 453498 59334
rect 455505 59331 455571 59334
rect 454033 59258 454099 59261
rect 453438 59256 454099 59258
rect 453438 59200 454038 59256
rect 454094 59200 454099 59256
rect 453438 59198 454099 59200
rect 457486 59258 457546 59606
rect 457732 59394 457792 60044
rect 458560 59530 458620 60044
rect 459185 59530 459251 59533
rect 458560 59528 459251 59530
rect 458560 59472 459190 59528
rect 459246 59472 459251 59528
rect 458560 59470 459251 59472
rect 459185 59467 459251 59470
rect 459388 59394 459448 60044
rect 460216 59666 460276 60044
rect 461044 59802 461104 60044
rect 461577 59802 461643 59805
rect 461044 59800 461643 59802
rect 461044 59744 461582 59800
rect 461638 59744 461643 59800
rect 461044 59742 461643 59744
rect 461577 59739 461643 59742
rect 461669 59666 461735 59669
rect 460216 59664 461735 59666
rect 460216 59608 461674 59664
rect 461730 59608 461735 59664
rect 460216 59606 461735 59608
rect 461669 59603 461735 59606
rect 461872 59530 461932 60044
rect 462700 59666 462760 60044
rect 463528 59802 463588 60044
rect 464153 59802 464219 59805
rect 463528 59800 464219 59802
rect 463528 59744 464158 59800
rect 464214 59744 464219 59800
rect 463528 59742 464219 59744
rect 464153 59739 464219 59742
rect 462700 59606 464170 59666
rect 463969 59530 464035 59533
rect 461872 59528 464035 59530
rect 461872 59472 463974 59528
rect 464030 59472 464035 59528
rect 461872 59470 464035 59472
rect 463969 59467 464035 59470
rect 461577 59394 461643 59397
rect 463785 59394 463851 59397
rect 457732 59334 459202 59394
rect 459388 59334 460950 59394
rect 458265 59258 458331 59261
rect 457486 59256 458331 59258
rect 457486 59200 458270 59256
rect 458326 59200 458331 59256
rect 457486 59198 458331 59200
rect 459142 59258 459202 59334
rect 459737 59258 459803 59261
rect 459142 59256 459803 59258
rect 459142 59200 459742 59256
rect 459798 59200 459803 59256
rect 459142 59198 459803 59200
rect 460890 59258 460950 59334
rect 461577 59392 463851 59394
rect 461577 59336 461582 59392
rect 461638 59336 463790 59392
rect 463846 59336 463851 59392
rect 461577 59334 463851 59336
rect 461577 59331 461643 59334
rect 463785 59331 463851 59334
rect 461025 59258 461091 59261
rect 460890 59256 461091 59258
rect 460890 59200 461030 59256
rect 461086 59200 461091 59256
rect 460890 59198 461091 59200
rect 464110 59258 464170 59606
rect 464356 59394 464416 60044
rect 465184 59530 465244 60044
rect 467833 59530 467899 59533
rect 465184 59528 467899 59530
rect 465184 59472 467838 59528
rect 467894 59472 467899 59528
rect 583520 59516 584960 59756
rect 465184 59470 467899 59472
rect 467833 59467 467899 59470
rect 466545 59394 466611 59397
rect 464356 59392 466611 59394
rect 464356 59336 466550 59392
rect 466606 59336 466611 59392
rect 464356 59334 466611 59336
rect 466545 59331 466611 59334
rect 465073 59258 465139 59261
rect 464110 59256 465139 59258
rect 464110 59200 465078 59256
rect 465134 59200 465139 59256
rect 464110 59198 465139 59200
rect 452745 59195 452811 59198
rect 454033 59195 454099 59198
rect 458265 59195 458331 59198
rect 459737 59195 459803 59198
rect 461025 59195 461091 59198
rect 465073 59195 465139 59198
rect 452929 59122 452995 59125
rect 451598 59120 452995 59122
rect 451598 59064 452934 59120
rect 452990 59064 452995 59120
rect 451598 59062 452995 59064
rect 180812 59060 180818 59062
rect 181989 59059 182055 59062
rect 183369 59059 183435 59062
rect 191741 59059 191807 59062
rect 220629 59059 220695 59062
rect 231117 59059 231183 59062
rect 242157 59059 242223 59062
rect 305913 59059 305979 59062
rect 308581 59059 308647 59062
rect 328637 59059 328703 59062
rect 335445 59059 335511 59062
rect 367737 59059 367803 59062
rect 452929 59059 452995 59062
rect 72969 58984 74274 58986
rect 72969 58928 72974 58984
rect 73030 58928 74274 58984
rect 72969 58926 74274 58928
rect 72969 58923 73035 58926
rect 291878 58924 291884 58988
rect 291948 58986 291954 58988
rect 294505 58986 294571 58989
rect 291948 58984 294571 58986
rect 291948 58928 294510 58984
rect 294566 58928 294571 58984
rect 291948 58926 294571 58928
rect 291948 58924 291954 58926
rect 294505 58923 294571 58926
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
rect 19425 3362 19491 3365
rect 86217 3362 86283 3365
rect 19425 3360 86283 3362
rect 19425 3304 19430 3360
rect 19486 3304 86222 3360
rect 86278 3304 86283 3360
rect 19425 3302 86283 3304
rect 19425 3299 19491 3302
rect 86217 3299 86283 3302
rect 144821 3362 144887 3365
rect 583385 3362 583451 3365
rect 144821 3360 583451 3362
rect 144821 3304 144826 3360
rect 144882 3304 583390 3360
rect 583446 3304 583451 3360
rect 144821 3302 583451 3304
rect 144821 3299 144887 3302
rect 583385 3299 583451 3302
<< via3 >>
rect 180748 59392 180812 59396
rect 180748 59336 180762 59392
rect 180762 59336 180812 59392
rect 180748 59332 180812 59336
rect 180748 59060 180812 59124
rect 291884 59740 291948 59804
rect 291884 58924 291948 58988
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 447968 60134 456618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 447968 63854 460338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 447968 67574 464058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 447968 74414 470898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 447968 78134 474618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 447968 81854 478338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 447968 85574 482058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 447968 92414 452898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 447968 96134 456618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 447968 99854 460338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 447968 103574 464058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 447968 110414 470898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 447968 114134 474618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 447968 117854 478338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 447968 121574 482058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 447968 128414 452898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 447968 132134 456618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 447968 135854 460338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 447968 139574 464058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 447968 146414 470898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 447968 150134 474618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 447968 153854 478338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 447968 157574 482058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 447968 164414 452898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 447968 168134 456618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 447968 171854 460338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 447968 175574 464058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 447968 182414 470898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 447968 186134 474618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 447968 189854 478338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 447968 193574 482058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 447968 200414 452898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 447968 204134 456618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 447968 207854 460338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 447968 211574 464058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 447968 218414 470898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 447968 222134 474618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 447968 225854 478338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 447968 229574 482058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 447968 236414 452898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 447968 240134 456618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 447968 243854 460338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 447968 247574 464058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 447968 254414 470898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 447968 258134 474618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 447968 261854 478338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 447968 265574 482058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 447968 272414 452898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 447968 276134 456618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 447968 279854 460338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 447968 283574 464058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 447968 290414 470898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 447968 294134 474618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 447968 297854 478338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 447968 301574 482058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 447968 308414 452898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 447968 312134 456618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 447968 315854 460338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 447968 319574 464058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 447968 326414 470898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 447968 330134 474618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 447968 333854 478338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 447968 337574 482058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 447968 344414 452898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 447968 348134 456618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 447968 351854 460338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 447968 355574 464058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 447968 362414 470898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 447968 366134 474618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 447968 369854 478338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 447968 373574 482058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 447968 380414 452898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 447968 384134 456618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 447968 387854 460338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 447968 391574 464058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 447968 398414 470898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 447968 402134 474618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 447968 405854 478338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 447968 409574 482058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 447968 416414 452898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 447968 420134 456618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 447968 423854 460338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 447968 427574 464058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 447968 434414 470898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 447968 438134 474618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 447968 441854 478338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 447968 445574 482058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 447968 452414 452898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 447968 456134 456618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 447968 459854 460338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 447968 463574 464058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 291883 59804 291949 59805
rect 291883 59740 291884 59804
rect 291948 59740 291949 59804
rect 291883 59739 291949 59740
rect 180747 59396 180813 59397
rect 180747 59332 180748 59396
rect 180812 59332 180813 59396
rect 180747 59331 180813 59332
rect 180750 59125 180810 59331
rect 180747 59124 180813 59125
rect 180747 59060 180748 59124
rect 180812 59060 180813 59124
rect 180747 59059 180813 59060
rect 291886 58989 291946 59739
rect 291883 58988 291949 58989
rect 291883 58924 291884 58988
rect 291948 58924 291949 58988
rect 291883 58923 291949 58924
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 58000
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 28894 63854 58000
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 32614 67574 58000
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 39454 74414 58000
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 43174 78134 58000
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 46894 81854 58000
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 50614 85574 58000
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 58000
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 58000
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 28894 99854 58000
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 32614 103574 58000
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 39454 110414 58000
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 43174 114134 58000
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 46894 117854 58000
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 50614 121574 58000
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 58000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 58000
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 28894 135854 58000
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 32614 139574 58000
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 39454 146414 58000
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 43174 150134 58000
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 46894 153854 58000
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 50614 157574 58000
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 57454 164414 58000
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 25174 168134 58000
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 28894 171854 58000
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 32614 175574 58000
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 39454 182414 58000
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 43174 186134 58000
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 46894 189854 58000
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 50614 193574 58000
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 57454 200414 58000
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 58000
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 28894 207854 58000
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 32614 211574 58000
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 39454 218414 58000
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 43174 222134 58000
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 46894 225854 58000
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 50614 229574 58000
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 57454 236414 58000
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 58000
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 28894 243854 58000
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 32614 247574 58000
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 39454 254414 58000
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 43174 258134 58000
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 46894 261854 58000
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 50614 265574 58000
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 57454 272414 58000
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 25174 276134 58000
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 28894 279854 58000
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 32614 283574 58000
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 39454 290414 58000
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 43174 294134 58000
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 46894 297854 58000
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 50614 301574 58000
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 57454 308414 58000
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 25174 312134 58000
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 28894 315854 58000
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 32614 319574 58000
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 39454 326414 58000
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 43174 330134 58000
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 46894 333854 58000
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 50614 337574 58000
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 57454 344414 58000
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 25174 348134 58000
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 28894 351854 58000
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 32614 355574 58000
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 39454 362414 58000
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 43174 366134 58000
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 46894 369854 58000
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 50614 373574 58000
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 57454 380414 58000
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 25174 384134 58000
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 28894 387854 58000
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 32614 391574 58000
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 39454 398414 58000
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 43174 402134 58000
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 46894 405854 58000
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 50614 409574 58000
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 57454 416414 58000
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 25174 420134 58000
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 28894 423854 58000
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 32614 427574 58000
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 39454 434414 58000
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 43174 438134 58000
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 46894 441854 58000
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 50614 445574 58000
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 57454 452414 58000
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 25174 456134 58000
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 28894 459854 58000
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 32614 463574 58000
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 58000 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 58000 446614
rect -8726 446294 58000 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 58000 446294
rect -8726 446026 58000 446058
rect 467996 446614 592650 446646
rect 467996 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect 467996 446294 592650 446378
rect 467996 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect 467996 446026 592650 446058
rect -6806 442894 58000 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 58000 442894
rect -6806 442574 58000 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 58000 442574
rect -6806 442306 58000 442338
rect 467996 442894 590730 442926
rect 467996 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect 467996 442574 590730 442658
rect 467996 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect 467996 442306 590730 442338
rect -4886 439174 58000 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 58000 439174
rect -4886 438854 58000 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 58000 438854
rect -4886 438586 58000 438618
rect 467996 439174 588810 439206
rect 467996 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect 467996 438854 588810 438938
rect 467996 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect 467996 438586 588810 438618
rect -2966 435454 58000 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 58000 435454
rect -2966 435134 58000 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 58000 435134
rect -2966 434866 58000 434898
rect 467996 435454 586890 435486
rect 467996 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect 467996 435134 586890 435218
rect 467996 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect 467996 434866 586890 434898
rect -8726 428614 58000 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 58000 428614
rect -8726 428294 58000 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 58000 428294
rect -8726 428026 58000 428058
rect 467996 428614 592650 428646
rect 467996 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 467996 428294 592650 428378
rect 467996 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 467996 428026 592650 428058
rect -6806 424894 58000 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 58000 424894
rect -6806 424574 58000 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 58000 424574
rect -6806 424306 58000 424338
rect 467996 424894 590730 424926
rect 467996 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 467996 424574 590730 424658
rect 467996 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 467996 424306 590730 424338
rect -4886 421174 58000 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 58000 421174
rect -4886 420854 58000 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 58000 420854
rect -4886 420586 58000 420618
rect 467996 421174 588810 421206
rect 467996 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 467996 420854 588810 420938
rect 467996 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 467996 420586 588810 420618
rect -2966 417454 58000 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 58000 417454
rect -2966 417134 58000 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 58000 417134
rect -2966 416866 58000 416898
rect 467996 417454 586890 417486
rect 467996 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 467996 417134 586890 417218
rect 467996 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 467996 416866 586890 416898
rect -8726 410614 58000 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 58000 410614
rect -8726 410294 58000 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 58000 410294
rect -8726 410026 58000 410058
rect 467996 410614 592650 410646
rect 467996 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect 467996 410294 592650 410378
rect 467996 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect 467996 410026 592650 410058
rect -6806 406894 58000 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 58000 406894
rect -6806 406574 58000 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 58000 406574
rect -6806 406306 58000 406338
rect 467996 406894 590730 406926
rect 467996 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect 467996 406574 590730 406658
rect 467996 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect 467996 406306 590730 406338
rect -4886 403174 58000 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 58000 403174
rect -4886 402854 58000 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 58000 402854
rect -4886 402586 58000 402618
rect 467996 403174 588810 403206
rect 467996 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect 467996 402854 588810 402938
rect 467996 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect 467996 402586 588810 402618
rect -2966 399454 58000 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 58000 399454
rect -2966 399134 58000 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 58000 399134
rect -2966 398866 58000 398898
rect 467996 399454 586890 399486
rect 467996 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect 467996 399134 586890 399218
rect 467996 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect 467996 398866 586890 398898
rect -8726 392614 58000 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 58000 392614
rect -8726 392294 58000 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 58000 392294
rect -8726 392026 58000 392058
rect 467996 392614 592650 392646
rect 467996 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 467996 392294 592650 392378
rect 467996 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 467996 392026 592650 392058
rect -6806 388894 58000 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 58000 388894
rect -6806 388574 58000 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 58000 388574
rect -6806 388306 58000 388338
rect 467996 388894 590730 388926
rect 467996 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 467996 388574 590730 388658
rect 467996 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 467996 388306 590730 388338
rect -4886 385174 58000 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 58000 385174
rect -4886 384854 58000 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 58000 384854
rect -4886 384586 58000 384618
rect 467996 385174 588810 385206
rect 467996 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 467996 384854 588810 384938
rect 467996 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 467996 384586 588810 384618
rect -2966 381454 58000 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 58000 381454
rect -2966 381134 58000 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 58000 381134
rect -2966 380866 58000 380898
rect 467996 381454 586890 381486
rect 467996 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 467996 381134 586890 381218
rect 467996 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 467996 380866 586890 380898
rect -8726 374614 58000 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 58000 374614
rect -8726 374294 58000 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 58000 374294
rect -8726 374026 58000 374058
rect 467996 374614 592650 374646
rect 467996 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect 467996 374294 592650 374378
rect 467996 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect 467996 374026 592650 374058
rect -6806 370894 58000 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 58000 370894
rect -6806 370574 58000 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 58000 370574
rect -6806 370306 58000 370338
rect 467996 370894 590730 370926
rect 467996 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect 467996 370574 590730 370658
rect 467996 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect 467996 370306 590730 370338
rect -4886 367174 58000 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 58000 367174
rect -4886 366854 58000 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 58000 366854
rect -4886 366586 58000 366618
rect 467996 367174 588810 367206
rect 467996 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect 467996 366854 588810 366938
rect 467996 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect 467996 366586 588810 366618
rect -2966 363454 58000 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 58000 363454
rect -2966 363134 58000 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 58000 363134
rect -2966 362866 58000 362898
rect 467996 363454 586890 363486
rect 467996 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect 467996 363134 586890 363218
rect 467996 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect 467996 362866 586890 362898
rect -8726 356614 58000 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 58000 356614
rect -8726 356294 58000 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 58000 356294
rect -8726 356026 58000 356058
rect 467996 356614 592650 356646
rect 467996 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 467996 356294 592650 356378
rect 467996 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 467996 356026 592650 356058
rect -6806 352894 58000 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 58000 352894
rect -6806 352574 58000 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 58000 352574
rect -6806 352306 58000 352338
rect 467996 352894 590730 352926
rect 467996 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 467996 352574 590730 352658
rect 467996 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 467996 352306 590730 352338
rect -4886 349174 58000 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 58000 349174
rect -4886 348854 58000 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 58000 348854
rect -4886 348586 58000 348618
rect 467996 349174 588810 349206
rect 467996 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 467996 348854 588810 348938
rect 467996 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 467996 348586 588810 348618
rect -2966 345454 58000 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 58000 345454
rect -2966 345134 58000 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 58000 345134
rect -2966 344866 58000 344898
rect 467996 345454 586890 345486
rect 467996 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 467996 345134 586890 345218
rect 467996 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 467996 344866 586890 344898
rect -8726 338614 58000 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 58000 338614
rect -8726 338294 58000 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 58000 338294
rect -8726 338026 58000 338058
rect 467996 338614 592650 338646
rect 467996 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect 467996 338294 592650 338378
rect 467996 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect 467996 338026 592650 338058
rect -6806 334894 58000 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 58000 334894
rect -6806 334574 58000 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 58000 334574
rect -6806 334306 58000 334338
rect 467996 334894 590730 334926
rect 467996 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect 467996 334574 590730 334658
rect 467996 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect 467996 334306 590730 334338
rect -4886 331174 58000 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 58000 331174
rect -4886 330854 58000 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 58000 330854
rect -4886 330586 58000 330618
rect 467996 331174 588810 331206
rect 467996 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect 467996 330854 588810 330938
rect 467996 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect 467996 330586 588810 330618
rect -2966 327454 58000 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 58000 327454
rect -2966 327134 58000 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 58000 327134
rect -2966 326866 58000 326898
rect 467996 327454 586890 327486
rect 467996 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect 467996 327134 586890 327218
rect 467996 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect 467996 326866 586890 326898
rect -8726 320614 58000 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 58000 320614
rect -8726 320294 58000 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 58000 320294
rect -8726 320026 58000 320058
rect 467996 320614 592650 320646
rect 467996 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 467996 320294 592650 320378
rect 467996 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 467996 320026 592650 320058
rect -6806 316894 58000 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 58000 316894
rect -6806 316574 58000 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 58000 316574
rect -6806 316306 58000 316338
rect 467996 316894 590730 316926
rect 467996 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 467996 316574 590730 316658
rect 467996 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 467996 316306 590730 316338
rect -4886 313174 58000 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 58000 313174
rect -4886 312854 58000 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 58000 312854
rect -4886 312586 58000 312618
rect 467996 313174 588810 313206
rect 467996 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 467996 312854 588810 312938
rect 467996 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 467996 312586 588810 312618
rect -2966 309454 58000 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 58000 309454
rect -2966 309134 58000 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 58000 309134
rect -2966 308866 58000 308898
rect 467996 309454 586890 309486
rect 467996 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 467996 309134 586890 309218
rect 467996 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 467996 308866 586890 308898
rect -8726 302614 58000 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 58000 302614
rect -8726 302294 58000 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 58000 302294
rect -8726 302026 58000 302058
rect 467996 302614 592650 302646
rect 467996 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect 467996 302294 592650 302378
rect 467996 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect 467996 302026 592650 302058
rect -6806 298894 58000 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 58000 298894
rect -6806 298574 58000 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 58000 298574
rect -6806 298306 58000 298338
rect 467996 298894 590730 298926
rect 467996 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect 467996 298574 590730 298658
rect 467996 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect 467996 298306 590730 298338
rect -4886 295174 58000 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 58000 295174
rect -4886 294854 58000 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 58000 294854
rect -4886 294586 58000 294618
rect 467996 295174 588810 295206
rect 467996 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect 467996 294854 588810 294938
rect 467996 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect 467996 294586 588810 294618
rect -2966 291454 58000 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 58000 291454
rect -2966 291134 58000 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 58000 291134
rect -2966 290866 58000 290898
rect 467996 291454 586890 291486
rect 467996 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect 467996 291134 586890 291218
rect 467996 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect 467996 290866 586890 290898
rect -8726 284614 58000 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 58000 284614
rect -8726 284294 58000 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 58000 284294
rect -8726 284026 58000 284058
rect 467996 284614 592650 284646
rect 467996 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 467996 284294 592650 284378
rect 467996 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 467996 284026 592650 284058
rect -6806 280894 58000 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 58000 280894
rect -6806 280574 58000 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 58000 280574
rect -6806 280306 58000 280338
rect 467996 280894 590730 280926
rect 467996 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 467996 280574 590730 280658
rect 467996 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 467996 280306 590730 280338
rect -4886 277174 58000 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 58000 277174
rect -4886 276854 58000 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 58000 276854
rect -4886 276586 58000 276618
rect 467996 277174 588810 277206
rect 467996 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 467996 276854 588810 276938
rect 467996 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 467996 276586 588810 276618
rect -2966 273454 58000 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 58000 273454
rect -2966 273134 58000 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 58000 273134
rect -2966 272866 58000 272898
rect 467996 273454 586890 273486
rect 467996 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 467996 273134 586890 273218
rect 467996 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 467996 272866 586890 272898
rect -8726 266614 58000 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 58000 266614
rect -8726 266294 58000 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 58000 266294
rect -8726 266026 58000 266058
rect 467996 266614 592650 266646
rect 467996 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect 467996 266294 592650 266378
rect 467996 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect 467996 266026 592650 266058
rect -6806 262894 58000 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 58000 262894
rect -6806 262574 58000 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 58000 262574
rect -6806 262306 58000 262338
rect 467996 262894 590730 262926
rect 467996 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect 467996 262574 590730 262658
rect 467996 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect 467996 262306 590730 262338
rect -4886 259174 58000 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 58000 259174
rect -4886 258854 58000 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 58000 258854
rect -4886 258586 58000 258618
rect 467996 259174 588810 259206
rect 467996 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect 467996 258854 588810 258938
rect 467996 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect 467996 258586 588810 258618
rect -2966 255454 58000 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 58000 255454
rect -2966 255134 58000 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 58000 255134
rect -2966 254866 58000 254898
rect 467996 255454 586890 255486
rect 467996 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect 467996 255134 586890 255218
rect 467996 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect 467996 254866 586890 254898
rect -8726 248614 58000 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 58000 248614
rect -8726 248294 58000 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 58000 248294
rect -8726 248026 58000 248058
rect 467996 248614 592650 248646
rect 467996 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 467996 248294 592650 248378
rect 467996 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 467996 248026 592650 248058
rect -6806 244894 58000 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 58000 244894
rect -6806 244574 58000 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 58000 244574
rect -6806 244306 58000 244338
rect 467996 244894 590730 244926
rect 467996 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 467996 244574 590730 244658
rect 467996 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 467996 244306 590730 244338
rect -4886 241174 58000 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 58000 241174
rect -4886 240854 58000 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 58000 240854
rect -4886 240586 58000 240618
rect 467996 241174 588810 241206
rect 467996 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 467996 240854 588810 240938
rect 467996 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 467996 240586 588810 240618
rect -2966 237454 58000 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 58000 237454
rect -2966 237134 58000 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 58000 237134
rect -2966 236866 58000 236898
rect 467996 237454 586890 237486
rect 467996 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 467996 237134 586890 237218
rect 467996 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 467996 236866 586890 236898
rect -8726 230614 58000 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 58000 230614
rect -8726 230294 58000 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 58000 230294
rect -8726 230026 58000 230058
rect 467996 230614 592650 230646
rect 467996 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect 467996 230294 592650 230378
rect 467996 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect 467996 230026 592650 230058
rect -6806 226894 58000 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 58000 226894
rect -6806 226574 58000 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 58000 226574
rect -6806 226306 58000 226338
rect 467996 226894 590730 226926
rect 467996 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect 467996 226574 590730 226658
rect 467996 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect 467996 226306 590730 226338
rect -4886 223174 58000 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 58000 223174
rect -4886 222854 58000 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 58000 222854
rect -4886 222586 58000 222618
rect 467996 223174 588810 223206
rect 467996 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect 467996 222854 588810 222938
rect 467996 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect 467996 222586 588810 222618
rect -2966 219454 58000 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 58000 219454
rect -2966 219134 58000 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 58000 219134
rect -2966 218866 58000 218898
rect 467996 219454 586890 219486
rect 467996 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect 467996 219134 586890 219218
rect 467996 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect 467996 218866 586890 218898
rect -8726 212614 58000 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 58000 212614
rect -8726 212294 58000 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 58000 212294
rect -8726 212026 58000 212058
rect 467996 212614 592650 212646
rect 467996 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 467996 212294 592650 212378
rect 467996 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 467996 212026 592650 212058
rect -6806 208894 58000 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 58000 208894
rect -6806 208574 58000 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 58000 208574
rect -6806 208306 58000 208338
rect 467996 208894 590730 208926
rect 467996 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 467996 208574 590730 208658
rect 467996 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 467996 208306 590730 208338
rect -4886 205174 58000 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 58000 205174
rect -4886 204854 58000 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 58000 204854
rect -4886 204586 58000 204618
rect 467996 205174 588810 205206
rect 467996 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 467996 204854 588810 204938
rect 467996 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 467996 204586 588810 204618
rect -2966 201454 58000 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 58000 201454
rect -2966 201134 58000 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 58000 201134
rect -2966 200866 58000 200898
rect 467996 201454 586890 201486
rect 467996 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 467996 201134 586890 201218
rect 467996 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 467996 200866 586890 200898
rect -8726 194614 58000 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 58000 194614
rect -8726 194294 58000 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 58000 194294
rect -8726 194026 58000 194058
rect 467996 194614 592650 194646
rect 467996 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect 467996 194294 592650 194378
rect 467996 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect 467996 194026 592650 194058
rect -6806 190894 58000 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 58000 190894
rect -6806 190574 58000 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 58000 190574
rect -6806 190306 58000 190338
rect 467996 190894 590730 190926
rect 467996 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect 467996 190574 590730 190658
rect 467996 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect 467996 190306 590730 190338
rect -4886 187174 58000 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 58000 187174
rect -4886 186854 58000 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 58000 186854
rect -4886 186586 58000 186618
rect 467996 187174 588810 187206
rect 467996 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect 467996 186854 588810 186938
rect 467996 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect 467996 186586 588810 186618
rect -2966 183454 58000 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 58000 183454
rect -2966 183134 58000 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 58000 183134
rect -2966 182866 58000 182898
rect 467996 183454 586890 183486
rect 467996 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect 467996 183134 586890 183218
rect 467996 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect 467996 182866 586890 182898
rect -8726 176614 58000 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 58000 176614
rect -8726 176294 58000 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 58000 176294
rect -8726 176026 58000 176058
rect 467996 176614 592650 176646
rect 467996 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 467996 176294 592650 176378
rect 467996 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 467996 176026 592650 176058
rect -6806 172894 58000 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 58000 172894
rect -6806 172574 58000 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 58000 172574
rect -6806 172306 58000 172338
rect 467996 172894 590730 172926
rect 467996 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 467996 172574 590730 172658
rect 467996 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 467996 172306 590730 172338
rect -4886 169174 58000 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 58000 169174
rect -4886 168854 58000 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 58000 168854
rect -4886 168586 58000 168618
rect 467996 169174 588810 169206
rect 467996 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 467996 168854 588810 168938
rect 467996 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 467996 168586 588810 168618
rect -2966 165454 58000 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 58000 165454
rect -2966 165134 58000 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 58000 165134
rect -2966 164866 58000 164898
rect 467996 165454 586890 165486
rect 467996 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 467996 165134 586890 165218
rect 467996 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 467996 164866 586890 164898
rect -8726 158614 58000 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 58000 158614
rect -8726 158294 58000 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 58000 158294
rect -8726 158026 58000 158058
rect 467996 158614 592650 158646
rect 467996 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect 467996 158294 592650 158378
rect 467996 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect 467996 158026 592650 158058
rect -6806 154894 58000 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 58000 154894
rect -6806 154574 58000 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 58000 154574
rect -6806 154306 58000 154338
rect 467996 154894 590730 154926
rect 467996 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect 467996 154574 590730 154658
rect 467996 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect 467996 154306 590730 154338
rect -4886 151174 58000 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 58000 151174
rect -4886 150854 58000 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 58000 150854
rect -4886 150586 58000 150618
rect 467996 151174 588810 151206
rect 467996 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect 467996 150854 588810 150938
rect 467996 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect 467996 150586 588810 150618
rect -2966 147454 58000 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 58000 147454
rect -2966 147134 58000 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 58000 147134
rect -2966 146866 58000 146898
rect 467996 147454 586890 147486
rect 467996 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect 467996 147134 586890 147218
rect 467996 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect 467996 146866 586890 146898
rect -8726 140614 58000 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 58000 140614
rect -8726 140294 58000 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 58000 140294
rect -8726 140026 58000 140058
rect 467996 140614 592650 140646
rect 467996 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 467996 140294 592650 140378
rect 467996 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 467996 140026 592650 140058
rect -6806 136894 58000 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 58000 136894
rect -6806 136574 58000 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 58000 136574
rect -6806 136306 58000 136338
rect 467996 136894 590730 136926
rect 467996 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 467996 136574 590730 136658
rect 467996 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 467996 136306 590730 136338
rect -4886 133174 58000 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 58000 133174
rect -4886 132854 58000 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 58000 132854
rect -4886 132586 58000 132618
rect 467996 133174 588810 133206
rect 467996 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 467996 132854 588810 132938
rect 467996 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 467996 132586 588810 132618
rect -2966 129454 58000 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 58000 129454
rect -2966 129134 58000 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 58000 129134
rect -2966 128866 58000 128898
rect 467996 129454 586890 129486
rect 467996 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 467996 129134 586890 129218
rect 467996 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 467996 128866 586890 128898
rect -8726 122614 58000 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 58000 122614
rect -8726 122294 58000 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 58000 122294
rect -8726 122026 58000 122058
rect 467996 122614 592650 122646
rect 467996 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect 467996 122294 592650 122378
rect 467996 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect 467996 122026 592650 122058
rect -6806 118894 58000 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 58000 118894
rect -6806 118574 58000 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 58000 118574
rect -6806 118306 58000 118338
rect 467996 118894 590730 118926
rect 467996 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect 467996 118574 590730 118658
rect 467996 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect 467996 118306 590730 118338
rect -4886 115174 58000 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 58000 115174
rect -4886 114854 58000 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 58000 114854
rect -4886 114586 58000 114618
rect 467996 115174 588810 115206
rect 467996 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect 467996 114854 588810 114938
rect 467996 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect 467996 114586 588810 114618
rect -2966 111454 58000 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 58000 111454
rect -2966 111134 58000 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 58000 111134
rect -2966 110866 58000 110898
rect 467996 111454 586890 111486
rect 467996 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect 467996 111134 586890 111218
rect 467996 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect 467996 110866 586890 110898
rect -8726 104614 58000 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 58000 104614
rect -8726 104294 58000 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 58000 104294
rect -8726 104026 58000 104058
rect 467996 104614 592650 104646
rect 467996 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 467996 104294 592650 104378
rect 467996 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 467996 104026 592650 104058
rect -6806 100894 58000 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 58000 100894
rect -6806 100574 58000 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 58000 100574
rect -6806 100306 58000 100338
rect 467996 100894 590730 100926
rect 467996 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 467996 100574 590730 100658
rect 467996 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 467996 100306 590730 100338
rect -4886 97174 58000 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 58000 97174
rect -4886 96854 58000 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 58000 96854
rect -4886 96586 58000 96618
rect 467996 97174 588810 97206
rect 467996 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 467996 96854 588810 96938
rect 467996 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 467996 96586 588810 96618
rect -2966 93454 58000 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 58000 93454
rect -2966 93134 58000 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 58000 93134
rect -2966 92866 58000 92898
rect 467996 93454 586890 93486
rect 467996 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 467996 93134 586890 93218
rect 467996 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 467996 92866 586890 92898
rect -8726 86614 58000 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 58000 86614
rect -8726 86294 58000 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 58000 86294
rect -8726 86026 58000 86058
rect 467996 86614 592650 86646
rect 467996 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect 467996 86294 592650 86378
rect 467996 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect 467996 86026 592650 86058
rect -6806 82894 58000 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 58000 82894
rect -6806 82574 58000 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 58000 82574
rect -6806 82306 58000 82338
rect 467996 82894 590730 82926
rect 467996 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect 467996 82574 590730 82658
rect 467996 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect 467996 82306 590730 82338
rect -4886 79174 58000 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 58000 79174
rect -4886 78854 58000 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 58000 78854
rect -4886 78586 58000 78618
rect 467996 79174 588810 79206
rect 467996 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect 467996 78854 588810 78938
rect 467996 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect 467996 78586 588810 78618
rect -2966 75454 58000 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 58000 75454
rect -2966 75134 58000 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 58000 75134
rect -2966 74866 58000 74898
rect 467996 75454 586890 75486
rect 467996 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect 467996 75134 586890 75218
rect 467996 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect 467996 74866 586890 74898
rect -8726 68614 58000 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 58000 68614
rect -8726 68294 58000 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 58000 68294
rect -8726 68026 58000 68058
rect 467996 68614 592650 68646
rect 467996 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 467996 68294 592650 68378
rect 467996 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 467996 68026 592650 68058
rect -6806 64894 58000 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 58000 64894
rect -6806 64574 58000 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 58000 64574
rect -6806 64306 58000 64338
rect 467996 64894 590730 64926
rect 467996 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 467996 64574 590730 64658
rect 467996 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 467996 64306 590730 64338
rect -4886 61174 58000 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 58000 61174
rect -4886 60854 58000 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 58000 60854
rect -4886 60586 58000 60618
rect 467996 61174 588810 61206
rect 467996 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 467996 60854 588810 60938
rect 467996 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 467996 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use azadi_soc_top_caravel  mprj
timestamp 0
transform 1 0 60000 0 1 60000
box 0 0 405996 385968
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 58000 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s 467996 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 58000 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s 467996 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 58000 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s 467996 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 58000 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s 467996 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 58000 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s 467996 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 58000 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s 467996 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 58000 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s 467996 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 58000 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s 467996 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 58000 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s 467996 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 58000 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s 467996 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 58000 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s 467996 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 447968 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 447968 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 447968 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 447968 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 447968 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 447968 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 447968 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 447968 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 447968 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 447968 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 447968 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 58000 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s 467996 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 58000 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s 467996 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 58000 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s 467996 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 58000 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s 467996 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 58000 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s 467996 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 58000 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s 467996 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 58000 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s 467996 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 58000 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s 467996 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 58000 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s 467996 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 58000 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s 467996 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 58000 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s 467996 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 447968 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 447968 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 447968 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 447968 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 447968 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 447968 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 447968 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 447968 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 447968 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 447968 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 447968 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 58000 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s 467996 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 58000 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s 467996 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 58000 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s 467996 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 58000 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s 467996 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 58000 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s 467996 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 58000 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s 467996 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 58000 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s 467996 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 58000 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s 467996 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 58000 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s 467996 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 58000 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s 467996 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 58000 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s 467996 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 447968 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 447968 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 447968 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 447968 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 447968 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 447968 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 447968 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 447968 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 447968 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 447968 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 447968 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 58000 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s 467996 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 58000 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s 467996 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 58000 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s 467996 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 58000 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s 467996 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 58000 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s 467996 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 58000 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s 467996 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 58000 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s 467996 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 58000 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s 467996 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 58000 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s 467996 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 58000 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s 467996 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 58000 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s 467996 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 447968 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 447968 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 447968 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 447968 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 447968 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 447968 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 447968 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 447968 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 447968 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 447968 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 447968 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 58000 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 467996 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 58000 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 467996 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 58000 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 467996 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 58000 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 467996 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 58000 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 467996 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 58000 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 467996 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 58000 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 467996 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 58000 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 467996 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 58000 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 467996 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 58000 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 467996 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 58000 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 467996 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 447968 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 447968 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 447968 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 447968 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 447968 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 447968 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 447968 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 447968 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 447968 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 447968 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 447968 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 447968 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 58000 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 467996 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 58000 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 467996 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 58000 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 467996 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 58000 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 467996 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 58000 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 467996 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 58000 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 467996 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 58000 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 467996 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 58000 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 467996 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 58000 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 467996 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 58000 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 467996 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 58000 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 467996 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 447968 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 447968 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 447968 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 447968 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 447968 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 447968 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 447968 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 447968 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 447968 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 447968 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 447968 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 447968 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 58000 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 467996 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 58000 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 467996 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 58000 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 467996 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 58000 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 467996 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 58000 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 467996 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 58000 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 467996 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 58000 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 467996 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 58000 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 467996 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 58000 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 467996 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 58000 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 467996 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 447968 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 447968 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 447968 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 447968 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 447968 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 447968 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 447968 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 447968 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 447968 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 447968 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 447968 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 58000 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 467996 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 58000 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 467996 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 58000 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 467996 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 58000 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 467996 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 58000 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 467996 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 58000 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 467996 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 58000 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 467996 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 58000 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 467996 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 58000 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 467996 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 58000 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 467996 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 58000 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 467996 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 447968 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 447968 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 447968 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 447968 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 447968 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 447968 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 447968 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 447968 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 447968 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 447968 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 447968 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 447968 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
