magic
tech sky130A
magscale 1 2
timestamp 1653833104
<< metal1 >>
rect 256602 49784 256608 49836
rect 256660 49824 256666 49836
rect 257798 49824 257804 49836
rect 256660 49796 257804 49824
rect 256660 49784 256666 49796
rect 257798 49784 257804 49796
rect 257856 49784 257862 49836
rect 351822 49784 351828 49836
rect 351880 49824 351886 49836
rect 353294 49824 353300 49836
rect 351880 49796 353300 49824
rect 351880 49784 351886 49796
rect 353294 49784 353300 49796
rect 353352 49784 353358 49836
rect 3418 49716 3424 49768
rect 3476 49756 3482 49768
rect 97994 49756 98000 49768
rect 3476 49728 98000 49756
rect 3476 49716 3482 49728
rect 97994 49716 98000 49728
rect 98052 49716 98058 49768
rect 299474 49240 299480 49292
rect 299532 49280 299538 49292
rect 375374 49280 375380 49292
rect 299532 49252 375380 49280
rect 299532 49240 299538 49252
rect 375374 49240 375380 49252
rect 375432 49240 375438 49292
rect 436462 49240 436468 49292
rect 436520 49280 436526 49292
rect 520274 49280 520280 49292
rect 436520 49252 520280 49280
rect 436520 49240 436526 49252
rect 520274 49240 520280 49252
rect 520332 49240 520338 49292
rect 150434 49172 150440 49224
rect 150492 49212 150498 49224
rect 208118 49212 208124 49224
rect 150492 49184 208124 49212
rect 150492 49172 150498 49184
rect 208118 49172 208124 49184
rect 208176 49172 208182 49224
rect 282730 49172 282736 49224
rect 282788 49212 282794 49224
rect 412634 49212 412640 49224
rect 282788 49184 412640 49212
rect 282788 49172 282794 49184
rect 412634 49172 412640 49184
rect 412692 49172 412698 49224
rect 78674 49104 78680 49156
rect 78732 49144 78738 49156
rect 118602 49144 118608 49156
rect 78732 49116 118608 49144
rect 78732 49104 78738 49116
rect 118602 49104 118608 49116
rect 118660 49104 118666 49156
rect 197354 49104 197360 49156
rect 197412 49144 197418 49156
rect 346394 49144 346400 49156
rect 197412 49116 346400 49144
rect 197412 49104 197418 49116
rect 346394 49104 346400 49116
rect 346452 49104 346458 49156
rect 378778 49104 378784 49156
rect 378836 49144 378842 49156
rect 517698 49144 517704 49156
rect 378836 49116 517704 49144
rect 378836 49104 378842 49116
rect 517698 49104 517704 49116
rect 517756 49104 517762 49156
rect 92474 49036 92480 49088
rect 92532 49076 92538 49088
rect 184842 49076 184848 49088
rect 92532 49048 184848 49076
rect 92532 49036 92538 49048
rect 184842 49036 184848 49048
rect 184900 49036 184906 49088
rect 246942 49036 246948 49088
rect 247000 49076 247006 49088
rect 281534 49076 281540 49088
rect 247000 49048 281540 49076
rect 247000 49036 247006 49048
rect 281534 49036 281540 49048
rect 281592 49036 281598 49088
rect 311710 49036 311716 49088
rect 311768 49076 311774 49088
rect 518894 49076 518900 49088
rect 311768 49048 518900 49076
rect 311768 49036 311774 49048
rect 518894 49036 518900 49048
rect 518952 49036 518958 49088
rect 6914 48968 6920 49020
rect 6972 49008 6978 49020
rect 99374 49008 99380 49020
rect 6972 48980 99380 49008
rect 6972 48968 6978 48980
rect 99374 48968 99380 48980
rect 99432 48968 99438 49020
rect 198734 48968 198740 49020
rect 198792 49008 198798 49020
rect 470594 49008 470600 49020
rect 198792 48980 470600 49008
rect 198792 48968 198798 48980
rect 470594 48968 470600 48980
rect 470652 48968 470658 49020
rect 521746 48968 521752 49020
rect 521804 49008 521810 49020
rect 560386 49008 560392 49020
rect 521804 48980 560392 49008
rect 521804 48968 521810 48980
rect 560386 48968 560392 48980
rect 560444 48968 560450 49020
rect 346394 47880 346400 47932
rect 346452 47920 346458 47932
rect 387794 47920 387800 47932
rect 346452 47892 387800 47920
rect 346452 47880 346458 47892
rect 387794 47880 387800 47892
rect 387852 47880 387858 47932
rect 276014 47812 276020 47864
rect 276072 47852 276078 47864
rect 368750 47852 368756 47864
rect 276072 47824 368756 47852
rect 276072 47812 276078 47824
rect 368750 47812 368756 47824
rect 368808 47812 368814 47864
rect 286318 47744 286324 47796
rect 286376 47784 286382 47796
rect 426434 47784 426440 47796
rect 286376 47756 426440 47784
rect 286376 47744 286382 47756
rect 426434 47744 426440 47756
rect 426492 47744 426498 47796
rect 434622 47744 434628 47796
rect 434680 47784 434686 47796
rect 502426 47784 502432 47796
rect 434680 47756 502432 47784
rect 434680 47744 434686 47756
rect 502426 47744 502432 47756
rect 502484 47744 502490 47796
rect 190454 47676 190460 47728
rect 190512 47716 190518 47728
rect 345014 47716 345020 47728
rect 190512 47688 345020 47716
rect 190512 47676 190518 47688
rect 345014 47676 345020 47688
rect 345072 47676 345078 47728
rect 382918 47676 382924 47728
rect 382976 47716 382982 47728
rect 519170 47716 519176 47728
rect 382976 47688 519176 47716
rect 382976 47676 382982 47688
rect 519170 47676 519176 47688
rect 519228 47676 519234 47728
rect 93854 47608 93860 47660
rect 93912 47648 93918 47660
rect 122466 47648 122472 47660
rect 93912 47620 122472 47648
rect 93912 47608 93918 47620
rect 122466 47608 122472 47620
rect 122524 47608 122530 47660
rect 200114 47608 200120 47660
rect 200172 47648 200178 47660
rect 221826 47648 221832 47660
rect 200172 47620 221832 47648
rect 200172 47608 200178 47620
rect 221826 47608 221832 47620
rect 221884 47608 221890 47660
rect 242710 47608 242716 47660
rect 242768 47648 242774 47660
rect 267734 47648 267740 47660
rect 242768 47620 267740 47648
rect 242768 47608 242774 47620
rect 267734 47608 267740 47620
rect 267792 47608 267798 47660
rect 304902 47608 304908 47660
rect 304960 47648 304966 47660
rect 494054 47648 494060 47660
rect 304960 47620 494060 47648
rect 304960 47608 304966 47620
rect 494054 47608 494060 47620
rect 494112 47608 494118 47660
rect 1394 47540 1400 47592
rect 1452 47580 1458 47592
rect 99650 47580 99656 47592
rect 1452 47552 99656 47580
rect 1452 47540 1458 47552
rect 99650 47540 99656 47552
rect 99708 47540 99714 47592
rect 138014 47540 138020 47592
rect 138072 47580 138078 47592
rect 454402 47580 454408 47592
rect 138072 47552 454408 47580
rect 138072 47540 138078 47552
rect 454402 47540 454408 47552
rect 454460 47540 454466 47592
rect 510614 47540 510620 47592
rect 510672 47580 510678 47592
rect 557626 47580 557632 47592
rect 510672 47552 557632 47580
rect 510672 47540 510678 47552
rect 557626 47540 557632 47552
rect 557684 47540 557690 47592
rect 396074 46928 396080 46980
rect 396132 46968 396138 46980
rect 402974 46968 402980 46980
rect 396132 46940 402980 46968
rect 396132 46928 396138 46940
rect 402974 46928 402980 46940
rect 403032 46928 403038 46980
rect 282914 46452 282920 46504
rect 282972 46492 282978 46504
rect 369854 46492 369860 46504
rect 282972 46464 369860 46492
rect 282972 46452 282978 46464
rect 369854 46452 369860 46464
rect 369912 46452 369918 46504
rect 277302 46384 277308 46436
rect 277360 46424 277366 46436
rect 405734 46424 405740 46436
rect 277360 46396 405740 46424
rect 277360 46384 277366 46396
rect 405734 46384 405740 46396
rect 405792 46384 405798 46436
rect 201494 46316 201500 46368
rect 201552 46356 201558 46368
rect 348142 46356 348148 46368
rect 201552 46328 348148 46356
rect 201552 46316 201558 46328
rect 348142 46316 348148 46328
rect 348200 46316 348206 46368
rect 371234 46316 371240 46368
rect 371292 46356 371298 46368
rect 394694 46356 394700 46368
rect 371292 46328 394700 46356
rect 371292 46316 371298 46328
rect 394694 46316 394700 46328
rect 394752 46316 394758 46368
rect 416682 46316 416688 46368
rect 416740 46356 416746 46368
rect 438854 46356 438860 46368
rect 416740 46328 438860 46356
rect 416740 46316 416746 46328
rect 438854 46316 438860 46328
rect 438912 46316 438918 46368
rect 445662 46316 445668 46368
rect 445720 46356 445726 46368
rect 540974 46356 540980 46368
rect 445720 46328 540980 46356
rect 445720 46316 445726 46328
rect 540974 46316 540980 46328
rect 541032 46316 541038 46368
rect 46934 46248 46940 46300
rect 46992 46288 46998 46300
rect 109034 46288 109040 46300
rect 46992 46260 109040 46288
rect 46992 46248 46998 46260
rect 109034 46248 109040 46260
rect 109092 46248 109098 46300
rect 246758 46248 246764 46300
rect 246816 46288 246822 46300
rect 284294 46288 284300 46300
rect 246816 46260 284300 46288
rect 246816 46248 246822 46260
rect 284294 46248 284300 46260
rect 284352 46248 284358 46300
rect 315942 46248 315948 46300
rect 316000 46288 316006 46300
rect 543734 46288 543740 46300
rect 316000 46260 543740 46288
rect 316000 46248 316006 46260
rect 543734 46248 543740 46260
rect 543792 46248 543798 46300
rect 80054 46180 80060 46232
rect 80112 46220 80118 46232
rect 150526 46220 150532 46232
rect 80112 46192 150532 46220
rect 80112 46180 80118 46192
rect 150526 46180 150532 46192
rect 150584 46180 150590 46232
rect 175274 46180 175280 46232
rect 175332 46220 175338 46232
rect 214926 46220 214932 46232
rect 175332 46192 214932 46220
rect 175332 46180 175338 46192
rect 214926 46180 214932 46192
rect 214984 46180 214990 46232
rect 253198 46180 253204 46232
rect 253256 46220 253262 46232
rect 484578 46220 484584 46232
rect 253256 46192 484584 46220
rect 253256 46180 253262 46192
rect 484578 46180 484584 46192
rect 484636 46180 484642 46232
rect 321554 45160 321560 45212
rect 321612 45200 321618 45212
rect 383930 45200 383936 45212
rect 321612 45172 383936 45200
rect 321612 45160 321618 45172
rect 383930 45160 383936 45172
rect 383988 45160 383994 45212
rect 278682 45092 278688 45144
rect 278740 45132 278746 45144
rect 408494 45132 408500 45144
rect 278740 45104 408500 45132
rect 278740 45092 278746 45104
rect 408494 45092 408500 45104
rect 408552 45092 408558 45144
rect 329098 45024 329104 45076
rect 329156 45064 329162 45076
rect 502334 45064 502340 45076
rect 329156 45036 502340 45064
rect 329156 45024 329162 45036
rect 502334 45024 502340 45036
rect 502392 45024 502398 45076
rect 297910 44956 297916 45008
rect 297968 44996 297974 45008
rect 476114 44996 476120 45008
rect 297968 44968 476120 44996
rect 297968 44956 297974 44968
rect 476114 44956 476120 44968
rect 476172 44956 476178 45008
rect 53834 44888 53840 44940
rect 53892 44928 53898 44940
rect 112622 44928 112628 44940
rect 53892 44900 112628 44928
rect 53892 44888 53898 44900
rect 112622 44888 112628 44900
rect 112680 44888 112686 44940
rect 154574 44888 154580 44940
rect 154632 44928 154638 44940
rect 333422 44928 333428 44940
rect 154632 44900 333428 44928
rect 154632 44888 154638 44900
rect 333422 44888 333428 44900
rect 333480 44888 333486 44940
rect 418890 44888 418896 44940
rect 418948 44928 418954 44940
rect 528554 44928 528560 44940
rect 418948 44900 528560 44928
rect 418948 44888 418954 44900
rect 528554 44888 528560 44900
rect 528612 44888 528618 44940
rect 93946 44820 93952 44872
rect 94004 44860 94010 44872
rect 155402 44860 155408 44872
rect 94004 44832 155408 44860
rect 94004 44820 94010 44832
rect 155402 44820 155408 44832
rect 155460 44820 155466 44872
rect 168374 44820 168380 44872
rect 168432 44860 168438 44872
rect 211798 44860 211804 44872
rect 168432 44832 211804 44860
rect 168432 44820 168438 44832
rect 211798 44820 211804 44832
rect 211856 44820 211862 44872
rect 248230 44820 248236 44872
rect 248288 44860 248294 44872
rect 295334 44860 295340 44872
rect 248288 44832 295340 44860
rect 248288 44820 248294 44832
rect 295334 44820 295340 44832
rect 295392 44820 295398 44872
rect 319990 44820 319996 44872
rect 320048 44860 320054 44872
rect 557534 44860 557540 44872
rect 320048 44832 557540 44860
rect 320048 44820 320054 44832
rect 557534 44820 557540 44832
rect 557592 44820 557598 44872
rect 310514 43732 310520 43784
rect 310572 43772 310578 43784
rect 380894 43772 380900 43784
rect 310572 43744 380900 43772
rect 310572 43732 310578 43744
rect 380894 43732 380900 43744
rect 380952 43732 380958 43784
rect 262122 43664 262128 43716
rect 262180 43704 262186 43716
rect 349154 43704 349160 43716
rect 262180 43676 349160 43704
rect 262180 43664 262186 43676
rect 349154 43664 349160 43676
rect 349212 43664 349218 43716
rect 286870 43596 286876 43648
rect 286928 43636 286934 43648
rect 440234 43636 440240 43648
rect 286928 43608 440240 43636
rect 286928 43596 286934 43608
rect 440234 43596 440240 43608
rect 440292 43596 440298 43648
rect 443638 43596 443644 43648
rect 443696 43636 443702 43648
rect 532694 43636 532700 43648
rect 443696 43608 532700 43636
rect 443696 43596 443702 43608
rect 532694 43596 532700 43608
rect 532752 43596 532758 43648
rect 129734 43528 129740 43580
rect 129792 43568 129798 43580
rect 326522 43568 326528 43580
rect 129792 43540 326528 43568
rect 129792 43528 129798 43540
rect 326522 43528 326528 43540
rect 326580 43528 326586 43580
rect 348418 43528 348424 43580
rect 348476 43568 348482 43580
rect 509326 43568 509332 43580
rect 348476 43540 509332 43568
rect 348476 43528 348482 43540
rect 509326 43528 509332 43540
rect 509384 43528 509390 43580
rect 60734 43460 60740 43512
rect 60792 43500 60798 43512
rect 113818 43500 113824 43512
rect 60792 43472 113824 43500
rect 60792 43460 60798 43472
rect 113818 43460 113824 43472
rect 113876 43460 113882 43512
rect 319806 43460 319812 43512
rect 319864 43500 319870 43512
rect 561674 43500 561680 43512
rect 319864 43472 561680 43500
rect 319864 43460 319870 43472
rect 561674 43460 561680 43472
rect 561732 43460 561738 43512
rect 67634 43392 67640 43444
rect 67692 43432 67698 43444
rect 177482 43432 177488 43444
rect 67692 43404 177488 43432
rect 67692 43392 67698 43404
rect 177482 43392 177488 43404
rect 177540 43392 177546 43444
rect 219434 43392 219440 43444
rect 219492 43432 219498 43444
rect 480346 43432 480352 43444
rect 219492 43404 480352 43432
rect 219492 43392 219498 43404
rect 480346 43392 480352 43404
rect 480404 43392 480410 43444
rect 307754 42372 307760 42424
rect 307812 42412 307818 42424
rect 379514 42412 379520 42424
rect 307812 42384 379520 42412
rect 307812 42372 307818 42384
rect 379514 42372 379520 42384
rect 379572 42372 379578 42424
rect 284018 42304 284024 42356
rect 284076 42344 284082 42356
rect 430574 42344 430580 42356
rect 284076 42316 430580 42344
rect 284076 42304 284082 42316
rect 430574 42304 430580 42316
rect 430632 42304 430638 42356
rect 204254 42236 204260 42288
rect 204312 42276 204318 42288
rect 352006 42276 352012 42288
rect 204312 42248 352012 42276
rect 204312 42236 204318 42248
rect 352006 42236 352012 42248
rect 352064 42236 352070 42288
rect 429930 42236 429936 42288
rect 429988 42276 429994 42288
rect 530210 42276 530216 42288
rect 429988 42248 530216 42276
rect 429988 42236 429994 42248
rect 530210 42236 530216 42248
rect 530268 42236 530274 42288
rect 64874 42168 64880 42220
rect 64932 42208 64938 42220
rect 115382 42208 115388 42220
rect 64932 42180 115388 42208
rect 64932 42168 64938 42180
rect 115382 42168 115388 42180
rect 115440 42168 115446 42220
rect 342898 42168 342904 42220
rect 342956 42208 342962 42220
rect 509510 42208 509516 42220
rect 342956 42180 509516 42208
rect 342956 42168 342962 42180
rect 509510 42168 509516 42180
rect 509568 42168 509574 42220
rect 106274 42100 106280 42152
rect 106332 42140 106338 42152
rect 188522 42140 188528 42152
rect 106332 42112 188528 42140
rect 106332 42100 106338 42112
rect 188522 42100 188528 42112
rect 188580 42100 188586 42152
rect 253750 42100 253756 42152
rect 253808 42140 253814 42152
rect 320174 42140 320180 42152
rect 253808 42112 320180 42140
rect 253808 42100 253814 42112
rect 320174 42100 320180 42112
rect 320232 42100 320238 42152
rect 321462 42100 321468 42152
rect 321520 42140 321526 42152
rect 564434 42140 564440 42152
rect 321520 42112 564440 42140
rect 321520 42100 321526 42112
rect 564434 42100 564440 42112
rect 564492 42100 564498 42152
rect 34514 42032 34520 42084
rect 34572 42072 34578 42084
rect 138842 42072 138848 42084
rect 34572 42044 138848 42072
rect 34572 42032 34578 42044
rect 138842 42032 138848 42044
rect 138900 42032 138906 42084
rect 194594 42032 194600 42084
rect 194652 42072 194658 42084
rect 473354 42072 473360 42084
rect 194652 42044 473360 42072
rect 194652 42032 194658 42044
rect 473354 42032 473360 42044
rect 473412 42032 473418 42084
rect 349246 41012 349252 41064
rect 349304 41052 349310 41064
rect 390738 41052 390744 41064
rect 349304 41024 390744 41052
rect 349304 41012 349310 41024
rect 390738 41012 390744 41024
rect 390796 41012 390802 41064
rect 264790 40944 264796 40996
rect 264848 40984 264854 40996
rect 358814 40984 358820 40996
rect 264848 40956 358820 40984
rect 264848 40944 264854 40956
rect 358814 40944 358820 40956
rect 358872 40944 358878 40996
rect 215294 40876 215300 40928
rect 215352 40916 215358 40928
rect 354858 40916 354864 40928
rect 215352 40888 354864 40916
rect 215352 40876 215358 40888
rect 354858 40876 354864 40888
rect 354916 40876 354922 40928
rect 376018 40876 376024 40928
rect 376076 40916 376082 40928
rect 516318 40916 516324 40928
rect 376076 40888 516324 40916
rect 376076 40876 376082 40888
rect 516318 40876 516324 40888
rect 516376 40876 516382 40928
rect 75914 40808 75920 40860
rect 75972 40848 75978 40860
rect 117958 40848 117964 40860
rect 75972 40820 117964 40848
rect 75972 40808 75978 40820
rect 117958 40808 117964 40820
rect 118016 40808 118022 40860
rect 289722 40808 289728 40860
rect 289780 40848 289786 40860
rect 448514 40848 448520 40860
rect 289780 40820 448520 40848
rect 289780 40808 289786 40820
rect 448514 40808 448520 40820
rect 448572 40808 448578 40860
rect 113174 40740 113180 40792
rect 113232 40780 113238 40792
rect 191282 40780 191288 40792
rect 113232 40752 191288 40780
rect 113232 40740 113238 40752
rect 191282 40740 191288 40752
rect 191340 40740 191346 40792
rect 318702 40740 318708 40792
rect 318760 40780 318766 40792
rect 554774 40780 554780 40792
rect 318760 40752 554780 40780
rect 318760 40740 318766 40752
rect 554774 40740 554780 40752
rect 554832 40740 554838 40792
rect 27614 40672 27620 40724
rect 27672 40712 27678 40724
rect 135898 40712 135904 40724
rect 27672 40684 135904 40712
rect 27672 40672 27678 40684
rect 135898 40672 135904 40684
rect 135956 40672 135962 40724
rect 241514 40672 241520 40724
rect 241572 40712 241578 40724
rect 485774 40712 485780 40724
rect 241572 40684 485780 40712
rect 241572 40672 241578 40684
rect 485774 40672 485780 40684
rect 485832 40672 485838 40724
rect 292574 39652 292580 39704
rect 292632 39692 292638 39704
rect 375374 39692 375380 39704
rect 292632 39664 375380 39692
rect 292632 39652 292638 39664
rect 375374 39652 375380 39664
rect 375432 39652 375438 39704
rect 277302 39584 277308 39636
rect 277360 39624 277366 39636
rect 401594 39624 401600 39636
rect 277360 39596 401600 39624
rect 277360 39584 277366 39596
rect 401594 39584 401600 39596
rect 401652 39584 401658 39636
rect 186314 39516 186320 39568
rect 186372 39556 186378 39568
rect 346486 39556 346492 39568
rect 186372 39528 346492 39556
rect 186372 39516 186378 39528
rect 346486 39516 346492 39528
rect 346544 39516 346550 39568
rect 403618 39516 403624 39568
rect 403676 39556 403682 39568
rect 523218 39556 523224 39568
rect 403676 39528 523224 39556
rect 403676 39516 403682 39528
rect 523218 39516 523224 39528
rect 523276 39516 523282 39568
rect 331950 39448 331956 39500
rect 332008 39488 332014 39500
rect 503898 39488 503904 39500
rect 332008 39460 503904 39488
rect 332008 39448 332014 39460
rect 503898 39448 503904 39460
rect 503956 39448 503962 39500
rect 85574 39380 85580 39432
rect 85632 39420 85638 39432
rect 120718 39420 120724 39432
rect 85632 39392 120724 39420
rect 85632 39380 85638 39392
rect 120718 39380 120724 39392
rect 120776 39380 120782 39432
rect 248046 39380 248052 39432
rect 248104 39420 248110 39432
rect 299566 39420 299572 39432
rect 248104 39392 299572 39420
rect 248104 39380 248110 39392
rect 299566 39380 299572 39392
rect 299624 39380 299630 39432
rect 317138 39380 317144 39432
rect 317196 39420 317202 39432
rect 550634 39420 550640 39432
rect 317196 39392 550640 39420
rect 317196 39380 317202 39392
rect 550634 39380 550640 39392
rect 550692 39380 550698 39432
rect 22094 39312 22100 39364
rect 22152 39352 22158 39364
rect 134702 39352 134708 39364
rect 22152 39324 134708 39352
rect 22152 39312 22158 39324
rect 134702 39312 134708 39324
rect 134760 39312 134766 39364
rect 191834 39312 191840 39364
rect 191892 39352 191898 39364
rect 471974 39352 471980 39364
rect 191892 39324 471980 39352
rect 191892 39312 191898 39324
rect 471974 39312 471980 39324
rect 472032 39312 472038 39364
rect 303614 38156 303620 38208
rect 303672 38196 303678 38208
rect 378318 38196 378324 38208
rect 303672 38168 378324 38196
rect 303672 38156 303678 38168
rect 378318 38156 378324 38168
rect 378376 38156 378382 38208
rect 281350 38088 281356 38140
rect 281408 38128 281414 38140
rect 415394 38128 415400 38140
rect 281408 38100 415400 38128
rect 281408 38088 281414 38100
rect 415394 38088 415400 38100
rect 415452 38088 415458 38140
rect 443730 38088 443736 38140
rect 443788 38128 443794 38140
rect 538214 38128 538220 38140
rect 443788 38100 538220 38128
rect 443788 38088 443794 38100
rect 538214 38088 538220 38100
rect 538272 38088 538278 38140
rect 193214 38020 193220 38072
rect 193272 38060 193278 38072
rect 347958 38060 347964 38072
rect 193272 38032 347964 38060
rect 193272 38020 193278 38032
rect 347958 38020 347964 38032
rect 348016 38020 348022 38072
rect 392578 38020 392584 38072
rect 392636 38060 392642 38072
rect 523034 38060 523040 38072
rect 392636 38032 523040 38060
rect 392636 38020 392642 38032
rect 523034 38020 523040 38032
rect 523092 38020 523098 38072
rect 89714 37952 89720 38004
rect 89772 37992 89778 38004
rect 122098 37992 122104 38004
rect 89772 37964 122104 37992
rect 89772 37952 89778 37964
rect 122098 37952 122104 37964
rect 122156 37952 122162 38004
rect 253566 37952 253572 38004
rect 253624 37992 253630 38004
rect 316034 37992 316040 38004
rect 253624 37964 316040 37992
rect 253624 37952 253630 37964
rect 316034 37952 316040 37964
rect 316092 37952 316098 38004
rect 317322 37952 317328 38004
rect 317380 37992 317386 38004
rect 547874 37992 547880 38004
rect 317380 37964 547880 37992
rect 317380 37952 317386 37964
rect 547874 37952 547880 37964
rect 547932 37952 547938 38004
rect 17954 37884 17960 37936
rect 18012 37924 18018 37936
rect 134518 37924 134524 37936
rect 18012 37896 134524 37924
rect 18012 37884 18018 37896
rect 134518 37884 134524 37896
rect 134576 37884 134582 37936
rect 244274 37884 244280 37936
rect 244332 37924 244338 37936
rect 487430 37924 487436 37936
rect 244332 37896 487436 37924
rect 244332 37884 244338 37896
rect 487430 37884 487436 37896
rect 487488 37884 487494 37936
rect 266262 36864 266268 36916
rect 266320 36904 266326 36916
rect 362954 36904 362960 36916
rect 266320 36876 362960 36904
rect 266320 36864 266326 36876
rect 362954 36864 362960 36876
rect 363012 36864 363018 36916
rect 240134 36796 240140 36848
rect 240192 36836 240198 36848
rect 361758 36836 361764 36848
rect 240192 36808 361764 36836
rect 240192 36796 240198 36808
rect 361758 36796 361764 36808
rect 361816 36796 361822 36848
rect 353938 36728 353944 36780
rect 353996 36768 354002 36780
rect 510706 36768 510712 36780
rect 353996 36740 510712 36768
rect 353996 36728 354002 36740
rect 510706 36728 510712 36740
rect 510764 36728 510770 36780
rect 77294 36660 77300 36712
rect 77352 36700 77358 36712
rect 149698 36700 149704 36712
rect 77352 36672 149704 36700
rect 77352 36660 77358 36672
rect 149698 36660 149704 36672
rect 149756 36660 149762 36712
rect 291010 36660 291016 36712
rect 291068 36700 291074 36712
rect 451274 36700 451280 36712
rect 291068 36672 451280 36700
rect 291068 36660 291074 36672
rect 451274 36660 451280 36672
rect 451332 36660 451338 36712
rect 99374 36592 99380 36644
rect 99432 36632 99438 36644
rect 186958 36632 186964 36644
rect 99432 36604 186964 36632
rect 99432 36592 99438 36604
rect 186958 36592 186964 36604
rect 187016 36592 187022 36644
rect 313182 36592 313188 36644
rect 313240 36632 313246 36644
rect 532694 36632 532700 36644
rect 313240 36604 532700 36632
rect 313240 36592 313246 36604
rect 532694 36592 532700 36604
rect 532752 36592 532758 36644
rect 16574 36524 16580 36576
rect 16632 36564 16638 36576
rect 101582 36564 101588 36576
rect 16632 36536 101588 36564
rect 16632 36524 16638 36536
rect 101582 36524 101588 36536
rect 101640 36524 101646 36576
rect 176654 36524 176660 36576
rect 176712 36564 176718 36576
rect 467834 36564 467840 36576
rect 176712 36536 467840 36564
rect 176712 36524 176718 36536
rect 467834 36524 467840 36536
rect 467892 36524 467898 36576
rect 267550 35504 267556 35556
rect 267608 35544 267614 35556
rect 369854 35544 369860 35556
rect 267608 35516 369860 35544
rect 267608 35504 267614 35516
rect 369854 35504 369860 35516
rect 369912 35504 369918 35556
rect 251174 35436 251180 35488
rect 251232 35476 251238 35488
rect 364426 35476 364432 35488
rect 251232 35448 364432 35476
rect 251232 35436 251238 35448
rect 364426 35436 364432 35448
rect 364484 35436 364490 35488
rect 360838 35368 360844 35420
rect 360896 35408 360902 35420
rect 513466 35408 513472 35420
rect 360896 35380 513472 35408
rect 360896 35368 360902 35380
rect 513466 35368 513472 35380
rect 513524 35368 513530 35420
rect 290826 35300 290832 35352
rect 290884 35340 290890 35352
rect 455414 35340 455420 35352
rect 290884 35312 455420 35340
rect 290884 35300 290890 35312
rect 455414 35300 455420 35312
rect 455472 35300 455478 35352
rect 86954 35232 86960 35284
rect 87012 35272 87018 35284
rect 152458 35272 152464 35284
rect 87012 35244 152464 35272
rect 87012 35232 87018 35244
rect 152458 35232 152464 35244
rect 152516 35232 152522 35284
rect 311802 35232 311808 35284
rect 311860 35272 311866 35284
rect 529934 35272 529940 35284
rect 311860 35244 529940 35272
rect 311860 35232 311866 35244
rect 529934 35232 529940 35244
rect 529992 35232 529998 35284
rect 20714 35164 20720 35216
rect 20772 35204 20778 35216
rect 102778 35204 102784 35216
rect 20772 35176 102784 35204
rect 20772 35164 20778 35176
rect 102778 35164 102784 35176
rect 102836 35164 102842 35216
rect 180794 35164 180800 35216
rect 180852 35204 180858 35216
rect 469214 35204 469220 35216
rect 180852 35176 469220 35204
rect 180852 35164 180858 35176
rect 469214 35164 469220 35176
rect 469272 35164 469278 35216
rect 273162 34008 273168 34060
rect 273220 34048 273226 34060
rect 387794 34048 387800 34060
rect 273220 34020 387800 34048
rect 273220 34008 273226 34020
rect 387794 34008 387800 34020
rect 387852 34008 387858 34060
rect 293770 33940 293776 33992
rect 293828 33980 293834 33992
rect 465074 33980 465080 33992
rect 293828 33952 465080 33980
rect 293828 33940 293834 33952
rect 465074 33940 465080 33952
rect 465132 33940 465138 33992
rect 133874 33872 133880 33924
rect 133932 33912 133938 33924
rect 326338 33912 326344 33924
rect 133932 33884 326344 33912
rect 133932 33872 133938 33884
rect 326338 33872 326344 33884
rect 326396 33872 326402 33924
rect 378870 33872 378876 33924
rect 378928 33912 378934 33924
rect 518986 33912 518992 33924
rect 378928 33884 518992 33912
rect 378928 33872 378934 33884
rect 518986 33872 518992 33884
rect 519044 33872 519050 33924
rect 28994 33804 29000 33856
rect 29052 33844 29058 33856
rect 105722 33844 105728 33856
rect 29052 33816 105728 33844
rect 29052 33804 29058 33816
rect 105722 33804 105728 33816
rect 105780 33804 105786 33856
rect 310238 33804 310244 33856
rect 310296 33844 310302 33856
rect 525794 33844 525800 33856
rect 310296 33816 525800 33844
rect 310296 33804 310302 33816
rect 525794 33804 525800 33816
rect 525852 33804 525858 33856
rect 56594 33736 56600 33788
rect 56652 33776 56658 33788
rect 174722 33776 174728 33788
rect 56652 33748 174728 33776
rect 56652 33736 56658 33748
rect 174722 33736 174728 33748
rect 174780 33736 174786 33788
rect 184934 33736 184940 33788
rect 184992 33776 184998 33788
rect 470686 33776 470692 33788
rect 184992 33748 470692 33776
rect 184992 33736 184998 33748
rect 470686 33736 470692 33748
rect 470744 33736 470750 33788
rect 524414 33736 524420 33788
rect 524472 33776 524478 33788
rect 563238 33776 563244 33788
rect 524472 33748 563244 33776
rect 524472 33736 524478 33748
rect 563238 33736 563244 33748
rect 563296 33736 563302 33788
rect 270218 32648 270224 32700
rect 270276 32688 270282 32700
rect 376754 32688 376760 32700
rect 270276 32660 376760 32688
rect 270276 32648 270282 32660
rect 376754 32648 376760 32660
rect 376812 32648 376818 32700
rect 445018 32648 445024 32700
rect 445076 32688 445082 32700
rect 545114 32688 545120 32700
rect 445076 32660 545120 32688
rect 445076 32648 445082 32660
rect 545114 32648 545120 32660
rect 545172 32648 545178 32700
rect 247034 32580 247040 32632
rect 247092 32620 247098 32632
rect 363046 32620 363052 32632
rect 247092 32592 363052 32620
rect 247092 32580 247098 32592
rect 363046 32580 363052 32592
rect 363104 32580 363110 32632
rect 425790 32580 425796 32632
rect 425848 32620 425854 32632
rect 531314 32620 531320 32632
rect 425848 32592 531320 32620
rect 425848 32580 425854 32592
rect 531314 32580 531320 32592
rect 531372 32580 531378 32632
rect 292482 32512 292488 32564
rect 292540 32552 292546 32564
rect 458174 32552 458180 32564
rect 292540 32524 458180 32552
rect 292540 32512 292546 32524
rect 458174 32512 458180 32524
rect 458232 32512 458238 32564
rect 81434 32444 81440 32496
rect 81492 32484 81498 32496
rect 181622 32484 181628 32496
rect 81492 32456 181628 32484
rect 81492 32444 81498 32456
rect 181622 32444 181628 32456
rect 181680 32444 181686 32496
rect 310422 32444 310428 32496
rect 310480 32484 310486 32496
rect 523034 32484 523040 32496
rect 310480 32456 523040 32484
rect 310480 32444 310486 32456
rect 523034 32444 523040 32456
rect 523092 32444 523098 32496
rect 40034 32376 40040 32428
rect 40092 32416 40098 32428
rect 108482 32416 108488 32428
rect 40092 32388 108488 32416
rect 40092 32376 40098 32388
rect 108482 32376 108488 32388
rect 108540 32376 108546 32428
rect 135254 32376 135260 32428
rect 135312 32416 135318 32428
rect 456978 32416 456984 32428
rect 135312 32388 456984 32416
rect 135312 32376 135318 32388
rect 456978 32376 456984 32388
rect 457036 32376 457042 32428
rect 253934 31356 253940 31408
rect 253992 31396 253998 31408
rect 364610 31396 364616 31408
rect 253992 31368 364616 31396
rect 253992 31356 253998 31368
rect 364610 31356 364616 31368
rect 364668 31356 364674 31408
rect 275922 31288 275928 31340
rect 275980 31328 275986 31340
rect 398834 31328 398840 31340
rect 275980 31300 398840 31328
rect 275980 31288 275986 31300
rect 398834 31288 398840 31300
rect 398892 31288 398898 31340
rect 340138 31220 340144 31272
rect 340196 31260 340202 31272
rect 506750 31260 506756 31272
rect 340196 31232 506756 31260
rect 340196 31220 340202 31232
rect 506750 31220 506756 31232
rect 506808 31220 506814 31272
rect 172514 31152 172520 31204
rect 172572 31192 172578 31204
rect 342254 31192 342260 31204
rect 172572 31164 342260 31192
rect 172572 31152 172578 31164
rect 342254 31152 342260 31164
rect 342312 31152 342318 31204
rect 441062 31152 441068 31204
rect 441120 31192 441126 31204
rect 531314 31192 531320 31204
rect 441120 31164 531320 31192
rect 441120 31152 441126 31164
rect 531314 31152 531320 31164
rect 531372 31152 531378 31204
rect 91094 31084 91100 31136
rect 91152 31124 91158 31136
rect 153838 31124 153844 31136
rect 91152 31096 153844 31124
rect 91152 31084 91158 31096
rect 153838 31084 153844 31096
rect 153896 31084 153902 31136
rect 307478 31084 307484 31136
rect 307536 31124 307542 31136
rect 514754 31124 514760 31136
rect 307536 31096 514760 31124
rect 307536 31084 307542 31096
rect 514754 31084 514760 31096
rect 514812 31084 514818 31136
rect 44174 31016 44180 31068
rect 44232 31056 44238 31068
rect 108298 31056 108304 31068
rect 44232 31028 108304 31056
rect 44232 31016 44238 31028
rect 108298 31016 108304 31028
rect 108356 31016 108362 31068
rect 187694 31016 187700 31068
rect 187752 31056 187758 31068
rect 470870 31056 470876 31068
rect 187752 31028 470876 31056
rect 187752 31016 187758 31028
rect 470870 31016 470876 31028
rect 470928 31016 470934 31068
rect 258074 29928 258080 29980
rect 258132 29968 258138 29980
rect 365714 29968 365720 29980
rect 258132 29940 365720 29968
rect 258132 29928 258138 29940
rect 365714 29928 365720 29940
rect 365772 29928 365778 29980
rect 274358 29860 274364 29912
rect 274416 29900 274422 29912
rect 394694 29900 394700 29912
rect 274416 29872 394700 29900
rect 274416 29860 274422 29872
rect 394694 29860 394700 29872
rect 394752 29860 394758 29912
rect 338758 29792 338764 29844
rect 338816 29832 338822 29844
rect 505094 29832 505100 29844
rect 338816 29804 505100 29832
rect 338816 29792 338822 29804
rect 505094 29792 505100 29804
rect 505152 29792 505158 29844
rect 176746 29724 176752 29776
rect 176804 29764 176810 29776
rect 343634 29764 343640 29776
rect 176804 29736 343640 29764
rect 176804 29724 176810 29736
rect 343634 29724 343640 29736
rect 343692 29724 343698 29776
rect 440878 29724 440884 29776
rect 440936 29764 440942 29776
rect 527174 29764 527180 29776
rect 440936 29736 527180 29764
rect 440936 29724 440942 29736
rect 527174 29724 527180 29736
rect 527232 29724 527238 29776
rect 49694 29656 49700 29708
rect 49752 29696 49758 29708
rect 173158 29696 173164 29708
rect 49752 29668 173164 29696
rect 49752 29656 49758 29668
rect 173158 29656 173164 29668
rect 173216 29656 173222 29708
rect 307662 29656 307668 29708
rect 307720 29696 307726 29708
rect 511994 29696 512000 29708
rect 307720 29668 512000 29696
rect 307720 29656 307726 29668
rect 511994 29656 512000 29668
rect 512052 29656 512058 29708
rect 4798 29588 4804 29640
rect 4856 29628 4862 29640
rect 131942 29628 131948 29640
rect 4856 29600 131948 29628
rect 4856 29588 4862 29600
rect 131942 29588 131948 29600
rect 132000 29588 132006 29640
rect 166994 29588 167000 29640
rect 167052 29628 167058 29640
rect 465166 29628 465172 29640
rect 167052 29600 465172 29628
rect 167052 29588 167058 29600
rect 465166 29588 465172 29600
rect 465224 29588 465230 29640
rect 274542 28500 274548 28552
rect 274600 28540 274606 28552
rect 390554 28540 390560 28552
rect 274600 28512 390560 28540
rect 274600 28500 274606 28512
rect 390554 28500 390560 28512
rect 390612 28500 390618 28552
rect 242894 28432 242900 28484
rect 242952 28472 242958 28484
rect 361574 28472 361580 28484
rect 242952 28444 361580 28472
rect 242952 28432 242958 28444
rect 361574 28432 361580 28444
rect 361632 28432 361638 28484
rect 364978 28432 364984 28484
rect 365036 28472 365042 28484
rect 516134 28472 516140 28484
rect 365036 28444 516140 28472
rect 365036 28432 365042 28444
rect 516134 28432 516140 28444
rect 516192 28432 516198 28484
rect 296622 28364 296628 28416
rect 296680 28404 296686 28416
rect 473354 28404 473360 28416
rect 296680 28376 473360 28404
rect 296680 28364 296686 28376
rect 473354 28364 473360 28376
rect 473412 28364 473418 28416
rect 10318 28296 10324 28348
rect 10376 28336 10382 28348
rect 131758 28336 131764 28348
rect 10376 28308 131764 28336
rect 10376 28296 10382 28308
rect 131758 28296 131764 28308
rect 131816 28296 131822 28348
rect 306282 28296 306288 28348
rect 306340 28336 306346 28348
rect 507854 28336 507860 28348
rect 306340 28308 507860 28336
rect 306340 28296 306346 28308
rect 507854 28296 507860 28308
rect 507912 28296 507918 28348
rect 131114 28228 131120 28280
rect 131172 28268 131178 28280
rect 455506 28268 455512 28280
rect 131172 28240 455512 28268
rect 131172 28228 131178 28240
rect 455506 28228 455512 28240
rect 455564 28228 455570 28280
rect 260834 27140 260840 27192
rect 260892 27180 260898 27192
rect 367278 27180 367284 27192
rect 260892 27152 367284 27180
rect 260892 27140 260898 27152
rect 367278 27140 367284 27152
rect 367336 27140 367342 27192
rect 270402 27072 270408 27124
rect 270460 27112 270466 27124
rect 380894 27112 380900 27124
rect 270460 27084 380900 27112
rect 270460 27072 270466 27084
rect 380894 27072 380900 27084
rect 380952 27072 380958 27124
rect 442258 27072 442264 27124
rect 442316 27112 442322 27124
rect 534074 27112 534080 27124
rect 442316 27084 534080 27112
rect 442316 27072 442322 27084
rect 534074 27072 534080 27084
rect 534132 27072 534138 27124
rect 293586 27004 293592 27056
rect 293644 27044 293650 27056
rect 462314 27044 462320 27056
rect 293644 27016 462320 27044
rect 293644 27004 293650 27016
rect 462314 27004 462320 27016
rect 462372 27004 462378 27056
rect 48314 26936 48320 26988
rect 48372 26976 48378 26988
rect 141602 26976 141608 26988
rect 48372 26948 141608 26976
rect 48372 26936 48378 26948
rect 141602 26936 141608 26948
rect 141660 26936 141666 26988
rect 304902 26936 304908 26988
rect 304960 26976 304966 26988
rect 505094 26976 505100 26988
rect 304960 26948 505100 26976
rect 304960 26936 304966 26948
rect 505094 26936 505100 26948
rect 505152 26936 505158 26988
rect 74534 26868 74540 26920
rect 74592 26908 74598 26920
rect 180058 26908 180064 26920
rect 74592 26880 180064 26908
rect 74592 26868 74598 26880
rect 180058 26868 180064 26880
rect 180116 26868 180122 26920
rect 266354 26868 266360 26920
rect 266412 26908 266418 26920
rect 492858 26908 492864 26920
rect 266412 26880 492864 26908
rect 266412 26868 266418 26880
rect 492858 26868 492864 26880
rect 492916 26868 492922 26920
rect 269022 25780 269028 25832
rect 269080 25820 269086 25832
rect 373994 25820 374000 25832
rect 269080 25792 374000 25820
rect 269080 25780 269086 25792
rect 373994 25780 374000 25792
rect 374052 25780 374058 25832
rect 286686 25712 286692 25764
rect 286744 25752 286750 25764
rect 437474 25752 437480 25764
rect 286744 25724 437480 25752
rect 286744 25712 286750 25724
rect 437474 25712 437480 25724
rect 437532 25712 437538 25764
rect 438118 25712 438124 25764
rect 438176 25752 438182 25764
rect 516134 25752 516140 25764
rect 438176 25724 516140 25752
rect 438176 25712 438182 25724
rect 516134 25712 516140 25724
rect 516192 25712 516198 25764
rect 140774 25644 140780 25696
rect 140832 25684 140838 25696
rect 329190 25684 329196 25696
rect 140832 25656 329196 25684
rect 140832 25644 140838 25656
rect 329190 25644 329196 25656
rect 329248 25644 329254 25696
rect 410610 25644 410616 25696
rect 410668 25684 410674 25696
rect 524506 25684 524512 25696
rect 410668 25656 524512 25684
rect 410668 25644 410674 25656
rect 524506 25644 524512 25656
rect 524564 25644 524570 25696
rect 153194 25576 153200 25628
rect 153252 25616 153258 25628
rect 207658 25616 207664 25628
rect 153252 25588 207664 25616
rect 153252 25576 153258 25588
rect 207658 25576 207664 25588
rect 207716 25576 207722 25628
rect 303338 25576 303344 25628
rect 303396 25616 303402 25628
rect 500954 25616 500960 25628
rect 303396 25588 500960 25616
rect 303396 25576 303402 25588
rect 500954 25576 500960 25588
rect 501012 25576 501018 25628
rect 35894 25508 35900 25560
rect 35952 25548 35958 25560
rect 106918 25548 106924 25560
rect 35952 25520 106924 25548
rect 35952 25508 35958 25520
rect 106918 25508 106924 25520
rect 106976 25508 106982 25560
rect 201586 25508 201592 25560
rect 201644 25548 201650 25560
rect 474734 25548 474740 25560
rect 201644 25520 474740 25548
rect 201644 25508 201650 25520
rect 474734 25508 474740 25520
rect 474792 25508 474798 25560
rect 267366 24420 267372 24472
rect 267424 24460 267430 24472
rect 365714 24460 365720 24472
rect 267424 24432 365720 24460
rect 267424 24420 267430 24432
rect 365714 24420 365720 24432
rect 365772 24420 365778 24472
rect 264974 24352 264980 24404
rect 265032 24392 265038 24404
rect 367094 24392 367100 24404
rect 265032 24364 367100 24392
rect 265032 24352 265038 24364
rect 367094 24352 367100 24364
rect 367152 24352 367158 24404
rect 285582 24284 285588 24336
rect 285640 24324 285646 24336
rect 433334 24324 433340 24336
rect 285640 24296 433340 24324
rect 285640 24284 285646 24296
rect 433334 24284 433340 24296
rect 433392 24284 433398 24336
rect 433978 24284 433984 24336
rect 434036 24324 434042 24336
rect 506474 24324 506480 24336
rect 434036 24296 506480 24324
rect 434036 24284 434042 24296
rect 506474 24284 506480 24296
rect 506532 24284 506538 24336
rect 303522 24216 303528 24268
rect 303580 24256 303586 24268
rect 498194 24256 498200 24268
rect 303580 24228 498200 24256
rect 303580 24216 303586 24228
rect 498194 24216 498200 24228
rect 498252 24216 498258 24268
rect 135346 24148 135352 24200
rect 135404 24188 135410 24200
rect 203518 24188 203524 24200
rect 135404 24160 203524 24188
rect 135404 24148 135410 24160
rect 203518 24148 203524 24160
rect 203576 24148 203582 24200
rect 266998 24148 267004 24200
rect 267056 24188 267062 24200
rect 490006 24188 490012 24200
rect 267056 24160 490012 24188
rect 267056 24148 267062 24160
rect 490006 24148 490012 24160
rect 490064 24148 490070 24200
rect 26234 24080 26240 24132
rect 26292 24120 26298 24132
rect 104158 24120 104164 24132
rect 26292 24092 104164 24120
rect 26292 24080 26298 24092
rect 104158 24080 104164 24092
rect 104216 24080 104222 24132
rect 149054 24080 149060 24132
rect 149112 24120 149118 24132
rect 461026 24120 461032 24132
rect 149112 24092 461032 24120
rect 149112 24080 149118 24092
rect 461026 24080 461032 24092
rect 461084 24080 461090 24132
rect 271782 22992 271788 23044
rect 271840 23032 271846 23044
rect 383654 23032 383660 23044
rect 271840 23004 383660 23032
rect 271840 22992 271846 23004
rect 383654 22992 383660 23004
rect 383712 22992 383718 23044
rect 439498 22992 439504 23044
rect 439556 23032 439562 23044
rect 523126 23032 523132 23044
rect 439556 23004 523132 23032
rect 439556 22992 439562 23004
rect 523126 22992 523132 23004
rect 523184 22992 523190 23044
rect 288342 22924 288348 22976
rect 288400 22964 288406 22976
rect 444374 22964 444380 22976
rect 288400 22936 444380 22964
rect 288400 22924 288406 22936
rect 444374 22924 444380 22936
rect 444432 22924 444438 22976
rect 132494 22856 132500 22908
rect 132552 22896 132558 22908
rect 202138 22896 202144 22908
rect 132552 22868 202144 22896
rect 132552 22856 132558 22868
rect 202138 22856 202144 22868
rect 202196 22856 202202 22908
rect 242802 22856 242808 22908
rect 242860 22896 242866 22908
rect 277394 22896 277400 22908
rect 242860 22868 277400 22896
rect 242860 22856 242866 22868
rect 277394 22856 277400 22868
rect 277452 22856 277458 22908
rect 300670 22856 300676 22908
rect 300728 22896 300734 22908
rect 489914 22896 489920 22908
rect 300728 22868 489920 22896
rect 300728 22856 300734 22868
rect 489914 22856 489920 22868
rect 489972 22856 489978 22908
rect 158714 22788 158720 22840
rect 158772 22828 158778 22840
rect 333238 22828 333244 22840
rect 158772 22800 333244 22828
rect 158772 22788 158778 22800
rect 333238 22788 333244 22800
rect 333296 22788 333302 22840
rect 411254 22788 411260 22840
rect 411312 22828 411318 22840
rect 532878 22828 532884 22840
rect 411312 22800 532884 22828
rect 411312 22788 411318 22800
rect 532878 22788 532884 22800
rect 532936 22788 532942 22840
rect 52454 22720 52460 22772
rect 52512 22760 52518 22772
rect 142798 22760 142804 22772
rect 52512 22732 142804 22760
rect 52512 22720 52518 22732
rect 142798 22720 142804 22732
rect 142856 22720 142862 22772
rect 262858 22720 262864 22772
rect 262916 22760 262922 22772
rect 490190 22760 490196 22772
rect 262916 22732 490196 22760
rect 262916 22720 262922 22732
rect 490190 22720 490196 22732
rect 490248 22720 490254 22772
rect 235994 21632 236000 21684
rect 236052 21672 236058 21684
rect 360194 21672 360200 21684
rect 236052 21644 360200 21672
rect 236052 21632 236058 21644
rect 360194 21632 360200 21644
rect 360252 21632 360258 21684
rect 179414 21564 179420 21616
rect 179472 21604 179478 21616
rect 345198 21604 345204 21616
rect 179472 21576 345204 21604
rect 179472 21564 179478 21576
rect 345198 21564 345204 21576
rect 345256 21564 345262 21616
rect 356698 21564 356704 21616
rect 356756 21604 356762 21616
rect 514846 21604 514852 21616
rect 356756 21576 514852 21604
rect 356756 21564 356762 21576
rect 514846 21564 514852 21576
rect 514904 21564 514910 21616
rect 300486 21496 300492 21548
rect 300544 21536 300550 21548
rect 487154 21536 487160 21548
rect 300544 21508 487160 21536
rect 300544 21496 300550 21508
rect 487154 21496 487160 21508
rect 487212 21496 487218 21548
rect 242158 21428 242164 21480
rect 242216 21468 242222 21480
rect 484394 21468 484400 21480
rect 242216 21440 484400 21468
rect 242216 21428 242222 21440
rect 484394 21428 484400 21440
rect 484452 21428 484458 21480
rect 33134 21360 33140 21412
rect 33192 21400 33198 21412
rect 105538 21400 105544 21412
rect 33192 21372 105544 21400
rect 33192 21360 33198 21372
rect 105538 21360 105544 21372
rect 105596 21360 105602 21412
rect 128354 21360 128360 21412
rect 128412 21400 128418 21412
rect 200942 21400 200948 21412
rect 128412 21372 200948 21400
rect 128412 21360 128418 21372
rect 200942 21360 200948 21372
rect 201000 21360 201006 21412
rect 241238 21360 241244 21412
rect 241296 21400 241302 21412
rect 270494 21400 270500 21412
rect 241296 21372 270500 21400
rect 241296 21360 241302 21372
rect 270494 21360 270500 21372
rect 270552 21360 270558 21412
rect 324130 21360 324136 21412
rect 324188 21400 324194 21412
rect 574738 21400 574744 21412
rect 324188 21372 574744 21400
rect 324188 21360 324194 21372
rect 574738 21360 574744 21372
rect 574796 21360 574802 21412
rect 271874 20272 271880 20324
rect 271932 20312 271938 20324
rect 369946 20312 369952 20324
rect 271932 20284 369952 20312
rect 271932 20272 271938 20284
rect 369946 20272 369952 20284
rect 370004 20272 370010 20324
rect 218054 20204 218060 20256
rect 218112 20244 218118 20256
rect 354674 20244 354680 20256
rect 218112 20216 354680 20244
rect 218112 20204 218118 20216
rect 354674 20204 354680 20216
rect 354732 20204 354738 20256
rect 299382 20136 299388 20188
rect 299440 20176 299446 20188
rect 483014 20176 483020 20188
rect 299440 20148 483020 20176
rect 299440 20136 299446 20148
rect 483014 20136 483020 20148
rect 483072 20136 483078 20188
rect 302878 20068 302884 20120
rect 302936 20108 302942 20120
rect 491294 20108 491300 20120
rect 302936 20080 491300 20108
rect 302936 20068 302942 20080
rect 491294 20068 491300 20080
rect 491352 20068 491358 20120
rect 103514 20000 103520 20052
rect 103572 20040 103578 20052
rect 125042 20040 125048 20052
rect 103572 20012 125048 20040
rect 103572 20000 103578 20012
rect 125042 20000 125048 20012
rect 125100 20000 125106 20052
rect 126974 20000 126980 20052
rect 127032 20040 127038 20052
rect 324958 20040 324964 20052
rect 127032 20012 324964 20040
rect 127032 20000 127038 20012
rect 324958 20000 324964 20012
rect 325016 20000 325022 20052
rect 404998 20000 405004 20052
rect 405056 20040 405062 20052
rect 526070 20040 526076 20052
rect 405056 20012 526076 20040
rect 405056 20000 405062 20012
rect 526070 20000 526076 20012
rect 526128 20000 526134 20052
rect 14458 19932 14464 19984
rect 14516 19972 14522 19984
rect 133138 19972 133144 19984
rect 14516 19944 133144 19972
rect 14516 19932 14522 19944
rect 133138 19932 133144 19944
rect 133196 19932 133202 19984
rect 185026 19932 185032 19984
rect 185084 19972 185090 19984
rect 217502 19972 217508 19984
rect 185084 19944 217508 19972
rect 185084 19932 185090 19944
rect 217502 19932 217508 19944
rect 217560 19932 217566 19984
rect 238478 19932 238484 19984
rect 238536 19972 238542 19984
rect 263594 19972 263600 19984
rect 238536 19944 263600 19972
rect 238536 19932 238542 19944
rect 263594 19932 263600 19944
rect 263652 19932 263658 19984
rect 323946 19932 323952 19984
rect 324004 19972 324010 19984
rect 572714 19972 572720 19984
rect 324004 19944 572720 19972
rect 324004 19932 324010 19944
rect 572714 19932 572720 19944
rect 572772 19932 572778 19984
rect 233234 18844 233240 18896
rect 233292 18884 233298 18896
rect 358906 18884 358912 18896
rect 233292 18856 358912 18884
rect 233292 18844 233298 18856
rect 358906 18844 358912 18856
rect 358964 18844 358970 18896
rect 183554 18776 183560 18828
rect 183612 18816 183618 18828
rect 345014 18816 345020 18828
rect 183612 18788 345020 18816
rect 183612 18776 183618 18788
rect 345014 18776 345020 18788
rect 345072 18776 345078 18828
rect 345658 18776 345664 18828
rect 345716 18816 345722 18828
rect 512086 18816 512092 18828
rect 345716 18788 512092 18816
rect 345716 18776 345722 18788
rect 512086 18776 512092 18788
rect 512144 18776 512150 18828
rect 297726 18708 297732 18760
rect 297784 18748 297790 18760
rect 480254 18748 480260 18760
rect 297784 18720 480260 18748
rect 297784 18708 297790 18720
rect 480254 18708 480260 18720
rect 480312 18708 480318 18760
rect 100754 18640 100760 18692
rect 100812 18680 100818 18692
rect 124858 18680 124864 18692
rect 100812 18652 124864 18680
rect 100812 18640 100818 18652
rect 124858 18640 124864 18652
rect 124916 18640 124922 18692
rect 238662 18640 238668 18692
rect 238720 18680 238726 18692
rect 259454 18680 259460 18692
rect 238720 18652 259460 18680
rect 238720 18640 238726 18652
rect 259454 18640 259460 18652
rect 259512 18640 259518 18692
rect 322842 18640 322848 18692
rect 322900 18680 322906 18692
rect 568574 18680 568580 18692
rect 322900 18652 568580 18680
rect 322900 18640 322906 18652
rect 568574 18640 568580 18652
rect 568632 18640 568638 18692
rect 4890 18572 4896 18624
rect 4948 18612 4954 18624
rect 98638 18612 98644 18624
rect 4948 18584 98644 18612
rect 4948 18572 4954 18584
rect 98638 18572 98644 18584
rect 98696 18572 98702 18624
rect 109034 18572 109040 18624
rect 109092 18612 109098 18624
rect 158162 18612 158168 18624
rect 109092 18584 158168 18612
rect 109092 18572 109098 18584
rect 158162 18572 158168 18584
rect 158220 18572 158226 18624
rect 178034 18572 178040 18624
rect 178092 18612 178098 18624
rect 214558 18612 214564 18624
rect 178092 18584 214564 18612
rect 178092 18572 178098 18584
rect 214558 18572 214564 18584
rect 214616 18572 214622 18624
rect 223574 18572 223580 18624
rect 223632 18612 223638 18624
rect 480530 18612 480536 18624
rect 223632 18584 480536 18612
rect 223632 18572 223638 18584
rect 480530 18572 480536 18584
rect 480588 18572 480594 18624
rect 322934 17688 322940 17740
rect 322992 17728 322998 17740
rect 507946 17728 507952 17740
rect 322992 17700 507952 17728
rect 322992 17688 322998 17700
rect 507946 17688 507952 17700
rect 508004 17688 508010 17740
rect 316126 17620 316132 17672
rect 316184 17660 316190 17672
rect 506566 17660 506572 17672
rect 316184 17632 506572 17660
rect 316184 17620 316190 17632
rect 506566 17620 506572 17632
rect 506624 17620 506630 17672
rect 304994 17552 305000 17604
rect 305052 17592 305058 17604
rect 503714 17592 503720 17604
rect 305052 17564 503720 17592
rect 305052 17552 305058 17564
rect 503714 17552 503720 17564
rect 503772 17552 503778 17604
rect 160094 17484 160100 17536
rect 160152 17524 160158 17536
rect 463786 17524 463792 17536
rect 160152 17496 463792 17524
rect 160152 17484 160158 17496
rect 463786 17484 463792 17496
rect 463844 17484 463850 17536
rect 155954 17416 155960 17468
rect 156012 17456 156018 17468
rect 462406 17456 462412 17468
rect 156012 17428 462412 17456
rect 156012 17416 156018 17428
rect 462406 17416 462412 17428
rect 462464 17416 462470 17468
rect 151814 17348 151820 17400
rect 151872 17388 151878 17400
rect 461210 17388 461216 17400
rect 151872 17360 461216 17388
rect 151872 17348 151878 17360
rect 461210 17348 461216 17360
rect 461268 17348 461274 17400
rect 55214 17280 55220 17332
rect 55272 17320 55278 17332
rect 144362 17320 144368 17332
rect 55272 17292 144368 17320
rect 55272 17280 55278 17292
rect 144362 17280 144368 17292
rect 144420 17280 144426 17332
rect 144914 17280 144920 17332
rect 144972 17320 144978 17332
rect 459554 17320 459560 17332
rect 144972 17292 459560 17320
rect 144972 17280 144978 17292
rect 459554 17280 459560 17292
rect 459612 17280 459618 17332
rect 96614 17212 96620 17264
rect 96672 17252 96678 17264
rect 123478 17252 123484 17264
rect 96672 17224 123484 17252
rect 96672 17212 96678 17224
rect 123478 17212 123484 17224
rect 123536 17212 123542 17264
rect 142154 17212 142160 17264
rect 142212 17252 142218 17264
rect 458266 17252 458272 17264
rect 142212 17224 458272 17252
rect 142212 17212 142218 17224
rect 458266 17212 458272 17224
rect 458324 17212 458330 17264
rect 298094 16396 298100 16448
rect 298152 16436 298158 16448
rect 501046 16436 501052 16448
rect 298152 16408 501052 16436
rect 298152 16396 298158 16408
rect 501046 16396 501052 16408
rect 501104 16396 501110 16448
rect 294874 16328 294880 16380
rect 294932 16368 294938 16380
rect 499666 16368 499672 16380
rect 294932 16340 499672 16368
rect 294932 16328 294938 16340
rect 499666 16328 499672 16340
rect 499724 16328 499730 16380
rect 291378 16260 291384 16312
rect 291436 16300 291442 16312
rect 499850 16300 499856 16312
rect 291436 16272 499856 16300
rect 291436 16260 291442 16272
rect 499850 16260 499856 16272
rect 499908 16260 499914 16312
rect 287330 16192 287336 16244
rect 287388 16232 287394 16244
rect 498286 16232 498292 16244
rect 287388 16204 498292 16232
rect 287388 16192 287394 16204
rect 498286 16192 498292 16204
rect 498344 16192 498350 16244
rect 284386 16124 284392 16176
rect 284444 16164 284450 16176
rect 497090 16164 497096 16176
rect 284444 16136 497096 16164
rect 284444 16124 284450 16136
rect 497090 16124 497096 16136
rect 497148 16124 497154 16176
rect 280706 16056 280712 16108
rect 280764 16096 280770 16108
rect 496906 16096 496912 16108
rect 280764 16068 496912 16096
rect 280764 16056 280770 16068
rect 496906 16056 496912 16068
rect 496964 16056 496970 16108
rect 83274 15988 83280 16040
rect 83332 16028 83338 16040
rect 119338 16028 119344 16040
rect 83332 16000 119344 16028
rect 83332 15988 83338 16000
rect 119338 15988 119344 16000
rect 119396 15988 119402 16040
rect 276658 15988 276664 16040
rect 276716 16028 276722 16040
rect 495434 16028 495440 16040
rect 276716 16000 495440 16028
rect 276716 15988 276722 16000
rect 495434 15988 495440 16000
rect 495492 15988 495498 16040
rect 102226 15920 102232 15972
rect 102284 15960 102290 15972
rect 156598 15960 156604 15972
rect 102284 15932 156604 15960
rect 102284 15920 102290 15932
rect 156598 15920 156604 15932
rect 156656 15920 156662 15972
rect 160646 15920 160652 15972
rect 160704 15960 160710 15972
rect 210602 15960 210608 15972
rect 160704 15932 210608 15960
rect 160704 15920 160710 15932
rect 210602 15920 210608 15932
rect 210660 15920 210666 15972
rect 273254 15920 273260 15972
rect 273312 15960 273318 15972
rect 494146 15960 494152 15972
rect 273312 15932 494152 15960
rect 273312 15920 273318 15932
rect 494146 15920 494152 15932
rect 494204 15920 494210 15972
rect 15838 15852 15844 15904
rect 15896 15892 15902 15904
rect 165062 15892 165068 15904
rect 15896 15864 165068 15892
rect 15896 15852 15902 15864
rect 165062 15852 165068 15864
rect 165120 15852 165126 15904
rect 209774 15852 209780 15904
rect 209832 15892 209838 15904
rect 224402 15892 224408 15904
rect 209832 15864 224408 15892
rect 209832 15852 209838 15864
rect 224402 15852 224408 15864
rect 224460 15852 224466 15904
rect 235902 15852 235908 15904
rect 235960 15892 235966 15904
rect 253106 15892 253112 15904
rect 235960 15864 253112 15892
rect 235960 15852 235966 15864
rect 253106 15852 253112 15864
rect 253164 15852 253170 15904
rect 270034 15852 270040 15904
rect 270092 15892 270098 15904
rect 492674 15892 492680 15904
rect 270092 15864 492680 15892
rect 270092 15852 270098 15864
rect 492674 15852 492680 15864
rect 492732 15852 492738 15904
rect 528554 15852 528560 15904
rect 528612 15892 528618 15904
rect 564526 15892 564532 15904
rect 528612 15864 564532 15892
rect 528612 15852 528618 15864
rect 564526 15852 564532 15864
rect 564584 15852 564590 15904
rect 234614 14832 234620 14884
rect 234672 14872 234678 14884
rect 483106 14872 483112 14884
rect 234672 14844 483112 14872
rect 234672 14832 234678 14844
rect 483106 14832 483112 14844
rect 483164 14832 483170 14884
rect 231026 14764 231032 14816
rect 231084 14804 231090 14816
rect 483290 14804 483296 14816
rect 231084 14776 483296 14804
rect 231084 14764 231090 14776
rect 483290 14764 483296 14776
rect 483348 14764 483354 14816
rect 226334 14696 226340 14748
rect 226392 14736 226398 14748
rect 481634 14736 481640 14748
rect 226392 14708 481640 14736
rect 226392 14696 226398 14708
rect 481634 14696 481640 14708
rect 481692 14696 481698 14748
rect 216858 14628 216864 14680
rect 216916 14668 216922 14680
rect 478874 14668 478880 14680
rect 216916 14640 478880 14668
rect 216916 14628 216922 14640
rect 478874 14628 478880 14640
rect 478932 14628 478938 14680
rect 164418 14560 164424 14612
rect 164476 14600 164482 14612
rect 210418 14600 210424 14612
rect 164476 14572 210424 14600
rect 164476 14560 164482 14572
rect 210418 14560 210424 14572
rect 210476 14560 210482 14612
rect 213362 14560 213368 14612
rect 213420 14600 213426 14612
rect 477494 14600 477500 14612
rect 213420 14572 477500 14600
rect 213420 14560 213426 14572
rect 477494 14560 477500 14572
rect 477552 14560 477558 14612
rect 72602 14492 72608 14544
rect 72660 14532 72666 14544
rect 116578 14532 116584 14544
rect 72660 14504 116584 14532
rect 72660 14492 72666 14504
rect 116578 14492 116584 14504
rect 116636 14492 116642 14544
rect 209866 14492 209872 14544
rect 209924 14532 209930 14544
rect 476298 14532 476304 14544
rect 209924 14504 476304 14532
rect 209924 14492 209930 14504
rect 476298 14492 476304 14504
rect 476356 14492 476362 14544
rect 84194 14424 84200 14476
rect 84252 14464 84258 14476
rect 151078 14464 151084 14476
rect 84252 14436 151084 14464
rect 84252 14424 84258 14436
rect 151078 14424 151084 14436
rect 151136 14424 151142 14476
rect 206186 14424 206192 14476
rect 206244 14464 206250 14476
rect 476482 14464 476488 14476
rect 206244 14436 476488 14464
rect 206244 14424 206250 14436
rect 476482 14424 476488 14436
rect 476540 14424 476546 14476
rect 507210 14424 507216 14476
rect 507268 14464 507274 14476
rect 559098 14464 559104 14476
rect 507268 14436 559104 14464
rect 507268 14424 507274 14436
rect 559098 14424 559104 14436
rect 559156 14424 559162 14476
rect 151906 13472 151912 13524
rect 151964 13512 151970 13524
rect 331858 13512 331864 13524
rect 151964 13484 331864 13512
rect 151964 13472 151970 13484
rect 331858 13472 331864 13484
rect 331916 13472 331922 13524
rect 147858 13404 147864 13456
rect 147916 13444 147922 13456
rect 330478 13444 330484 13456
rect 147916 13416 330484 13444
rect 147916 13404 147922 13416
rect 330478 13404 330484 13416
rect 330536 13404 330542 13456
rect 143534 13336 143540 13388
rect 143592 13376 143598 13388
rect 330662 13376 330668 13388
rect 143592 13348 330668 13376
rect 143592 13336 143598 13348
rect 330662 13336 330668 13348
rect 330720 13336 330726 13388
rect 449158 13336 449164 13388
rect 449216 13376 449222 13388
rect 559282 13376 559288 13388
rect 449216 13348 559288 13376
rect 449216 13336 449222 13348
rect 559282 13336 559288 13348
rect 559340 13336 559346 13388
rect 173894 13268 173900 13320
rect 173952 13308 173958 13320
rect 466546 13308 466552 13320
rect 173952 13280 466552 13308
rect 173952 13268 173958 13280
rect 466546 13268 466552 13280
rect 466604 13268 466610 13320
rect 170306 13200 170312 13252
rect 170364 13240 170370 13252
rect 466730 13240 466736 13252
rect 170364 13212 466736 13240
rect 170364 13200 170370 13212
rect 466730 13200 466736 13212
rect 466788 13200 466794 13252
rect 41874 13132 41880 13184
rect 41932 13172 41938 13184
rect 140038 13172 140044 13184
rect 41932 13144 140044 13172
rect 41932 13132 41938 13144
rect 140038 13132 140044 13144
rect 140096 13132 140102 13184
rect 163682 13132 163688 13184
rect 163740 13172 163746 13184
rect 463970 13172 463976 13184
rect 163740 13144 463976 13172
rect 163740 13132 163746 13144
rect 463970 13132 463976 13144
rect 464028 13132 464034 13184
rect 58434 13064 58440 13116
rect 58492 13104 58498 13116
rect 112438 13104 112444 13116
rect 58492 13076 112444 13104
rect 58492 13064 58498 13076
rect 112438 13064 112444 13076
rect 112496 13064 112502 13116
rect 127526 13064 127532 13116
rect 127584 13104 127590 13116
rect 454034 13104 454040 13116
rect 127584 13076 454040 13104
rect 127584 13064 127590 13076
rect 454034 13064 454040 13076
rect 454092 13064 454098 13116
rect 374086 12112 374092 12164
rect 374144 12152 374150 12164
rect 397454 12152 397460 12164
rect 374144 12124 397460 12152
rect 374144 12112 374150 12124
rect 397454 12112 397460 12124
rect 397512 12112 397518 12164
rect 286594 11976 286600 12028
rect 286652 12016 286658 12028
rect 374362 12016 374368 12028
rect 286652 11988 374368 12016
rect 286652 11976 286658 11988
rect 374362 11976 374368 11988
rect 374420 11976 374426 12028
rect 279050 11908 279056 11960
rect 279108 11948 279114 11960
rect 371418 11948 371424 11960
rect 279108 11920 371424 11948
rect 279108 11908 279114 11920
rect 371418 11908 371424 11920
rect 371476 11908 371482 11960
rect 435358 11908 435364 11960
rect 435416 11948 435422 11960
rect 509602 11948 509608 11960
rect 435416 11920 509608 11948
rect 435416 11908 435422 11920
rect 509602 11908 509608 11920
rect 509660 11908 509666 11960
rect 268378 11840 268384 11892
rect 268436 11880 268442 11892
rect 368474 11880 368480 11892
rect 268436 11852 368480 11880
rect 268436 11840 268442 11852
rect 368474 11840 368480 11852
rect 368532 11840 368538 11892
rect 370498 11840 370504 11892
rect 370556 11880 370562 11892
rect 517514 11880 517520 11892
rect 370556 11852 517520 11880
rect 370556 11840 370562 11852
rect 517514 11840 517520 11852
rect 517572 11840 517578 11892
rect 108114 11772 108120 11824
rect 108172 11812 108178 11824
rect 126238 11812 126244 11824
rect 108172 11784 126244 11812
rect 108172 11772 108178 11784
rect 126238 11772 126244 11784
rect 126296 11772 126302 11824
rect 137186 11772 137192 11824
rect 137244 11812 137250 11824
rect 327718 11812 327724 11824
rect 137244 11784 327724 11812
rect 137244 11772 137250 11784
rect 327718 11772 327724 11784
rect 327776 11772 327782 11824
rect 340966 11772 340972 11824
rect 341024 11812 341030 11824
rect 513650 11812 513656 11824
rect 341024 11784 513656 11812
rect 341024 11772 341030 11784
rect 513650 11772 513656 11784
rect 513708 11772 513714 11824
rect 51074 11704 51080 11756
rect 51132 11744 51138 11756
rect 111058 11744 111064 11756
rect 51132 11716 111064 11744
rect 51132 11704 51138 11716
rect 111058 11704 111064 11716
rect 111116 11704 111122 11756
rect 176654 11704 176660 11756
rect 176712 11744 176718 11756
rect 177850 11744 177856 11756
rect 176712 11716 177856 11744
rect 176712 11704 176718 11716
rect 177850 11704 177856 11716
rect 177908 11704 177914 11756
rect 255958 11704 255964 11756
rect 256016 11744 256022 11756
rect 488534 11744 488540 11756
rect 256016 11716 488540 11744
rect 256016 11704 256022 11716
rect 488534 11704 488540 11716
rect 488592 11704 488598 11756
rect 517882 11704 517888 11756
rect 517940 11744 517946 11756
rect 561766 11744 561772 11756
rect 517940 11716 561772 11744
rect 517940 11704 517946 11716
rect 561766 11704 561772 11716
rect 561824 11704 561830 11756
rect 582374 11704 582380 11756
rect 582432 11744 582438 11756
rect 583386 11744 583392 11756
rect 582432 11716 583392 11744
rect 582432 11704 582438 11716
rect 583386 11704 583392 11716
rect 583444 11704 583450 11756
rect 425514 10616 425520 10668
rect 425572 10656 425578 10668
rect 536926 10656 536932 10668
rect 425572 10628 536932 10656
rect 425572 10616 425578 10628
rect 536926 10616 536932 10628
rect 536984 10616 536990 10668
rect 318058 10548 318064 10600
rect 318116 10588 318122 10600
rect 382274 10588 382280 10600
rect 318116 10560 382280 10588
rect 318116 10548 318122 10560
rect 382274 10548 382280 10560
rect 382332 10548 382338 10600
rect 418522 10548 418528 10600
rect 418580 10588 418586 10600
rect 534166 10588 534172 10600
rect 418580 10560 534172 10588
rect 418580 10548 418586 10560
rect 534166 10548 534172 10560
rect 534224 10548 534230 10600
rect 229370 10480 229376 10532
rect 229428 10520 229434 10532
rect 357526 10520 357532 10532
rect 229428 10492 357532 10520
rect 229428 10480 229434 10492
rect 357526 10480 357532 10492
rect 357584 10480 357590 10532
rect 400214 10480 400220 10532
rect 400272 10520 400278 10532
rect 530026 10520 530032 10532
rect 400272 10492 530032 10520
rect 400272 10480 400278 10492
rect 530026 10480 530032 10492
rect 530084 10480 530090 10532
rect 171686 10412 171692 10464
rect 171744 10452 171750 10464
rect 213178 10452 213184 10464
rect 171744 10424 213184 10452
rect 171744 10412 171750 10424
rect 213178 10412 213184 10424
rect 213236 10412 213242 10464
rect 222746 10412 222752 10464
rect 222804 10452 222810 10464
rect 356054 10452 356060 10464
rect 222804 10424 356060 10452
rect 222804 10412 222810 10424
rect 356054 10412 356060 10424
rect 356112 10412 356118 10464
rect 393314 10412 393320 10464
rect 393372 10452 393378 10464
rect 527266 10452 527272 10464
rect 393372 10424 527272 10452
rect 393372 10412 393378 10424
rect 527266 10412 527272 10424
rect 527324 10412 527330 10464
rect 69106 10344 69112 10396
rect 69164 10384 69170 10396
rect 115198 10384 115204 10396
rect 69164 10356 115204 10384
rect 69164 10344 69170 10356
rect 115198 10344 115204 10356
rect 115256 10344 115262 10396
rect 125594 10344 125600 10396
rect 125652 10384 125658 10396
rect 200758 10384 200764 10396
rect 125652 10356 200764 10384
rect 125652 10344 125658 10356
rect 200758 10344 200764 10356
rect 200816 10344 200822 10396
rect 211706 10344 211712 10396
rect 211764 10384 211770 10396
rect 353294 10384 353300 10396
rect 211764 10356 353300 10384
rect 211764 10344 211770 10356
rect 353294 10344 353300 10356
rect 353352 10344 353358 10396
rect 386414 10344 386420 10396
rect 386472 10384 386478 10396
rect 525886 10384 525892 10396
rect 386472 10356 525892 10384
rect 386472 10344 386478 10356
rect 525886 10344 525892 10356
rect 525944 10344 525950 10396
rect 30834 10276 30840 10328
rect 30892 10316 30898 10328
rect 137278 10316 137284 10328
rect 30892 10288 137284 10316
rect 30892 10276 30898 10288
rect 137278 10276 137284 10288
rect 137336 10276 137342 10328
rect 208578 10276 208584 10328
rect 208636 10316 208642 10328
rect 352190 10316 352196 10328
rect 208636 10288 352196 10316
rect 208636 10276 208642 10288
rect 352190 10276 352196 10288
rect 352248 10276 352254 10328
rect 369394 10276 369400 10328
rect 369452 10316 369458 10328
rect 520366 10316 520372 10328
rect 369452 10288 520372 10316
rect 369452 10276 369458 10288
rect 520366 10276 520372 10288
rect 520424 10276 520430 10328
rect 151722 9596 151728 9648
rect 151780 9636 151786 9648
rect 153010 9636 153016 9648
rect 151780 9608 153016 9636
rect 151780 9596 151786 9608
rect 153010 9596 153016 9608
rect 153068 9596 153074 9648
rect 209682 9596 209688 9648
rect 209740 9636 209746 9648
rect 210970 9636 210976 9648
rect 209740 9608 210976 9636
rect 209740 9596 209746 9608
rect 210970 9596 210976 9608
rect 211028 9596 211034 9648
rect 421742 9324 421748 9376
rect 421800 9364 421806 9376
rect 460382 9364 460388 9376
rect 421800 9336 460388 9364
rect 421800 9324 421806 9336
rect 460382 9324 460388 9336
rect 460440 9324 460446 9376
rect 422938 9256 422944 9308
rect 422996 9296 423002 9308
rect 463970 9296 463976 9308
rect 422996 9268 463976 9296
rect 422996 9256 423002 9268
rect 463970 9256 463976 9268
rect 464028 9256 464034 9308
rect 96246 9188 96252 9240
rect 96304 9228 96310 9240
rect 185578 9228 185584 9240
rect 96304 9200 185584 9228
rect 96304 9188 96310 9200
rect 185578 9188 185584 9200
rect 185636 9188 185642 9240
rect 297266 9188 297272 9240
rect 297324 9228 297330 9240
rect 376846 9228 376852 9240
rect 297324 9200 376852 9228
rect 297324 9188 297330 9200
rect 376846 9188 376852 9200
rect 376904 9188 376910 9240
rect 424502 9188 424508 9240
rect 424560 9228 424566 9240
rect 467466 9228 467472 9240
rect 424560 9200 467472 9228
rect 424560 9188 424566 9200
rect 467466 9188 467472 9200
rect 467524 9188 467530 9240
rect 24210 9120 24216 9172
rect 24268 9160 24274 9172
rect 166258 9160 166264 9172
rect 24268 9132 166264 9160
rect 24268 9120 24274 9132
rect 166258 9120 166264 9132
rect 166316 9120 166322 9172
rect 169570 9120 169576 9172
rect 169628 9160 169634 9172
rect 335998 9160 336004 9172
rect 169628 9132 336004 9160
rect 169628 9120 169634 9132
rect 335998 9120 336004 9132
rect 336056 9120 336062 9172
rect 424318 9120 424324 9172
rect 424376 9160 424382 9172
rect 471054 9160 471060 9172
rect 424376 9132 471060 9160
rect 424376 9120 424382 9132
rect 471054 9120 471060 9132
rect 471112 9120 471118 9172
rect 166074 9052 166080 9104
rect 166132 9092 166138 9104
rect 336182 9092 336188 9104
rect 166132 9064 336188 9092
rect 166132 9052 166138 9064
rect 336182 9052 336188 9064
rect 336240 9052 336246 9104
rect 427078 9052 427084 9104
rect 427136 9092 427142 9104
rect 478138 9092 478144 9104
rect 427136 9064 478144 9092
rect 427136 9052 427142 9064
rect 478138 9052 478144 9064
rect 478196 9052 478202 9104
rect 162486 8984 162492 9036
rect 162544 9024 162550 9036
rect 334618 9024 334624 9036
rect 162544 8996 334624 9024
rect 162544 8984 162550 8996
rect 334618 8984 334624 8996
rect 334676 8984 334682 9036
rect 450906 8984 450912 9036
rect 450964 9024 450970 9036
rect 542538 9024 542544 9036
rect 450964 8996 542544 9024
rect 450964 8984 450970 8996
rect 542538 8984 542544 8996
rect 542596 8984 542602 9036
rect 19426 8916 19432 8968
rect 19484 8956 19490 8968
rect 164878 8956 164884 8968
rect 19484 8928 164884 8956
rect 19484 8916 19490 8928
rect 164878 8916 164884 8928
rect 164936 8916 164942 8968
rect 295242 8916 295248 8968
rect 295300 8956 295306 8968
rect 469858 8956 469864 8968
rect 295300 8928 469864 8956
rect 295300 8916 295306 8928
rect 469858 8916 469864 8928
rect 469916 8916 469922 8968
rect 532510 8916 532516 8968
rect 532568 8956 532574 8968
rect 566090 8956 566096 8968
rect 532568 8928 566096 8956
rect 532568 8916 532574 8928
rect 566090 8916 566096 8928
rect 566148 8916 566154 8968
rect 400122 8304 400128 8356
rect 400180 8344 400186 8356
rect 404538 8344 404544 8356
rect 400180 8316 404544 8344
rect 400180 8304 400186 8316
rect 404538 8304 404544 8316
rect 404596 8304 404602 8356
rect 89162 8168 89168 8220
rect 89220 8208 89226 8220
rect 184198 8208 184204 8220
rect 89220 8180 184204 8208
rect 89220 8168 89226 8180
rect 184198 8168 184204 8180
rect 184256 8168 184262 8220
rect 85666 8100 85672 8152
rect 85724 8140 85730 8152
rect 182818 8140 182824 8152
rect 85724 8112 182824 8140
rect 85724 8100 85730 8112
rect 182818 8100 182824 8112
rect 182876 8100 182882 8152
rect 421558 8100 421564 8152
rect 421616 8140 421622 8152
rect 456886 8140 456892 8152
rect 421616 8112 456892 8140
rect 421616 8100 421622 8112
rect 456886 8100 456892 8112
rect 456944 8100 456950 8152
rect 45462 8032 45468 8084
rect 45520 8072 45526 8084
rect 141418 8072 141424 8084
rect 45520 8044 141424 8072
rect 45520 8032 45526 8044
rect 141418 8032 141424 8044
rect 141476 8032 141482 8084
rect 446398 8032 446404 8084
rect 446456 8072 446462 8084
rect 549070 8072 549076 8084
rect 446456 8044 549076 8072
rect 446456 8032 446462 8044
rect 549070 8032 549076 8044
rect 549128 8032 549134 8084
rect 38378 7964 38384 8016
rect 38436 8004 38442 8016
rect 138658 8004 138664 8016
rect 38436 7976 138664 8004
rect 38436 7964 38442 7976
rect 138658 7964 138664 7976
rect 138716 7964 138722 8016
rect 382366 7964 382372 8016
rect 382424 8004 382430 8016
rect 400490 8004 400496 8016
rect 382424 7976 400496 8004
rect 382424 7964 382430 7976
rect 400490 7964 400496 7976
rect 400548 7964 400554 8016
rect 447962 7964 447968 8016
rect 448020 8004 448026 8016
rect 552658 8004 552664 8016
rect 448020 7976 552664 8004
rect 448020 7964 448026 7976
rect 552658 7964 552664 7976
rect 552716 7964 552722 8016
rect 78582 7896 78588 7948
rect 78640 7936 78646 7948
rect 181438 7936 181444 7948
rect 78640 7908 181444 7936
rect 78640 7896 78646 7908
rect 181438 7896 181444 7908
rect 181496 7896 181502 7948
rect 378870 7896 378876 7948
rect 378928 7936 378934 7948
rect 398926 7936 398932 7948
rect 378928 7908 398932 7936
rect 378928 7896 378934 7908
rect 398926 7896 398932 7908
rect 398984 7896 398990 7948
rect 447778 7896 447784 7948
rect 447836 7936 447842 7948
rect 556154 7936 556160 7948
rect 447836 7908 556160 7936
rect 447836 7896 447842 7908
rect 556154 7896 556160 7908
rect 556212 7896 556218 7948
rect 71498 7828 71504 7880
rect 71556 7868 71562 7880
rect 178678 7868 178684 7880
rect 71556 7840 178684 7868
rect 71556 7828 71562 7840
rect 178678 7828 178684 7840
rect 178736 7828 178742 7880
rect 368198 7828 368204 7880
rect 368256 7868 368262 7880
rect 396166 7868 396172 7880
rect 368256 7840 396172 7868
rect 368256 7828 368262 7840
rect 396166 7828 396172 7840
rect 396224 7828 396230 7880
rect 417418 7828 417424 7880
rect 417476 7868 417482 7880
rect 442626 7868 442632 7880
rect 417476 7840 442632 7868
rect 417476 7828 417482 7840
rect 442626 7828 442632 7840
rect 442684 7828 442690 7880
rect 450538 7828 450544 7880
rect 450596 7868 450602 7880
rect 563238 7868 563244 7880
rect 450596 7840 563244 7868
rect 450596 7828 450602 7840
rect 563238 7828 563244 7840
rect 563296 7828 563302 7880
rect 64322 7760 64328 7812
rect 64380 7800 64386 7812
rect 177298 7800 177304 7812
rect 64380 7772 177304 7800
rect 64380 7760 64386 7772
rect 177298 7760 177304 7772
rect 177356 7760 177362 7812
rect 234338 7760 234344 7812
rect 234396 7800 234402 7812
rect 246390 7800 246396 7812
rect 234396 7772 246396 7800
rect 234396 7760 234402 7772
rect 246390 7760 246396 7772
rect 246448 7760 246454 7812
rect 364610 7760 364616 7812
rect 364668 7800 364674 7812
rect 394878 7800 394884 7812
rect 364668 7772 394884 7800
rect 364668 7760 364674 7772
rect 394878 7760 394884 7772
rect 394936 7760 394942 7812
rect 417602 7760 417608 7812
rect 417660 7800 417666 7812
rect 446214 7800 446220 7812
rect 417660 7772 446220 7800
rect 417660 7760 417666 7772
rect 446214 7760 446220 7772
rect 446272 7760 446278 7812
rect 450722 7760 450728 7812
rect 450780 7800 450786 7812
rect 566826 7800 566832 7812
rect 450780 7772 566832 7800
rect 450780 7760 450786 7772
rect 566826 7760 566832 7772
rect 566884 7760 566890 7812
rect 60826 7692 60832 7744
rect 60884 7732 60890 7744
rect 175918 7732 175924 7744
rect 60884 7704 175924 7732
rect 60884 7692 60890 7704
rect 175918 7692 175924 7704
rect 175976 7692 175982 7744
rect 226426 7692 226432 7744
rect 226484 7732 226490 7744
rect 357710 7732 357716 7744
rect 226484 7704 357716 7732
rect 226484 7692 226490 7704
rect 357710 7692 357716 7704
rect 357768 7692 357774 7744
rect 361114 7692 361120 7744
rect 361172 7732 361178 7744
rect 395062 7732 395068 7744
rect 361172 7704 395068 7732
rect 361172 7692 361178 7704
rect 395062 7692 395068 7704
rect 395120 7692 395126 7744
rect 418798 7692 418804 7744
rect 418856 7732 418862 7744
rect 449802 7732 449808 7744
rect 418856 7704 449808 7732
rect 418856 7692 418862 7704
rect 449802 7692 449808 7704
rect 449860 7692 449866 7744
rect 451918 7692 451924 7744
rect 451976 7732 451982 7744
rect 570322 7732 570328 7744
rect 451976 7704 570328 7732
rect 451976 7692 451982 7704
rect 570322 7692 570328 7704
rect 570380 7692 570386 7744
rect 53742 7624 53748 7676
rect 53800 7664 53806 7676
rect 174538 7664 174544 7676
rect 53800 7636 174544 7664
rect 53800 7624 53806 7636
rect 174538 7624 174544 7636
rect 174596 7624 174602 7676
rect 237282 7624 237288 7676
rect 237340 7664 237346 7676
rect 257062 7664 257068 7676
rect 237340 7636 257068 7664
rect 237340 7624 237346 7636
rect 257062 7624 257068 7636
rect 257120 7624 257126 7676
rect 281166 7624 281172 7676
rect 281224 7664 281230 7676
rect 420178 7664 420184 7676
rect 281224 7636 420184 7664
rect 281224 7624 281230 7636
rect 420178 7624 420184 7636
rect 420236 7624 420242 7676
rect 420270 7624 420276 7676
rect 420328 7664 420334 7676
rect 453298 7664 453304 7676
rect 420328 7636 453304 7664
rect 420328 7624 420334 7636
rect 453298 7624 453304 7636
rect 453356 7624 453362 7676
rect 453390 7624 453396 7676
rect 453448 7664 453454 7676
rect 573910 7664 573916 7676
rect 453448 7636 573916 7664
rect 453448 7624 453454 7636
rect 573910 7624 573916 7636
rect 573968 7624 573974 7676
rect 9950 7556 9956 7608
rect 10008 7596 10014 7608
rect 163498 7596 163504 7608
rect 10008 7568 163504 7596
rect 10008 7556 10014 7568
rect 163498 7556 163504 7568
rect 163556 7556 163562 7608
rect 182542 7556 182548 7608
rect 182600 7596 182606 7608
rect 215938 7596 215944 7608
rect 182600 7568 215944 7596
rect 182600 7556 182606 7568
rect 215938 7556 215944 7568
rect 215996 7556 216002 7608
rect 241422 7556 241428 7608
rect 241480 7596 241486 7608
rect 274818 7596 274824 7608
rect 241480 7568 274824 7596
rect 241480 7556 241486 7568
rect 274818 7556 274824 7568
rect 274876 7556 274882 7608
rect 282822 7556 282828 7608
rect 282880 7596 282886 7608
rect 423766 7596 423772 7608
rect 282880 7568 423772 7596
rect 282880 7556 282886 7568
rect 423766 7556 423772 7568
rect 423824 7556 423830 7608
rect 454678 7556 454684 7608
rect 454736 7596 454742 7608
rect 577406 7596 577412 7608
rect 454736 7568 577412 7596
rect 454736 7556 454742 7568
rect 577406 7556 577412 7568
rect 577464 7556 577470 7608
rect 365714 7488 365720 7540
rect 365772 7528 365778 7540
rect 367002 7528 367008 7540
rect 365772 7500 367008 7528
rect 365772 7488 365778 7500
rect 367002 7488 367008 7500
rect 367060 7488 367066 7540
rect 325602 6740 325608 6792
rect 325660 6780 325666 6792
rect 383746 6780 383752 6792
rect 325660 6752 383752 6780
rect 325660 6740 325666 6752
rect 383746 6740 383752 6752
rect 383804 6740 383810 6792
rect 255222 6672 255228 6724
rect 255280 6712 255286 6724
rect 324406 6712 324412 6724
rect 255280 6684 324412 6712
rect 255280 6672 255286 6684
rect 324406 6672 324412 6684
rect 324464 6672 324470 6724
rect 105722 6604 105728 6656
rect 105780 6644 105786 6656
rect 157978 6644 157984 6656
rect 105780 6616 157984 6644
rect 105780 6604 105786 6616
rect 157978 6604 157984 6616
rect 158036 6604 158042 6656
rect 256602 6604 256608 6656
rect 256660 6644 256666 6656
rect 327994 6644 328000 6656
rect 256660 6616 328000 6644
rect 256660 6604 256666 6616
rect 327994 6604 328000 6616
rect 328052 6604 328058 6656
rect 329190 6604 329196 6656
rect 329248 6644 329254 6656
rect 385034 6644 385040 6656
rect 329248 6616 385040 6644
rect 329248 6604 329254 6616
rect 385034 6604 385040 6616
rect 385092 6604 385098 6656
rect 73798 6536 73804 6588
rect 73856 6576 73862 6588
rect 148502 6576 148508 6588
rect 73856 6548 148508 6576
rect 73856 6536 73862 6548
rect 148502 6536 148508 6548
rect 148560 6536 148566 6588
rect 257706 6536 257712 6588
rect 257764 6576 257770 6588
rect 331582 6576 331588 6588
rect 257764 6548 331588 6576
rect 257764 6536 257770 6548
rect 331582 6536 331588 6548
rect 331640 6536 331646 6588
rect 332686 6536 332692 6588
rect 332744 6576 332750 6588
rect 386506 6576 386512 6588
rect 332744 6548 386512 6576
rect 332744 6536 332750 6548
rect 386506 6536 386512 6548
rect 386564 6536 386570 6588
rect 428458 6536 428464 6588
rect 428516 6576 428522 6588
rect 481726 6576 481732 6588
rect 428516 6548 481732 6576
rect 428516 6536 428522 6548
rect 481726 6536 481732 6548
rect 481784 6536 481790 6588
rect 70302 6468 70308 6520
rect 70360 6508 70366 6520
rect 148318 6508 148324 6520
rect 70360 6480 148324 6508
rect 70360 6468 70366 6480
rect 148318 6468 148324 6480
rect 148376 6468 148382 6520
rect 257890 6468 257896 6520
rect 257948 6508 257954 6520
rect 335078 6508 335084 6520
rect 257948 6480 335084 6508
rect 257948 6468 257954 6480
rect 335078 6468 335084 6480
rect 335136 6468 335142 6520
rect 336274 6468 336280 6520
rect 336332 6508 336338 6520
rect 388162 6508 388168 6520
rect 336332 6480 388168 6508
rect 336332 6468 336338 6480
rect 388162 6468 388168 6480
rect 388220 6468 388226 6520
rect 389450 6468 389456 6520
rect 389508 6508 389514 6520
rect 401686 6508 401692 6520
rect 389508 6480 401692 6508
rect 389508 6468 389514 6480
rect 401686 6468 401692 6480
rect 401744 6468 401750 6520
rect 410518 6468 410524 6520
rect 410576 6508 410582 6520
rect 417878 6508 417884 6520
rect 410576 6480 417884 6508
rect 410576 6468 410582 6480
rect 417878 6468 417884 6480
rect 417936 6468 417942 6520
rect 428642 6468 428648 6520
rect 428700 6508 428706 6520
rect 485222 6508 485228 6520
rect 428700 6480 485228 6508
rect 428700 6468 428706 6480
rect 485222 6468 485228 6480
rect 485280 6468 485286 6520
rect 110506 6400 110512 6452
rect 110564 6440 110570 6452
rect 189718 6440 189724 6452
rect 110564 6412 189724 6440
rect 110564 6400 110570 6412
rect 189718 6400 189724 6412
rect 189776 6400 189782 6452
rect 259362 6400 259368 6452
rect 259420 6440 259426 6452
rect 338666 6440 338672 6452
rect 259420 6412 338672 6440
rect 259420 6400 259426 6412
rect 338666 6400 338672 6412
rect 338724 6400 338730 6452
rect 339862 6400 339868 6452
rect 339920 6440 339926 6452
rect 387978 6440 387984 6452
rect 339920 6412 387984 6440
rect 339920 6400 339926 6412
rect 387978 6400 387984 6412
rect 388036 6400 388042 6452
rect 412082 6400 412088 6452
rect 412140 6440 412146 6452
rect 421374 6440 421380 6452
rect 412140 6412 421380 6440
rect 412140 6400 412146 6412
rect 421374 6400 421380 6412
rect 421432 6400 421438 6452
rect 429838 6400 429844 6452
rect 429896 6440 429902 6452
rect 488810 6440 488816 6452
rect 429896 6412 488816 6440
rect 429896 6400 429902 6412
rect 488810 6400 488816 6412
rect 488868 6400 488874 6452
rect 66714 6332 66720 6384
rect 66772 6372 66778 6384
rect 146938 6372 146944 6384
rect 66772 6344 146944 6372
rect 66772 6332 66778 6344
rect 146938 6332 146944 6344
rect 146996 6332 147002 6384
rect 260466 6332 260472 6384
rect 260524 6372 260530 6384
rect 342162 6372 342168 6384
rect 260524 6344 342168 6372
rect 260524 6332 260530 6344
rect 342162 6332 342168 6344
rect 342220 6332 342226 6384
rect 343358 6332 343364 6384
rect 343416 6372 343422 6384
rect 389174 6372 389180 6384
rect 343416 6344 389180 6372
rect 343416 6332 343422 6344
rect 389174 6332 389180 6344
rect 389232 6332 389238 6384
rect 393038 6332 393044 6384
rect 393096 6372 393102 6384
rect 402974 6372 402980 6384
rect 393096 6344 402980 6372
rect 393096 6332 393102 6344
rect 402974 6332 402980 6344
rect 403032 6332 403038 6384
rect 411990 6332 411996 6384
rect 412048 6372 412054 6384
rect 424962 6372 424968 6384
rect 412048 6344 424968 6372
rect 412048 6332 412054 6344
rect 424962 6332 424968 6344
rect 425020 6332 425026 6384
rect 431402 6332 431408 6384
rect 431460 6372 431466 6384
rect 492306 6372 492312 6384
rect 431460 6344 492312 6372
rect 431460 6332 431466 6344
rect 492306 6332 492312 6344
rect 492364 6332 492370 6384
rect 63218 6264 63224 6316
rect 63276 6304 63282 6316
rect 145558 6304 145564 6316
rect 63276 6276 145564 6304
rect 63276 6264 63282 6276
rect 145558 6264 145564 6276
rect 145616 6264 145622 6316
rect 260650 6264 260656 6316
rect 260708 6304 260714 6316
rect 345750 6304 345756 6316
rect 260708 6276 345756 6304
rect 260708 6264 260714 6276
rect 345750 6264 345756 6276
rect 345808 6264 345814 6316
rect 385954 6264 385960 6316
rect 386012 6304 386018 6316
rect 400306 6304 400312 6316
rect 386012 6276 400312 6304
rect 386012 6264 386018 6276
rect 400306 6264 400312 6276
rect 400364 6264 400370 6316
rect 413278 6264 413284 6316
rect 413336 6304 413342 6316
rect 428458 6304 428464 6316
rect 413336 6276 428464 6304
rect 413336 6264 413342 6276
rect 428458 6264 428464 6276
rect 428516 6264 428522 6316
rect 431218 6264 431224 6316
rect 431276 6304 431282 6316
rect 495894 6304 495900 6316
rect 431276 6276 495900 6304
rect 431276 6264 431282 6276
rect 495894 6264 495900 6276
rect 495952 6264 495958 6316
rect 59630 6196 59636 6248
rect 59688 6236 59694 6248
rect 144178 6236 144184 6248
rect 59688 6208 144184 6236
rect 59688 6196 59694 6208
rect 144178 6196 144184 6208
rect 144236 6196 144242 6248
rect 157794 6196 157800 6248
rect 157852 6236 157858 6248
rect 209038 6236 209044 6248
rect 157852 6208 209044 6236
rect 157852 6196 157858 6208
rect 209038 6196 209044 6208
rect 209096 6196 209102 6248
rect 233142 6196 233148 6248
rect 233200 6236 233206 6248
rect 242986 6236 242992 6248
rect 233200 6208 242992 6236
rect 233200 6196 233206 6208
rect 242986 6196 242992 6208
rect 243044 6196 243050 6248
rect 263502 6196 263508 6248
rect 263560 6236 263566 6248
rect 352834 6236 352840 6248
rect 263560 6208 352840 6236
rect 263560 6196 263566 6208
rect 352834 6196 352840 6208
rect 352892 6196 352898 6248
rect 354030 6196 354036 6248
rect 354088 6236 354094 6248
rect 391934 6236 391940 6248
rect 354088 6208 391940 6236
rect 354088 6196 354094 6208
rect 391934 6196 391940 6208
rect 391992 6196 391998 6248
rect 414842 6196 414848 6248
rect 414900 6236 414906 6248
rect 432046 6236 432052 6248
rect 414900 6208 432052 6236
rect 414900 6196 414906 6208
rect 432046 6196 432052 6208
rect 432104 6196 432110 6248
rect 432598 6196 432604 6248
rect 432656 6236 432662 6248
rect 499390 6236 499396 6248
rect 432656 6208 499396 6236
rect 432656 6196 432662 6208
rect 499390 6196 499396 6208
rect 499448 6196 499454 6248
rect 103330 6128 103336 6180
rect 103388 6168 103394 6180
rect 188338 6168 188344 6180
rect 103388 6140 188344 6168
rect 103388 6128 103394 6140
rect 188338 6128 188344 6140
rect 188396 6128 188402 6180
rect 203886 6128 203892 6180
rect 203944 6168 203950 6180
rect 221458 6168 221464 6180
rect 203944 6140 221464 6168
rect 203944 6128 203950 6140
rect 221458 6128 221464 6140
rect 221516 6128 221522 6180
rect 234522 6128 234528 6180
rect 234580 6168 234586 6180
rect 249978 6168 249984 6180
rect 234580 6140 249984 6168
rect 234580 6128 234586 6140
rect 249978 6128 249984 6140
rect 250036 6128 250042 6180
rect 264606 6128 264612 6180
rect 264664 6168 264670 6180
rect 356330 6168 356336 6180
rect 264664 6140 356336 6168
rect 264664 6128 264670 6140
rect 356330 6128 356336 6140
rect 356388 6128 356394 6180
rect 357526 6128 357532 6180
rect 357584 6168 357590 6180
rect 393406 6168 393412 6180
rect 357584 6140 393412 6168
rect 357584 6128 357590 6140
rect 393406 6128 393412 6140
rect 393464 6128 393470 6180
rect 414658 6128 414664 6180
rect 414716 6168 414722 6180
rect 435542 6168 435548 6180
rect 414716 6140 435548 6168
rect 414716 6128 414722 6140
rect 435542 6128 435548 6140
rect 435600 6128 435606 6180
rect 436738 6128 436744 6180
rect 436796 6168 436802 6180
rect 513558 6168 513564 6180
rect 436796 6140 513564 6168
rect 436796 6128 436802 6140
rect 513558 6128 513564 6140
rect 513616 6128 513622 6180
rect 514754 6128 514760 6180
rect 514812 6168 514818 6180
rect 560294 6168 560300 6180
rect 514812 6140 560300 6168
rect 514812 6128 514818 6140
rect 560294 6128 560300 6140
rect 560352 6128 560358 6180
rect 409230 5584 409236 5636
rect 409288 5624 409294 5636
rect 414290 5624 414296 5636
rect 409288 5596 414296 5624
rect 409288 5584 409294 5596
rect 414290 5584 414296 5596
rect 414348 5584 414354 5636
rect 221550 5516 221556 5568
rect 221608 5556 221614 5568
rect 227162 5556 227168 5568
rect 221608 5528 227168 5556
rect 221608 5516 221614 5528
rect 227162 5516 227168 5528
rect 227220 5516 227226 5568
rect 403618 5516 403624 5568
rect 403676 5556 403682 5568
rect 405826 5556 405832 5568
rect 403676 5528 405832 5556
rect 403676 5516 403682 5528
rect 405826 5516 405832 5528
rect 405884 5516 405890 5568
rect 407758 5516 407764 5568
rect 407816 5556 407822 5568
rect 410794 5556 410800 5568
rect 407816 5528 410800 5556
rect 407816 5516 407822 5528
rect 410794 5516 410800 5528
rect 410852 5516 410858 5568
rect 122282 5312 122288 5364
rect 122340 5352 122346 5364
rect 130378 5352 130384 5364
rect 122340 5324 130384 5352
rect 122340 5312 122346 5324
rect 130378 5312 130384 5324
rect 130436 5312 130442 5364
rect 504174 5312 504180 5364
rect 504232 5352 504238 5364
rect 557626 5352 557632 5364
rect 504232 5324 557632 5352
rect 504232 5312 504238 5324
rect 557626 5312 557632 5324
rect 557684 5312 557690 5364
rect 123478 5244 123484 5296
rect 123536 5284 123542 5296
rect 162118 5284 162124 5296
rect 123536 5256 162124 5284
rect 123536 5244 123542 5256
rect 162118 5244 162124 5256
rect 162176 5244 162182 5296
rect 500586 5244 500592 5296
rect 500644 5284 500650 5296
rect 556246 5284 556252 5296
rect 500644 5256 556252 5284
rect 500644 5244 500650 5256
rect 556246 5244 556252 5256
rect 556304 5244 556310 5296
rect 119890 5176 119896 5228
rect 119948 5216 119954 5228
rect 160738 5216 160744 5228
rect 119948 5188 160744 5216
rect 119948 5176 119954 5188
rect 160738 5176 160744 5188
rect 160796 5176 160802 5228
rect 497090 5176 497096 5228
rect 497148 5216 497154 5228
rect 556430 5216 556436 5228
rect 497148 5188 556436 5216
rect 497148 5176 497154 5188
rect 556430 5176 556436 5188
rect 556488 5176 556494 5228
rect 116394 5108 116400 5160
rect 116452 5148 116458 5160
rect 160922 5148 160928 5160
rect 116452 5120 160928 5148
rect 116452 5108 116458 5120
rect 160922 5108 160928 5120
rect 160980 5108 160986 5160
rect 196802 5108 196808 5160
rect 196860 5148 196866 5160
rect 220078 5148 220084 5160
rect 196860 5120 220084 5148
rect 196860 5108 196866 5120
rect 220078 5108 220084 5120
rect 220136 5108 220142 5160
rect 246942 5108 246948 5160
rect 247000 5148 247006 5160
rect 292574 5148 292580 5160
rect 247000 5120 292580 5148
rect 247000 5108 247006 5120
rect 292574 5108 292580 5120
rect 292632 5108 292638 5160
rect 493502 5108 493508 5160
rect 493560 5148 493566 5160
rect 554866 5148 554872 5160
rect 493560 5120 554872 5148
rect 493560 5108 493566 5120
rect 554866 5108 554872 5120
rect 554924 5108 554930 5160
rect 112806 5040 112812 5092
rect 112864 5080 112870 5092
rect 159358 5080 159364 5092
rect 112864 5052 159364 5080
rect 112864 5040 112870 5052
rect 159358 5040 159364 5052
rect 159416 5040 159422 5092
rect 193306 5040 193312 5092
rect 193364 5080 193370 5092
rect 218698 5080 218704 5092
rect 193364 5052 218704 5080
rect 193364 5040 193370 5052
rect 218698 5040 218704 5052
rect 218756 5040 218762 5092
rect 249702 5040 249708 5092
rect 249760 5080 249766 5092
rect 303154 5080 303160 5092
rect 249760 5052 303160 5080
rect 249760 5040 249766 5052
rect 303154 5040 303160 5052
rect 303212 5040 303218 5092
rect 362218 5040 362224 5092
rect 362276 5080 362282 5092
rect 374178 5080 374184 5092
rect 362276 5052 374184 5080
rect 362276 5040 362282 5052
rect 374178 5040 374184 5052
rect 374236 5040 374242 5092
rect 489914 5040 489920 5092
rect 489972 5080 489978 5092
rect 553486 5080 553492 5092
rect 489972 5052 553492 5080
rect 489972 5040 489978 5052
rect 553486 5040 553492 5052
rect 553544 5040 553550 5092
rect 98638 4972 98644 5024
rect 98696 5012 98702 5024
rect 155218 5012 155224 5024
rect 98696 4984 155224 5012
rect 98696 4972 98702 4984
rect 155218 4972 155224 4984
rect 155276 4972 155282 5024
rect 189718 4972 189724 5024
rect 189776 5012 189782 5024
rect 217318 5012 217324 5024
rect 189776 4984 217324 5012
rect 189776 4972 189782 4984
rect 217318 4972 217324 4984
rect 217376 4972 217382 5024
rect 250990 4972 250996 5024
rect 251048 5012 251054 5024
rect 306742 5012 306748 5024
rect 251048 4984 306748 5012
rect 251048 4972 251054 4984
rect 306742 4972 306748 4984
rect 306800 4972 306806 5024
rect 315022 4972 315028 5024
rect 315080 5012 315086 5024
rect 381078 5012 381084 5024
rect 315080 4984 362356 5012
rect 315080 4972 315086 4984
rect 118786 4904 118792 4956
rect 118844 4944 118850 4956
rect 129182 4944 129188 4956
rect 118844 4916 129188 4944
rect 118844 4904 118850 4916
rect 129182 4904 129188 4916
rect 129240 4904 129246 4956
rect 147122 4904 147128 4956
rect 147180 4944 147186 4956
rect 206278 4944 206284 4956
rect 147180 4916 206284 4944
rect 147180 4904 147186 4916
rect 206278 4904 206284 4916
rect 206336 4904 206342 4956
rect 218146 4904 218152 4956
rect 218204 4944 218210 4956
rect 225598 4944 225604 4956
rect 218204 4916 225604 4944
rect 218204 4904 218210 4916
rect 225598 4904 225604 4916
rect 225656 4904 225662 4956
rect 245562 4904 245568 4956
rect 245620 4944 245626 4956
rect 288986 4944 288992 4956
rect 245620 4916 288992 4944
rect 245620 4904 245626 4916
rect 288986 4904 288992 4916
rect 289044 4904 289050 4956
rect 290182 4904 290188 4956
rect 290240 4944 290246 4956
rect 362218 4944 362224 4956
rect 290240 4916 362224 4944
rect 290240 4904 290246 4916
rect 362218 4904 362224 4916
rect 362276 4904 362282 4956
rect 362328 4944 362356 4984
rect 367066 4984 381084 5012
rect 367066 4944 367094 4984
rect 381078 4972 381084 4984
rect 381136 4972 381142 5024
rect 486418 4972 486424 5024
rect 486476 5012 486482 5024
rect 553670 5012 553676 5024
rect 486476 4984 553676 5012
rect 486476 4972 486482 4984
rect 553670 4972 553676 4984
rect 553728 4972 553734 5024
rect 362328 4916 367094 4944
rect 425606 4904 425612 4956
rect 425664 4944 425670 4956
rect 474550 4944 474556 4956
rect 425664 4916 474556 4944
rect 425664 4904 425670 4916
rect 474550 4904 474556 4916
rect 474608 4904 474614 4956
rect 482830 4904 482836 4956
rect 482888 4944 482894 4956
rect 552014 4944 552020 4956
rect 482888 4916 552020 4944
rect 482888 4904 482894 4916
rect 552014 4904 552020 4916
rect 552072 4904 552078 4956
rect 115198 4836 115204 4888
rect 115256 4876 115262 4888
rect 128998 4876 129004 4888
rect 115256 4848 129004 4876
rect 115256 4836 115262 4848
rect 128998 4836 129004 4848
rect 129056 4836 129062 4888
rect 143626 4836 143632 4888
rect 143684 4876 143690 4888
rect 205174 4876 205180 4888
rect 143684 4848 205180 4876
rect 143684 4836 143690 4848
rect 205174 4836 205180 4848
rect 205232 4836 205238 4888
rect 250806 4836 250812 4888
rect 250864 4876 250870 4888
rect 310238 4876 310244 4888
rect 250864 4848 310244 4876
rect 250864 4836 250870 4848
rect 310238 4836 310244 4848
rect 310296 4836 310302 4888
rect 537202 4876 537208 4888
rect 316006 4848 537208 4876
rect 12342 4768 12348 4820
rect 12400 4808 12406 4820
rect 101398 4808 101404 4820
rect 12400 4780 101404 4808
rect 12400 4768 12406 4780
rect 101398 4768 101404 4780
rect 101456 4768 101462 4820
rect 111610 4768 111616 4820
rect 111668 4808 111674 4820
rect 127618 4808 127624 4820
rect 111668 4780 127624 4808
rect 111668 4768 111674 4780
rect 127618 4768 127624 4780
rect 127676 4768 127682 4820
rect 140038 4768 140044 4820
rect 140096 4808 140102 4820
rect 204898 4808 204904 4820
rect 140096 4780 204904 4808
rect 140096 4768 140102 4780
rect 204898 4768 204904 4780
rect 204956 4768 204962 4820
rect 207382 4768 207388 4820
rect 207440 4808 207446 4820
rect 222838 4808 222844 4820
rect 207440 4780 222844 4808
rect 207440 4768 207446 4780
rect 222838 4768 222844 4780
rect 222896 4768 222902 4820
rect 231486 4768 231492 4820
rect 231544 4808 231550 4820
rect 239306 4808 239312 4820
rect 231544 4780 239312 4808
rect 231544 4768 231550 4780
rect 239306 4768 239312 4780
rect 239364 4768 239370 4820
rect 313826 4808 313832 4820
rect 258046 4780 313832 4808
rect 214466 4700 214472 4752
rect 214524 4740 214530 4752
rect 224218 4740 224224 4752
rect 214524 4712 224224 4740
rect 214524 4700 214530 4712
rect 224218 4700 224224 4712
rect 224276 4700 224282 4752
rect 252462 4700 252468 4752
rect 252520 4740 252526 4752
rect 258046 4740 258074 4780
rect 313826 4768 313832 4780
rect 313884 4768 313890 4820
rect 314470 4768 314476 4820
rect 314528 4808 314534 4820
rect 316006 4808 316034 4848
rect 537202 4836 537208 4848
rect 537260 4836 537266 4888
rect 540790 4808 540796 4820
rect 314528 4780 316034 4808
rect 325666 4780 540796 4808
rect 314528 4768 314534 4780
rect 252520 4712 258074 4740
rect 252520 4700 252526 4712
rect 314286 4700 314292 4752
rect 314344 4740 314350 4752
rect 325666 4740 325694 4780
rect 540790 4768 540796 4780
rect 540848 4768 540854 4820
rect 314344 4712 325694 4740
rect 314344 4700 314350 4712
rect 231670 4224 231676 4276
rect 231728 4264 231734 4276
rect 235810 4264 235816 4276
rect 231728 4236 235816 4264
rect 231728 4224 231734 4236
rect 235810 4224 235816 4236
rect 235868 4224 235874 4276
rect 225138 4156 225144 4208
rect 225196 4196 225202 4208
rect 226978 4196 226984 4208
rect 225196 4168 226984 4196
rect 225196 4156 225202 4168
rect 226978 4156 226984 4168
rect 227036 4156 227042 4208
rect 230382 4156 230388 4208
rect 230440 4196 230446 4208
rect 232222 4196 232228 4208
rect 230440 4168 232228 4196
rect 230440 4156 230446 4168
rect 232222 4156 232228 4168
rect 232280 4156 232286 4208
rect 46658 4088 46664 4140
rect 46716 4128 46722 4140
rect 172054 4128 172060 4140
rect 46716 4100 172060 4128
rect 46716 4088 46722 4100
rect 172054 4088 172060 4100
rect 172112 4088 172118 4140
rect 348050 4088 348056 4140
rect 348108 4128 348114 4140
rect 356698 4128 356704 4140
rect 348108 4100 356704 4128
rect 348108 4088 348114 4100
rect 356698 4088 356704 4100
rect 356756 4088 356762 4140
rect 468662 4088 468668 4140
rect 468720 4128 468726 4140
rect 548058 4128 548064 4140
rect 468720 4100 548064 4128
rect 468720 4088 468726 4100
rect 548058 4088 548064 4100
rect 548116 4088 548122 4140
rect 43070 4020 43076 4072
rect 43128 4060 43134 4072
rect 171778 4060 171784 4072
rect 43128 4032 171784 4060
rect 43128 4020 43134 4032
rect 171778 4020 171784 4032
rect 171836 4020 171842 4072
rect 465166 4020 465172 4072
rect 465224 4060 465230 4072
rect 546586 4060 546592 4072
rect 465224 4032 546592 4060
rect 465224 4020 465230 4032
rect 546586 4020 546592 4032
rect 546644 4020 546650 4072
rect 39574 3952 39580 4004
rect 39632 3992 39638 4004
rect 170398 3992 170404 4004
rect 39632 3964 170404 3992
rect 39632 3952 39638 3964
rect 170398 3952 170404 3964
rect 170456 3952 170462 4004
rect 461578 3952 461584 4004
rect 461636 3992 461642 4004
rect 546770 3992 546776 4004
rect 461636 3964 546776 3992
rect 461636 3952 461642 3964
rect 546770 3952 546776 3964
rect 546828 3952 546834 4004
rect 35986 3884 35992 3936
rect 36044 3924 36050 3936
rect 169018 3924 169024 3936
rect 36044 3896 169024 3924
rect 36044 3884 36050 3896
rect 169018 3884 169024 3896
rect 169076 3884 169082 3936
rect 458082 3884 458088 3936
rect 458140 3924 458146 3936
rect 545206 3924 545212 3936
rect 458140 3896 545212 3924
rect 458140 3884 458146 3896
rect 545206 3884 545212 3896
rect 545264 3884 545270 3936
rect 564434 3884 564440 3936
rect 564492 3924 564498 3936
rect 574094 3924 574100 3936
rect 564492 3896 574100 3924
rect 564492 3884 564498 3896
rect 574094 3884 574100 3896
rect 574152 3884 574158 3936
rect 32398 3816 32404 3868
rect 32456 3856 32462 3868
rect 167822 3856 167828 3868
rect 32456 3828 167828 3856
rect 32456 3816 32462 3828
rect 167822 3816 167828 3828
rect 167880 3816 167886 3868
rect 337470 3816 337476 3868
rect 337528 3856 337534 3868
rect 345658 3856 345664 3868
rect 337528 3828 345664 3856
rect 337528 3816 337534 3828
rect 345658 3816 345664 3828
rect 345716 3816 345722 3868
rect 454494 3816 454500 3868
rect 454552 3856 454558 3868
rect 543826 3856 543832 3868
rect 454552 3828 543832 3856
rect 454552 3816 454558 3828
rect 543826 3816 543832 3828
rect 543884 3816 543890 3868
rect 560846 3816 560852 3868
rect 560904 3856 560910 3868
rect 573082 3856 573088 3868
rect 560904 3828 573088 3856
rect 560904 3816 560910 3828
rect 573082 3816 573088 3828
rect 573140 3816 573146 3868
rect 28902 3748 28908 3800
rect 28960 3788 28966 3800
rect 167638 3788 167644 3800
rect 28960 3760 167644 3788
rect 28960 3748 28966 3760
rect 167638 3748 167644 3760
rect 167696 3748 167702 3800
rect 198182 3788 198188 3800
rect 180766 3760 198188 3788
rect 25314 3680 25320 3732
rect 25372 3720 25378 3732
rect 180766 3720 180794 3760
rect 198182 3748 198188 3760
rect 198240 3748 198246 3800
rect 326798 3748 326804 3800
rect 326856 3788 326862 3800
rect 342898 3788 342904 3800
rect 326856 3760 342904 3788
rect 326856 3748 326862 3760
rect 342898 3748 342904 3760
rect 342956 3748 342962 3800
rect 382918 3788 382924 3800
rect 373966 3760 382924 3788
rect 196618 3720 196624 3732
rect 25372 3692 180794 3720
rect 190748 3692 196624 3720
rect 25372 3680 25378 3692
rect 20622 3612 20628 3664
rect 20680 3652 20686 3664
rect 190748 3652 190776 3692
rect 196618 3680 196624 3692
rect 196676 3680 196682 3732
rect 330386 3680 330392 3732
rect 330444 3720 330450 3732
rect 348418 3720 348424 3732
rect 330444 3692 348424 3720
rect 330444 3680 330450 3692
rect 348418 3680 348424 3692
rect 348476 3680 348482 3732
rect 358722 3680 358728 3732
rect 358780 3720 358786 3732
rect 370498 3720 370504 3732
rect 358780 3692 370504 3720
rect 358780 3680 358786 3692
rect 370498 3680 370504 3692
rect 370556 3680 370562 3732
rect 372890 3680 372896 3732
rect 372948 3720 372954 3732
rect 373966 3720 373994 3760
rect 382918 3748 382924 3760
rect 382976 3748 382982 3800
rect 415486 3748 415492 3800
rect 415544 3788 415550 3800
rect 443638 3788 443644 3800
rect 415544 3760 443644 3788
rect 415544 3748 415550 3760
rect 443638 3748 443644 3760
rect 443696 3748 443702 3800
rect 447410 3748 447416 3800
rect 447468 3788 447474 3800
rect 542354 3788 542360 3800
rect 447468 3760 542360 3788
rect 447468 3748 447474 3760
rect 542354 3748 542360 3760
rect 542412 3748 542418 3800
rect 557350 3748 557356 3800
rect 557408 3788 557414 3800
rect 572898 3788 572904 3800
rect 557408 3760 572904 3788
rect 557408 3748 557414 3760
rect 572898 3748 572904 3760
rect 572956 3748 572962 3800
rect 372948 3692 373994 3720
rect 372948 3680 372954 3692
rect 376478 3680 376484 3732
rect 376536 3720 376542 3732
rect 392578 3720 392584 3732
rect 376536 3692 392584 3720
rect 376536 3680 376542 3692
rect 392578 3680 392584 3692
rect 392636 3680 392642 3732
rect 443822 3680 443828 3732
rect 443880 3720 443886 3732
rect 541066 3720 541072 3732
rect 443880 3692 541072 3720
rect 443880 3680 443886 3692
rect 541066 3680 541072 3692
rect 541124 3680 541130 3732
rect 553762 3680 553768 3732
rect 553820 3720 553826 3732
rect 571334 3720 571340 3732
rect 553820 3692 571340 3720
rect 553820 3680 553826 3692
rect 571334 3680 571340 3692
rect 571392 3680 571398 3732
rect 195238 3652 195244 3664
rect 20680 3624 190776 3652
rect 191116 3624 195244 3652
rect 20680 3612 20686 3624
rect 15930 3544 15936 3596
rect 15988 3584 15994 3596
rect 191116 3584 191144 3624
rect 195238 3612 195244 3624
rect 195296 3612 195302 3664
rect 319714 3612 319720 3664
rect 319772 3652 319778 3664
rect 340138 3652 340144 3664
rect 319772 3624 340144 3652
rect 319772 3612 319778 3624
rect 340138 3612 340144 3624
rect 340196 3612 340202 3664
rect 351638 3612 351644 3664
rect 351696 3652 351702 3664
rect 364978 3652 364984 3664
rect 351696 3624 364984 3652
rect 351696 3612 351702 3624
rect 364978 3612 364984 3624
rect 365036 3612 365042 3664
rect 365806 3612 365812 3664
rect 365864 3652 365870 3664
rect 378778 3652 378784 3664
rect 365864 3624 378784 3652
rect 365864 3612 365870 3624
rect 378778 3612 378784 3624
rect 378836 3612 378842 3664
rect 390646 3612 390652 3664
rect 390704 3652 390710 3664
rect 404998 3652 405004 3664
rect 390704 3624 405004 3652
rect 390704 3612 390710 3624
rect 404998 3612 405004 3624
rect 405056 3612 405062 3664
rect 408402 3612 408408 3664
rect 408460 3652 408466 3664
rect 425790 3652 425796 3664
rect 408460 3624 425796 3652
rect 408460 3612 408466 3624
rect 425790 3612 425796 3624
rect 425848 3612 425854 3664
rect 440326 3612 440332 3664
rect 440384 3652 440390 3664
rect 539686 3652 539692 3664
rect 440384 3624 539692 3652
rect 440384 3612 440390 3624
rect 539686 3612 539692 3624
rect 539744 3612 539750 3664
rect 550266 3612 550272 3664
rect 550324 3652 550330 3664
rect 570046 3652 570052 3664
rect 550324 3624 570052 3652
rect 550324 3612 550330 3624
rect 570046 3612 570052 3624
rect 570104 3612 570110 3664
rect 193858 3584 193864 3596
rect 15988 3556 191144 3584
rect 191208 3556 193864 3584
rect 15988 3544 15994 3556
rect 4062 3476 4068 3528
rect 4120 3516 4126 3528
rect 4798 3516 4804 3528
rect 4120 3488 4804 3516
rect 4120 3476 4126 3488
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 8754 3476 8760 3528
rect 8812 3516 8818 3528
rect 10318 3516 10324 3528
rect 8812 3488 10324 3516
rect 8812 3476 8818 3488
rect 10318 3476 10324 3488
rect 10376 3476 10382 3528
rect 13538 3476 13544 3528
rect 13596 3516 13602 3528
rect 14458 3516 14464 3528
rect 13596 3488 14464 3516
rect 13596 3476 13602 3488
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 14734 3476 14740 3528
rect 14792 3516 14798 3528
rect 15838 3516 15844 3528
rect 14792 3488 15844 3516
rect 14792 3476 14798 3488
rect 15838 3476 15844 3488
rect 15896 3476 15902 3528
rect 191208 3516 191236 3556
rect 193858 3544 193864 3556
rect 193916 3544 193922 3596
rect 226334 3544 226340 3596
rect 226392 3584 226398 3596
rect 227530 3584 227536 3596
rect 226392 3556 227536 3584
rect 226392 3544 226398 3556
rect 227530 3544 227536 3556
rect 227588 3544 227594 3596
rect 248782 3544 248788 3596
rect 248840 3584 248846 3596
rect 253198 3584 253204 3596
rect 248840 3556 253204 3584
rect 248840 3544 248846 3556
rect 253198 3544 253204 3556
rect 253256 3544 253262 3596
rect 262858 3584 262864 3596
rect 258046 3556 262864 3584
rect 16040 3488 191236 3516
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 3418 3448 3424 3460
rect 624 3420 3424 3448
rect 624 3408 630 3420
rect 3418 3408 3424 3420
rect 3476 3408 3482 3460
rect 5258 3408 5264 3460
rect 5316 3448 5322 3460
rect 5316 3420 6914 3448
rect 5316 3408 5322 3420
rect 6886 3312 6914 3420
rect 11146 3340 11152 3392
rect 11204 3380 11210 3392
rect 16040 3380 16068 3488
rect 193214 3476 193220 3528
rect 193272 3516 193278 3528
rect 194410 3516 194416 3528
rect 193272 3488 194416 3516
rect 193272 3476 193278 3488
rect 194410 3476 194416 3488
rect 194468 3476 194474 3528
rect 218054 3476 218060 3528
rect 218112 3516 218118 3528
rect 219250 3516 219256 3528
rect 218112 3488 219256 3516
rect 218112 3476 218118 3488
rect 219250 3476 219256 3488
rect 219308 3476 219314 3528
rect 242894 3476 242900 3528
rect 242952 3516 242958 3528
rect 244090 3516 244096 3528
rect 242952 3488 244096 3516
rect 242952 3476 242958 3488
rect 244090 3476 244096 3488
rect 244148 3476 244154 3528
rect 255866 3476 255872 3528
rect 255924 3516 255930 3528
rect 258046 3516 258074 3556
rect 262858 3544 262864 3556
rect 262916 3544 262922 3596
rect 284294 3544 284300 3596
rect 284352 3584 284358 3596
rect 285030 3584 285036 3596
rect 284352 3556 285036 3584
rect 284352 3544 284358 3556
rect 285030 3544 285036 3556
rect 285088 3544 285094 3596
rect 309042 3544 309048 3596
rect 309100 3584 309106 3596
rect 331950 3584 331956 3596
rect 309100 3556 331956 3584
rect 309100 3544 309106 3556
rect 331950 3544 331956 3556
rect 332008 3544 332014 3596
rect 344554 3544 344560 3596
rect 344612 3584 344618 3596
rect 360838 3584 360844 3596
rect 344612 3556 360844 3584
rect 344612 3544 344618 3556
rect 360838 3544 360844 3556
rect 360896 3544 360902 3596
rect 378962 3584 378968 3596
rect 373966 3556 378968 3584
rect 255924 3488 258074 3516
rect 255924 3476 255930 3488
rect 259454 3476 259460 3528
rect 259512 3516 259518 3528
rect 260650 3516 260656 3528
rect 259512 3488 260656 3516
rect 259512 3476 259518 3488
rect 260650 3476 260656 3488
rect 260708 3476 260714 3528
rect 299474 3476 299480 3528
rect 299532 3516 299538 3528
rect 300762 3516 300768 3528
rect 299532 3488 300768 3516
rect 299532 3476 299538 3488
rect 300762 3476 300768 3488
rect 300820 3476 300826 3528
rect 301958 3476 301964 3528
rect 302016 3516 302022 3528
rect 329098 3516 329104 3528
rect 302016 3488 329104 3516
rect 302016 3476 302022 3488
rect 329098 3476 329104 3488
rect 329156 3476 329162 3528
rect 333882 3476 333888 3528
rect 333940 3516 333946 3528
rect 333940 3488 345014 3516
rect 333940 3476 333946 3488
rect 197998 3448 198004 3460
rect 11204 3352 16068 3380
rect 16546 3420 198004 3448
rect 11204 3340 11210 3352
rect 16546 3312 16574 3420
rect 197998 3408 198004 3420
rect 198056 3408 198062 3460
rect 238110 3408 238116 3460
rect 238168 3448 238174 3460
rect 242158 3448 242164 3460
rect 238168 3420 242164 3448
rect 238168 3408 238174 3420
rect 242158 3408 242164 3420
rect 242216 3408 242222 3460
rect 262950 3408 262956 3460
rect 263008 3448 263014 3460
rect 302878 3448 302884 3460
rect 263008 3420 302884 3448
rect 263008 3408 263014 3420
rect 302878 3408 302884 3420
rect 302936 3408 302942 3460
rect 312630 3408 312636 3460
rect 312688 3448 312694 3460
rect 338758 3448 338764 3460
rect 312688 3420 338764 3448
rect 312688 3408 312694 3420
rect 338758 3408 338764 3420
rect 338816 3408 338822 3460
rect 344986 3448 345014 3488
rect 349246 3476 349252 3528
rect 349304 3516 349310 3528
rect 350442 3516 350448 3528
rect 349304 3488 350448 3516
rect 349304 3476 349310 3488
rect 350442 3476 350448 3488
rect 350500 3476 350506 3528
rect 362310 3476 362316 3528
rect 362368 3516 362374 3528
rect 373966 3516 373994 3556
rect 378962 3544 378968 3556
rect 379020 3544 379026 3596
rect 390554 3544 390560 3596
rect 390612 3584 390618 3596
rect 391842 3584 391848 3596
rect 390612 3556 391848 3584
rect 390612 3544 390618 3556
rect 391842 3544 391848 3556
rect 391900 3544 391906 3596
rect 397730 3544 397736 3596
rect 397788 3584 397794 3596
rect 418890 3584 418896 3596
rect 397788 3556 418896 3584
rect 397788 3544 397794 3556
rect 418890 3544 418896 3556
rect 418948 3544 418954 3596
rect 436738 3544 436744 3596
rect 436796 3584 436802 3596
rect 539870 3584 539876 3596
rect 436796 3556 539876 3584
rect 436796 3544 436802 3556
rect 539870 3544 539876 3556
rect 539928 3544 539934 3596
rect 546678 3544 546684 3596
rect 546736 3584 546742 3596
rect 570230 3584 570236 3596
rect 546736 3556 570236 3584
rect 546736 3544 546742 3556
rect 570230 3544 570236 3556
rect 570288 3544 570294 3596
rect 362368 3488 373994 3516
rect 362368 3476 362374 3488
rect 374086 3476 374092 3528
rect 374144 3516 374150 3528
rect 375282 3516 375288 3528
rect 374144 3488 375288 3516
rect 374144 3476 374150 3488
rect 375282 3476 375288 3488
rect 375340 3476 375346 3528
rect 379974 3476 379980 3528
rect 380032 3516 380038 3528
rect 403526 3516 403532 3528
rect 380032 3488 403532 3516
rect 380032 3476 380038 3488
rect 403526 3476 403532 3488
rect 403584 3476 403590 3528
rect 404814 3476 404820 3528
rect 404872 3516 404878 3528
rect 429930 3516 429936 3528
rect 404872 3488 429936 3516
rect 404872 3476 404878 3488
rect 429930 3476 429936 3488
rect 429988 3476 429994 3528
rect 433242 3476 433248 3528
rect 433300 3516 433306 3528
rect 538306 3516 538312 3528
rect 433300 3488 538312 3516
rect 433300 3476 433306 3488
rect 538306 3476 538312 3488
rect 538364 3476 538370 3528
rect 543182 3476 543188 3528
rect 543240 3516 543246 3528
rect 568758 3516 568764 3528
rect 543240 3488 568764 3516
rect 543240 3476 543246 3488
rect 568758 3476 568764 3488
rect 568816 3476 568822 3528
rect 575106 3476 575112 3528
rect 575164 3516 575170 3528
rect 576946 3516 576952 3528
rect 575164 3488 576952 3516
rect 575164 3476 575170 3488
rect 576946 3476 576952 3488
rect 577004 3476 577010 3528
rect 353938 3448 353944 3460
rect 344986 3420 353944 3448
rect 353938 3408 353944 3420
rect 353996 3408 354002 3460
rect 355226 3408 355232 3460
rect 355284 3448 355290 3460
rect 376018 3448 376024 3460
rect 355284 3420 376024 3448
rect 355284 3408 355290 3420
rect 376018 3408 376024 3420
rect 376076 3408 376082 3460
rect 383562 3408 383568 3460
rect 383620 3448 383626 3460
rect 410610 3448 410616 3460
rect 383620 3420 410616 3448
rect 383620 3408 383626 3420
rect 410610 3408 410616 3420
rect 410668 3408 410674 3460
rect 415394 3408 415400 3460
rect 415452 3448 415458 3460
rect 416682 3448 416688 3460
rect 415452 3420 416688 3448
rect 415452 3408 415458 3420
rect 416682 3408 416688 3420
rect 416740 3408 416746 3460
rect 422570 3408 422576 3460
rect 422628 3448 422634 3460
rect 535454 3448 535460 3460
rect 422628 3420 535460 3448
rect 422628 3408 422634 3420
rect 535454 3408 535460 3420
rect 535512 3408 535518 3460
rect 539594 3408 539600 3460
rect 539652 3448 539658 3460
rect 567194 3448 567200 3460
rect 539652 3420 567200 3448
rect 539652 3408 539658 3420
rect 567194 3408 567200 3420
rect 567252 3408 567258 3460
rect 574738 3408 574744 3460
rect 574796 3448 574802 3460
rect 576302 3448 576308 3460
rect 574796 3420 576308 3448
rect 574796 3408 574802 3420
rect 576302 3408 576308 3420
rect 576360 3408 576366 3460
rect 117590 3340 117596 3392
rect 117648 3380 117654 3392
rect 191098 3380 191104 3392
rect 117648 3352 191104 3380
rect 117648 3340 117654 3352
rect 191098 3340 191104 3352
rect 191156 3340 191162 3392
rect 259454 3340 259460 3392
rect 259512 3380 259518 3392
rect 266998 3380 267004 3392
rect 259512 3352 267004 3380
rect 259512 3340 259518 3352
rect 266998 3340 267004 3352
rect 267056 3340 267062 3392
rect 316034 3340 316040 3392
rect 316092 3380 316098 3392
rect 317322 3380 317328 3392
rect 316092 3352 317328 3380
rect 316092 3340 316098 3352
rect 317322 3340 317328 3352
rect 317380 3340 317386 3392
rect 440234 3340 440240 3392
rect 440292 3380 440298 3392
rect 441522 3380 441528 3392
rect 440292 3352 441528 3380
rect 440292 3340 440298 3352
rect 441522 3340 441528 3352
rect 441580 3340 441586 3392
rect 472250 3340 472256 3392
rect 472308 3380 472314 3392
rect 549530 3380 549536 3392
rect 472308 3352 549536 3380
rect 472308 3340 472314 3352
rect 549530 3340 549536 3352
rect 549588 3340 549594 3392
rect 568022 3340 568028 3392
rect 568080 3380 568086 3392
rect 575750 3380 575756 3392
rect 568080 3352 575756 3380
rect 568080 3340 568086 3352
rect 575750 3340 575756 3352
rect 575808 3340 575814 3392
rect 6886 3284 16574 3312
rect 121086 3272 121092 3324
rect 121144 3312 121150 3324
rect 192478 3312 192484 3324
rect 121144 3284 192484 3312
rect 121144 3272 121150 3284
rect 192478 3272 192484 3284
rect 192536 3272 192542 3324
rect 252370 3272 252376 3324
rect 252428 3312 252434 3324
rect 255958 3312 255964 3324
rect 252428 3284 255964 3312
rect 252428 3272 252434 3284
rect 255958 3272 255964 3284
rect 256016 3272 256022 3324
rect 475746 3272 475752 3324
rect 475804 3312 475810 3324
rect 549346 3312 549352 3324
rect 475804 3284 549352 3312
rect 475804 3272 475810 3284
rect 549346 3272 549352 3284
rect 549404 3272 549410 3324
rect 580258 3272 580264 3324
rect 580316 3312 580322 3324
rect 580994 3312 581000 3324
rect 580316 3284 581000 3312
rect 580316 3272 580322 3284
rect 580994 3272 581000 3284
rect 581052 3272 581058 3324
rect 124674 3204 124680 3256
rect 124732 3244 124738 3256
rect 194042 3244 194048 3256
rect 124732 3216 194048 3244
rect 124732 3204 124738 3216
rect 194042 3204 194048 3216
rect 194100 3204 194106 3256
rect 479334 3204 479340 3256
rect 479392 3244 479398 3256
rect 550726 3244 550732 3256
rect 479392 3216 550732 3244
rect 479392 3204 479398 3216
rect 550726 3204 550732 3216
rect 550784 3204 550790 3256
rect 143534 3136 143540 3188
rect 143592 3176 143598 3188
rect 144730 3176 144736 3188
rect 143592 3148 144736 3176
rect 143592 3136 143598 3148
rect 144730 3136 144736 3148
rect 144788 3136 144794 3188
rect 536098 3136 536104 3188
rect 536156 3176 536162 3188
rect 565906 3176 565912 3188
rect 536156 3148 565912 3176
rect 536156 3136 536162 3148
rect 565906 3136 565912 3148
rect 565964 3136 565970 3188
rect 571518 3000 571524 3052
rect 571576 3040 571582 3052
rect 575566 3040 575572 3052
rect 571576 3012 575572 3040
rect 571576 3000 571582 3012
rect 575566 3000 575572 3012
rect 575624 3000 575630 3052
rect 2866 2864 2872 2916
rect 2924 2904 2930 2916
rect 4890 2904 4896 2916
rect 2924 2876 4896 2904
rect 2924 2864 2930 2876
rect 4890 2864 4896 2876
rect 4948 2864 4954 2916
<< via1 >>
rect 256608 49784 256660 49836
rect 257804 49784 257856 49836
rect 351828 49784 351880 49836
rect 353300 49784 353352 49836
rect 3424 49716 3476 49768
rect 98000 49716 98052 49768
rect 299480 49240 299532 49292
rect 375380 49240 375432 49292
rect 436468 49240 436520 49292
rect 520280 49240 520332 49292
rect 150440 49172 150492 49224
rect 208124 49172 208176 49224
rect 282736 49172 282788 49224
rect 412640 49172 412692 49224
rect 78680 49104 78732 49156
rect 118608 49104 118660 49156
rect 197360 49104 197412 49156
rect 346400 49104 346452 49156
rect 378784 49104 378836 49156
rect 517704 49104 517756 49156
rect 92480 49036 92532 49088
rect 184848 49036 184900 49088
rect 246948 49036 247000 49088
rect 281540 49036 281592 49088
rect 311716 49036 311768 49088
rect 518900 49036 518952 49088
rect 6920 48968 6972 49020
rect 99380 48968 99432 49020
rect 198740 48968 198792 49020
rect 470600 48968 470652 49020
rect 521752 48968 521804 49020
rect 560392 48968 560444 49020
rect 346400 47880 346452 47932
rect 387800 47880 387852 47932
rect 276020 47812 276072 47864
rect 368756 47812 368808 47864
rect 286324 47744 286376 47796
rect 426440 47744 426492 47796
rect 434628 47744 434680 47796
rect 502432 47744 502484 47796
rect 190460 47676 190512 47728
rect 345020 47676 345072 47728
rect 382924 47676 382976 47728
rect 519176 47676 519228 47728
rect 93860 47608 93912 47660
rect 122472 47608 122524 47660
rect 200120 47608 200172 47660
rect 221832 47608 221884 47660
rect 242716 47608 242768 47660
rect 267740 47608 267792 47660
rect 304908 47608 304960 47660
rect 494060 47608 494112 47660
rect 1400 47540 1452 47592
rect 99656 47540 99708 47592
rect 138020 47540 138072 47592
rect 454408 47540 454460 47592
rect 510620 47540 510672 47592
rect 557632 47540 557684 47592
rect 396080 46928 396132 46980
rect 402980 46928 403032 46980
rect 282920 46452 282972 46504
rect 369860 46452 369912 46504
rect 277308 46384 277360 46436
rect 405740 46384 405792 46436
rect 201500 46316 201552 46368
rect 348148 46316 348200 46368
rect 371240 46316 371292 46368
rect 394700 46316 394752 46368
rect 416688 46316 416740 46368
rect 438860 46316 438912 46368
rect 445668 46316 445720 46368
rect 540980 46316 541032 46368
rect 46940 46248 46992 46300
rect 109040 46248 109092 46300
rect 246764 46248 246816 46300
rect 284300 46248 284352 46300
rect 315948 46248 316000 46300
rect 543740 46248 543792 46300
rect 80060 46180 80112 46232
rect 150532 46180 150584 46232
rect 175280 46180 175332 46232
rect 214932 46180 214984 46232
rect 253204 46180 253256 46232
rect 484584 46180 484636 46232
rect 321560 45160 321612 45212
rect 383936 45160 383988 45212
rect 278688 45092 278740 45144
rect 408500 45092 408552 45144
rect 329104 45024 329156 45076
rect 502340 45024 502392 45076
rect 297916 44956 297968 45008
rect 476120 44956 476172 45008
rect 53840 44888 53892 44940
rect 112628 44888 112680 44940
rect 154580 44888 154632 44940
rect 333428 44888 333480 44940
rect 418896 44888 418948 44940
rect 528560 44888 528612 44940
rect 93952 44820 94004 44872
rect 155408 44820 155460 44872
rect 168380 44820 168432 44872
rect 211804 44820 211856 44872
rect 248236 44820 248288 44872
rect 295340 44820 295392 44872
rect 319996 44820 320048 44872
rect 557540 44820 557592 44872
rect 310520 43732 310572 43784
rect 380900 43732 380952 43784
rect 262128 43664 262180 43716
rect 349160 43664 349212 43716
rect 286876 43596 286928 43648
rect 440240 43596 440292 43648
rect 443644 43596 443696 43648
rect 532700 43596 532752 43648
rect 129740 43528 129792 43580
rect 326528 43528 326580 43580
rect 348424 43528 348476 43580
rect 509332 43528 509384 43580
rect 60740 43460 60792 43512
rect 113824 43460 113876 43512
rect 319812 43460 319864 43512
rect 561680 43460 561732 43512
rect 67640 43392 67692 43444
rect 177488 43392 177540 43444
rect 219440 43392 219492 43444
rect 480352 43392 480404 43444
rect 307760 42372 307812 42424
rect 379520 42372 379572 42424
rect 284024 42304 284076 42356
rect 430580 42304 430632 42356
rect 204260 42236 204312 42288
rect 352012 42236 352064 42288
rect 429936 42236 429988 42288
rect 530216 42236 530268 42288
rect 64880 42168 64932 42220
rect 115388 42168 115440 42220
rect 342904 42168 342956 42220
rect 509516 42168 509568 42220
rect 106280 42100 106332 42152
rect 188528 42100 188580 42152
rect 253756 42100 253808 42152
rect 320180 42100 320232 42152
rect 321468 42100 321520 42152
rect 564440 42100 564492 42152
rect 34520 42032 34572 42084
rect 138848 42032 138900 42084
rect 194600 42032 194652 42084
rect 473360 42032 473412 42084
rect 349252 41012 349304 41064
rect 390744 41012 390796 41064
rect 264796 40944 264848 40996
rect 358820 40944 358872 40996
rect 215300 40876 215352 40928
rect 354864 40876 354916 40928
rect 376024 40876 376076 40928
rect 516324 40876 516376 40928
rect 75920 40808 75972 40860
rect 117964 40808 118016 40860
rect 289728 40808 289780 40860
rect 448520 40808 448572 40860
rect 113180 40740 113232 40792
rect 191288 40740 191340 40792
rect 318708 40740 318760 40792
rect 554780 40740 554832 40792
rect 27620 40672 27672 40724
rect 135904 40672 135956 40724
rect 241520 40672 241572 40724
rect 485780 40672 485832 40724
rect 292580 39652 292632 39704
rect 375380 39652 375432 39704
rect 277308 39584 277360 39636
rect 401600 39584 401652 39636
rect 186320 39516 186372 39568
rect 346492 39516 346544 39568
rect 403624 39516 403676 39568
rect 523224 39516 523276 39568
rect 331956 39448 332008 39500
rect 503904 39448 503956 39500
rect 85580 39380 85632 39432
rect 120724 39380 120776 39432
rect 248052 39380 248104 39432
rect 299572 39380 299624 39432
rect 317144 39380 317196 39432
rect 550640 39380 550692 39432
rect 22100 39312 22152 39364
rect 134708 39312 134760 39364
rect 191840 39312 191892 39364
rect 471980 39312 472032 39364
rect 303620 38156 303672 38208
rect 378324 38156 378376 38208
rect 281356 38088 281408 38140
rect 415400 38088 415452 38140
rect 443736 38088 443788 38140
rect 538220 38088 538272 38140
rect 193220 38020 193272 38072
rect 347964 38020 348016 38072
rect 392584 38020 392636 38072
rect 523040 38020 523092 38072
rect 89720 37952 89772 38004
rect 122104 37952 122156 38004
rect 253572 37952 253624 38004
rect 316040 37952 316092 38004
rect 317328 37952 317380 38004
rect 547880 37952 547932 38004
rect 17960 37884 18012 37936
rect 134524 37884 134576 37936
rect 244280 37884 244332 37936
rect 487436 37884 487488 37936
rect 266268 36864 266320 36916
rect 362960 36864 363012 36916
rect 240140 36796 240192 36848
rect 361764 36796 361816 36848
rect 353944 36728 353996 36780
rect 510712 36728 510764 36780
rect 77300 36660 77352 36712
rect 149704 36660 149756 36712
rect 291016 36660 291068 36712
rect 451280 36660 451332 36712
rect 99380 36592 99432 36644
rect 186964 36592 187016 36644
rect 313188 36592 313240 36644
rect 532700 36592 532752 36644
rect 16580 36524 16632 36576
rect 101588 36524 101640 36576
rect 176660 36524 176712 36576
rect 467840 36524 467892 36576
rect 267556 35504 267608 35556
rect 369860 35504 369912 35556
rect 251180 35436 251232 35488
rect 364432 35436 364484 35488
rect 360844 35368 360896 35420
rect 513472 35368 513524 35420
rect 290832 35300 290884 35352
rect 455420 35300 455472 35352
rect 86960 35232 87012 35284
rect 152464 35232 152516 35284
rect 311808 35232 311860 35284
rect 529940 35232 529992 35284
rect 20720 35164 20772 35216
rect 102784 35164 102836 35216
rect 180800 35164 180852 35216
rect 469220 35164 469272 35216
rect 273168 34008 273220 34060
rect 387800 34008 387852 34060
rect 293776 33940 293828 33992
rect 465080 33940 465132 33992
rect 133880 33872 133932 33924
rect 326344 33872 326396 33924
rect 378876 33872 378928 33924
rect 518992 33872 519044 33924
rect 29000 33804 29052 33856
rect 105728 33804 105780 33856
rect 310244 33804 310296 33856
rect 525800 33804 525852 33856
rect 56600 33736 56652 33788
rect 174728 33736 174780 33788
rect 184940 33736 184992 33788
rect 470692 33736 470744 33788
rect 524420 33736 524472 33788
rect 563244 33736 563296 33788
rect 270224 32648 270276 32700
rect 376760 32648 376812 32700
rect 445024 32648 445076 32700
rect 545120 32648 545172 32700
rect 247040 32580 247092 32632
rect 363052 32580 363104 32632
rect 425796 32580 425848 32632
rect 531320 32580 531372 32632
rect 292488 32512 292540 32564
rect 458180 32512 458232 32564
rect 81440 32444 81492 32496
rect 181628 32444 181680 32496
rect 310428 32444 310480 32496
rect 523040 32444 523092 32496
rect 40040 32376 40092 32428
rect 108488 32376 108540 32428
rect 135260 32376 135312 32428
rect 456984 32376 457036 32428
rect 253940 31356 253992 31408
rect 364616 31356 364668 31408
rect 275928 31288 275980 31340
rect 398840 31288 398892 31340
rect 340144 31220 340196 31272
rect 506756 31220 506808 31272
rect 172520 31152 172572 31204
rect 342260 31152 342312 31204
rect 441068 31152 441120 31204
rect 531320 31152 531372 31204
rect 91100 31084 91152 31136
rect 153844 31084 153896 31136
rect 307484 31084 307536 31136
rect 514760 31084 514812 31136
rect 44180 31016 44232 31068
rect 108304 31016 108356 31068
rect 187700 31016 187752 31068
rect 470876 31016 470928 31068
rect 258080 29928 258132 29980
rect 365720 29928 365772 29980
rect 274364 29860 274416 29912
rect 394700 29860 394752 29912
rect 338764 29792 338816 29844
rect 505100 29792 505152 29844
rect 176752 29724 176804 29776
rect 343640 29724 343692 29776
rect 440884 29724 440936 29776
rect 527180 29724 527232 29776
rect 49700 29656 49752 29708
rect 173164 29656 173216 29708
rect 307668 29656 307720 29708
rect 512000 29656 512052 29708
rect 4804 29588 4856 29640
rect 131948 29588 132000 29640
rect 167000 29588 167052 29640
rect 465172 29588 465224 29640
rect 274548 28500 274600 28552
rect 390560 28500 390612 28552
rect 242900 28432 242952 28484
rect 361580 28432 361632 28484
rect 364984 28432 365036 28484
rect 516140 28432 516192 28484
rect 296628 28364 296680 28416
rect 473360 28364 473412 28416
rect 10324 28296 10376 28348
rect 131764 28296 131816 28348
rect 306288 28296 306340 28348
rect 507860 28296 507912 28348
rect 131120 28228 131172 28280
rect 455512 28228 455564 28280
rect 260840 27140 260892 27192
rect 367284 27140 367336 27192
rect 270408 27072 270460 27124
rect 380900 27072 380952 27124
rect 442264 27072 442316 27124
rect 534080 27072 534132 27124
rect 293592 27004 293644 27056
rect 462320 27004 462372 27056
rect 48320 26936 48372 26988
rect 141608 26936 141660 26988
rect 304908 26936 304960 26988
rect 505100 26936 505152 26988
rect 74540 26868 74592 26920
rect 180064 26868 180116 26920
rect 266360 26868 266412 26920
rect 492864 26868 492916 26920
rect 269028 25780 269080 25832
rect 374000 25780 374052 25832
rect 286692 25712 286744 25764
rect 437480 25712 437532 25764
rect 438124 25712 438176 25764
rect 516140 25712 516192 25764
rect 140780 25644 140832 25696
rect 329196 25644 329248 25696
rect 410616 25644 410668 25696
rect 524512 25644 524564 25696
rect 153200 25576 153252 25628
rect 207664 25576 207716 25628
rect 303344 25576 303396 25628
rect 500960 25576 501012 25628
rect 35900 25508 35952 25560
rect 106924 25508 106976 25560
rect 201592 25508 201644 25560
rect 474740 25508 474792 25560
rect 267372 24420 267424 24472
rect 365720 24420 365772 24472
rect 264980 24352 265032 24404
rect 367100 24352 367152 24404
rect 285588 24284 285640 24336
rect 433340 24284 433392 24336
rect 433984 24284 434036 24336
rect 506480 24284 506532 24336
rect 303528 24216 303580 24268
rect 498200 24216 498252 24268
rect 135352 24148 135404 24200
rect 203524 24148 203576 24200
rect 267004 24148 267056 24200
rect 490012 24148 490064 24200
rect 26240 24080 26292 24132
rect 104164 24080 104216 24132
rect 149060 24080 149112 24132
rect 461032 24080 461084 24132
rect 271788 22992 271840 23044
rect 383660 22992 383712 23044
rect 439504 22992 439556 23044
rect 523132 22992 523184 23044
rect 288348 22924 288400 22976
rect 444380 22924 444432 22976
rect 132500 22856 132552 22908
rect 202144 22856 202196 22908
rect 242808 22856 242860 22908
rect 277400 22856 277452 22908
rect 300676 22856 300728 22908
rect 489920 22856 489972 22908
rect 158720 22788 158772 22840
rect 333244 22788 333296 22840
rect 411260 22788 411312 22840
rect 532884 22788 532936 22840
rect 52460 22720 52512 22772
rect 142804 22720 142856 22772
rect 262864 22720 262916 22772
rect 490196 22720 490248 22772
rect 236000 21632 236052 21684
rect 360200 21632 360252 21684
rect 179420 21564 179472 21616
rect 345204 21564 345256 21616
rect 356704 21564 356756 21616
rect 514852 21564 514904 21616
rect 300492 21496 300544 21548
rect 487160 21496 487212 21548
rect 242164 21428 242216 21480
rect 484400 21428 484452 21480
rect 33140 21360 33192 21412
rect 105544 21360 105596 21412
rect 128360 21360 128412 21412
rect 200948 21360 201000 21412
rect 241244 21360 241296 21412
rect 270500 21360 270552 21412
rect 324136 21360 324188 21412
rect 574744 21360 574796 21412
rect 271880 20272 271932 20324
rect 369952 20272 370004 20324
rect 218060 20204 218112 20256
rect 354680 20204 354732 20256
rect 299388 20136 299440 20188
rect 483020 20136 483072 20188
rect 302884 20068 302936 20120
rect 491300 20068 491352 20120
rect 103520 20000 103572 20052
rect 125048 20000 125100 20052
rect 126980 20000 127032 20052
rect 324964 20000 325016 20052
rect 405004 20000 405056 20052
rect 526076 20000 526128 20052
rect 14464 19932 14516 19984
rect 133144 19932 133196 19984
rect 185032 19932 185084 19984
rect 217508 19932 217560 19984
rect 238484 19932 238536 19984
rect 263600 19932 263652 19984
rect 323952 19932 324004 19984
rect 572720 19932 572772 19984
rect 233240 18844 233292 18896
rect 358912 18844 358964 18896
rect 183560 18776 183612 18828
rect 345020 18776 345072 18828
rect 345664 18776 345716 18828
rect 512092 18776 512144 18828
rect 297732 18708 297784 18760
rect 480260 18708 480312 18760
rect 100760 18640 100812 18692
rect 124864 18640 124916 18692
rect 238668 18640 238720 18692
rect 259460 18640 259512 18692
rect 322848 18640 322900 18692
rect 568580 18640 568632 18692
rect 4896 18572 4948 18624
rect 98644 18572 98696 18624
rect 109040 18572 109092 18624
rect 158168 18572 158220 18624
rect 178040 18572 178092 18624
rect 214564 18572 214616 18624
rect 223580 18572 223632 18624
rect 480536 18572 480588 18624
rect 322940 17688 322992 17740
rect 507952 17688 508004 17740
rect 316132 17620 316184 17672
rect 506572 17620 506624 17672
rect 305000 17552 305052 17604
rect 503720 17552 503772 17604
rect 160100 17484 160152 17536
rect 463792 17484 463844 17536
rect 155960 17416 156012 17468
rect 462412 17416 462464 17468
rect 151820 17348 151872 17400
rect 461216 17348 461268 17400
rect 55220 17280 55272 17332
rect 144368 17280 144420 17332
rect 144920 17280 144972 17332
rect 459560 17280 459612 17332
rect 96620 17212 96672 17264
rect 123484 17212 123536 17264
rect 142160 17212 142212 17264
rect 458272 17212 458324 17264
rect 298100 16396 298152 16448
rect 501052 16396 501104 16448
rect 294880 16328 294932 16380
rect 499672 16328 499724 16380
rect 291384 16260 291436 16312
rect 499856 16260 499908 16312
rect 287336 16192 287388 16244
rect 498292 16192 498344 16244
rect 284392 16124 284444 16176
rect 497096 16124 497148 16176
rect 280712 16056 280764 16108
rect 496912 16056 496964 16108
rect 83280 15988 83332 16040
rect 119344 15988 119396 16040
rect 276664 15988 276716 16040
rect 495440 15988 495492 16040
rect 102232 15920 102284 15972
rect 156604 15920 156656 15972
rect 160652 15920 160704 15972
rect 210608 15920 210660 15972
rect 273260 15920 273312 15972
rect 494152 15920 494204 15972
rect 15844 15852 15896 15904
rect 165068 15852 165120 15904
rect 209780 15852 209832 15904
rect 224408 15852 224460 15904
rect 235908 15852 235960 15904
rect 253112 15852 253164 15904
rect 270040 15852 270092 15904
rect 492680 15852 492732 15904
rect 528560 15852 528612 15904
rect 564532 15852 564584 15904
rect 234620 14832 234672 14884
rect 483112 14832 483164 14884
rect 231032 14764 231084 14816
rect 483296 14764 483348 14816
rect 226340 14696 226392 14748
rect 481640 14696 481692 14748
rect 216864 14628 216916 14680
rect 478880 14628 478932 14680
rect 164424 14560 164476 14612
rect 210424 14560 210476 14612
rect 213368 14560 213420 14612
rect 477500 14560 477552 14612
rect 72608 14492 72660 14544
rect 116584 14492 116636 14544
rect 209872 14492 209924 14544
rect 476304 14492 476356 14544
rect 84200 14424 84252 14476
rect 151084 14424 151136 14476
rect 206192 14424 206244 14476
rect 476488 14424 476540 14476
rect 507216 14424 507268 14476
rect 559104 14424 559156 14476
rect 151912 13472 151964 13524
rect 331864 13472 331916 13524
rect 147864 13404 147916 13456
rect 330484 13404 330536 13456
rect 143540 13336 143592 13388
rect 330668 13336 330720 13388
rect 449164 13336 449216 13388
rect 559288 13336 559340 13388
rect 173900 13268 173952 13320
rect 466552 13268 466604 13320
rect 170312 13200 170364 13252
rect 466736 13200 466788 13252
rect 41880 13132 41932 13184
rect 140044 13132 140096 13184
rect 163688 13132 163740 13184
rect 463976 13132 464028 13184
rect 58440 13064 58492 13116
rect 112444 13064 112496 13116
rect 127532 13064 127584 13116
rect 454040 13064 454092 13116
rect 374092 12112 374144 12164
rect 397460 12112 397512 12164
rect 286600 11976 286652 12028
rect 374368 11976 374420 12028
rect 279056 11908 279108 11960
rect 371424 11908 371476 11960
rect 435364 11908 435416 11960
rect 509608 11908 509660 11960
rect 268384 11840 268436 11892
rect 368480 11840 368532 11892
rect 370504 11840 370556 11892
rect 517520 11840 517572 11892
rect 108120 11772 108172 11824
rect 126244 11772 126296 11824
rect 137192 11772 137244 11824
rect 327724 11772 327776 11824
rect 340972 11772 341024 11824
rect 513656 11772 513708 11824
rect 51080 11704 51132 11756
rect 111064 11704 111116 11756
rect 176660 11704 176712 11756
rect 177856 11704 177908 11756
rect 255964 11704 256016 11756
rect 488540 11704 488592 11756
rect 517888 11704 517940 11756
rect 561772 11704 561824 11756
rect 582380 11704 582432 11756
rect 583392 11704 583444 11756
rect 425520 10616 425572 10668
rect 536932 10616 536984 10668
rect 318064 10548 318116 10600
rect 382280 10548 382332 10600
rect 418528 10548 418580 10600
rect 534172 10548 534224 10600
rect 229376 10480 229428 10532
rect 357532 10480 357584 10532
rect 400220 10480 400272 10532
rect 530032 10480 530084 10532
rect 171692 10412 171744 10464
rect 213184 10412 213236 10464
rect 222752 10412 222804 10464
rect 356060 10412 356112 10464
rect 393320 10412 393372 10464
rect 527272 10412 527324 10464
rect 69112 10344 69164 10396
rect 115204 10344 115256 10396
rect 125600 10344 125652 10396
rect 200764 10344 200816 10396
rect 211712 10344 211764 10396
rect 353300 10344 353352 10396
rect 386420 10344 386472 10396
rect 525892 10344 525944 10396
rect 30840 10276 30892 10328
rect 137284 10276 137336 10328
rect 208584 10276 208636 10328
rect 352196 10276 352248 10328
rect 369400 10276 369452 10328
rect 520372 10276 520424 10328
rect 151728 9596 151780 9648
rect 153016 9596 153068 9648
rect 209688 9596 209740 9648
rect 210976 9596 211028 9648
rect 421748 9324 421800 9376
rect 460388 9324 460440 9376
rect 422944 9256 422996 9308
rect 463976 9256 464028 9308
rect 96252 9188 96304 9240
rect 185584 9188 185636 9240
rect 297272 9188 297324 9240
rect 376852 9188 376904 9240
rect 424508 9188 424560 9240
rect 467472 9188 467524 9240
rect 24216 9120 24268 9172
rect 166264 9120 166316 9172
rect 169576 9120 169628 9172
rect 336004 9120 336056 9172
rect 424324 9120 424376 9172
rect 471060 9120 471112 9172
rect 166080 9052 166132 9104
rect 336188 9052 336240 9104
rect 427084 9052 427136 9104
rect 478144 9052 478196 9104
rect 162492 8984 162544 9036
rect 334624 8984 334676 9036
rect 450912 8984 450964 9036
rect 542544 8984 542596 9036
rect 19432 8916 19484 8968
rect 164884 8916 164936 8968
rect 295248 8916 295300 8968
rect 469864 8916 469916 8968
rect 532516 8916 532568 8968
rect 566096 8916 566148 8968
rect 400128 8304 400180 8356
rect 404544 8304 404596 8356
rect 89168 8168 89220 8220
rect 184204 8168 184256 8220
rect 85672 8100 85724 8152
rect 182824 8100 182876 8152
rect 421564 8100 421616 8152
rect 456892 8100 456944 8152
rect 45468 8032 45520 8084
rect 141424 8032 141476 8084
rect 446404 8032 446456 8084
rect 549076 8032 549128 8084
rect 38384 7964 38436 8016
rect 138664 7964 138716 8016
rect 382372 7964 382424 8016
rect 400496 7964 400548 8016
rect 447968 7964 448020 8016
rect 552664 7964 552716 8016
rect 78588 7896 78640 7948
rect 181444 7896 181496 7948
rect 378876 7896 378928 7948
rect 398932 7896 398984 7948
rect 447784 7896 447836 7948
rect 556160 7896 556212 7948
rect 71504 7828 71556 7880
rect 178684 7828 178736 7880
rect 368204 7828 368256 7880
rect 396172 7828 396224 7880
rect 417424 7828 417476 7880
rect 442632 7828 442684 7880
rect 450544 7828 450596 7880
rect 563244 7828 563296 7880
rect 64328 7760 64380 7812
rect 177304 7760 177356 7812
rect 234344 7760 234396 7812
rect 246396 7760 246448 7812
rect 364616 7760 364668 7812
rect 394884 7760 394936 7812
rect 417608 7760 417660 7812
rect 446220 7760 446272 7812
rect 450728 7760 450780 7812
rect 566832 7760 566884 7812
rect 60832 7692 60884 7744
rect 175924 7692 175976 7744
rect 226432 7692 226484 7744
rect 357716 7692 357768 7744
rect 361120 7692 361172 7744
rect 395068 7692 395120 7744
rect 418804 7692 418856 7744
rect 449808 7692 449860 7744
rect 451924 7692 451976 7744
rect 570328 7692 570380 7744
rect 53748 7624 53800 7676
rect 174544 7624 174596 7676
rect 237288 7624 237340 7676
rect 257068 7624 257120 7676
rect 281172 7624 281224 7676
rect 420184 7624 420236 7676
rect 420276 7624 420328 7676
rect 453304 7624 453356 7676
rect 453396 7624 453448 7676
rect 573916 7624 573968 7676
rect 9956 7556 10008 7608
rect 163504 7556 163556 7608
rect 182548 7556 182600 7608
rect 215944 7556 215996 7608
rect 241428 7556 241480 7608
rect 274824 7556 274876 7608
rect 282828 7556 282880 7608
rect 423772 7556 423824 7608
rect 454684 7556 454736 7608
rect 577412 7556 577464 7608
rect 365720 7488 365772 7540
rect 367008 7488 367060 7540
rect 325608 6740 325660 6792
rect 383752 6740 383804 6792
rect 255228 6672 255280 6724
rect 324412 6672 324464 6724
rect 105728 6604 105780 6656
rect 157984 6604 158036 6656
rect 256608 6604 256660 6656
rect 328000 6604 328052 6656
rect 329196 6604 329248 6656
rect 385040 6604 385092 6656
rect 73804 6536 73856 6588
rect 148508 6536 148560 6588
rect 257712 6536 257764 6588
rect 331588 6536 331640 6588
rect 332692 6536 332744 6588
rect 386512 6536 386564 6588
rect 428464 6536 428516 6588
rect 481732 6536 481784 6588
rect 70308 6468 70360 6520
rect 148324 6468 148376 6520
rect 257896 6468 257948 6520
rect 335084 6468 335136 6520
rect 336280 6468 336332 6520
rect 388168 6468 388220 6520
rect 389456 6468 389508 6520
rect 401692 6468 401744 6520
rect 410524 6468 410576 6520
rect 417884 6468 417936 6520
rect 428648 6468 428700 6520
rect 485228 6468 485280 6520
rect 110512 6400 110564 6452
rect 189724 6400 189776 6452
rect 259368 6400 259420 6452
rect 338672 6400 338724 6452
rect 339868 6400 339920 6452
rect 387984 6400 388036 6452
rect 412088 6400 412140 6452
rect 421380 6400 421432 6452
rect 429844 6400 429896 6452
rect 488816 6400 488868 6452
rect 66720 6332 66772 6384
rect 146944 6332 146996 6384
rect 260472 6332 260524 6384
rect 342168 6332 342220 6384
rect 343364 6332 343416 6384
rect 389180 6332 389232 6384
rect 393044 6332 393096 6384
rect 402980 6332 403032 6384
rect 411996 6332 412048 6384
rect 424968 6332 425020 6384
rect 431408 6332 431460 6384
rect 492312 6332 492364 6384
rect 63224 6264 63276 6316
rect 145564 6264 145616 6316
rect 260656 6264 260708 6316
rect 345756 6264 345808 6316
rect 385960 6264 386012 6316
rect 400312 6264 400364 6316
rect 413284 6264 413336 6316
rect 428464 6264 428516 6316
rect 431224 6264 431276 6316
rect 495900 6264 495952 6316
rect 59636 6196 59688 6248
rect 144184 6196 144236 6248
rect 157800 6196 157852 6248
rect 209044 6196 209096 6248
rect 233148 6196 233200 6248
rect 242992 6196 243044 6248
rect 263508 6196 263560 6248
rect 352840 6196 352892 6248
rect 354036 6196 354088 6248
rect 391940 6196 391992 6248
rect 414848 6196 414900 6248
rect 432052 6196 432104 6248
rect 432604 6196 432656 6248
rect 499396 6196 499448 6248
rect 103336 6128 103388 6180
rect 188344 6128 188396 6180
rect 203892 6128 203944 6180
rect 221464 6128 221516 6180
rect 234528 6128 234580 6180
rect 249984 6128 250036 6180
rect 264612 6128 264664 6180
rect 356336 6128 356388 6180
rect 357532 6128 357584 6180
rect 393412 6128 393464 6180
rect 414664 6128 414716 6180
rect 435548 6128 435600 6180
rect 436744 6128 436796 6180
rect 513564 6128 513616 6180
rect 514760 6128 514812 6180
rect 560300 6128 560352 6180
rect 409236 5584 409288 5636
rect 414296 5584 414348 5636
rect 221556 5516 221608 5568
rect 227168 5516 227220 5568
rect 403624 5516 403676 5568
rect 405832 5516 405884 5568
rect 407764 5516 407816 5568
rect 410800 5516 410852 5568
rect 122288 5312 122340 5364
rect 130384 5312 130436 5364
rect 504180 5312 504232 5364
rect 557632 5312 557684 5364
rect 123484 5244 123536 5296
rect 162124 5244 162176 5296
rect 500592 5244 500644 5296
rect 556252 5244 556304 5296
rect 119896 5176 119948 5228
rect 160744 5176 160796 5228
rect 497096 5176 497148 5228
rect 556436 5176 556488 5228
rect 116400 5108 116452 5160
rect 160928 5108 160980 5160
rect 196808 5108 196860 5160
rect 220084 5108 220136 5160
rect 246948 5108 247000 5160
rect 292580 5108 292632 5160
rect 493508 5108 493560 5160
rect 554872 5108 554924 5160
rect 112812 5040 112864 5092
rect 159364 5040 159416 5092
rect 193312 5040 193364 5092
rect 218704 5040 218756 5092
rect 249708 5040 249760 5092
rect 303160 5040 303212 5092
rect 362224 5040 362276 5092
rect 374184 5040 374236 5092
rect 489920 5040 489972 5092
rect 553492 5040 553544 5092
rect 98644 4972 98696 5024
rect 155224 4972 155276 5024
rect 189724 4972 189776 5024
rect 217324 4972 217376 5024
rect 250996 4972 251048 5024
rect 306748 4972 306800 5024
rect 315028 4972 315080 5024
rect 118792 4904 118844 4956
rect 129188 4904 129240 4956
rect 147128 4904 147180 4956
rect 206284 4904 206336 4956
rect 218152 4904 218204 4956
rect 225604 4904 225656 4956
rect 245568 4904 245620 4956
rect 288992 4904 289044 4956
rect 290188 4904 290240 4956
rect 362224 4904 362276 4956
rect 381084 4972 381136 5024
rect 486424 4972 486476 5024
rect 553676 4972 553728 5024
rect 425612 4904 425664 4956
rect 474556 4904 474608 4956
rect 482836 4904 482888 4956
rect 552020 4904 552072 4956
rect 115204 4836 115256 4888
rect 129004 4836 129056 4888
rect 143632 4836 143684 4888
rect 205180 4836 205232 4888
rect 250812 4836 250864 4888
rect 310244 4836 310296 4888
rect 12348 4768 12400 4820
rect 101404 4768 101456 4820
rect 111616 4768 111668 4820
rect 127624 4768 127676 4820
rect 140044 4768 140096 4820
rect 204904 4768 204956 4820
rect 207388 4768 207440 4820
rect 222844 4768 222896 4820
rect 231492 4768 231544 4820
rect 239312 4768 239364 4820
rect 214472 4700 214524 4752
rect 224224 4700 224276 4752
rect 252468 4700 252520 4752
rect 313832 4768 313884 4820
rect 314476 4768 314528 4820
rect 537208 4836 537260 4888
rect 314292 4700 314344 4752
rect 540796 4768 540848 4820
rect 231676 4224 231728 4276
rect 235816 4224 235868 4276
rect 225144 4156 225196 4208
rect 226984 4156 227036 4208
rect 230388 4156 230440 4208
rect 232228 4156 232280 4208
rect 46664 4088 46716 4140
rect 172060 4088 172112 4140
rect 348056 4088 348108 4140
rect 356704 4088 356756 4140
rect 468668 4088 468720 4140
rect 548064 4088 548116 4140
rect 43076 4020 43128 4072
rect 171784 4020 171836 4072
rect 465172 4020 465224 4072
rect 546592 4020 546644 4072
rect 39580 3952 39632 4004
rect 170404 3952 170456 4004
rect 461584 3952 461636 4004
rect 546776 3952 546828 4004
rect 35992 3884 36044 3936
rect 169024 3884 169076 3936
rect 458088 3884 458140 3936
rect 545212 3884 545264 3936
rect 564440 3884 564492 3936
rect 574100 3884 574152 3936
rect 32404 3816 32456 3868
rect 167828 3816 167880 3868
rect 337476 3816 337528 3868
rect 345664 3816 345716 3868
rect 454500 3816 454552 3868
rect 543832 3816 543884 3868
rect 560852 3816 560904 3868
rect 573088 3816 573140 3868
rect 28908 3748 28960 3800
rect 167644 3748 167696 3800
rect 25320 3680 25372 3732
rect 198188 3748 198240 3800
rect 326804 3748 326856 3800
rect 342904 3748 342956 3800
rect 20628 3612 20680 3664
rect 196624 3680 196676 3732
rect 330392 3680 330444 3732
rect 348424 3680 348476 3732
rect 358728 3680 358780 3732
rect 370504 3680 370556 3732
rect 372896 3680 372948 3732
rect 382924 3748 382976 3800
rect 415492 3748 415544 3800
rect 443644 3748 443696 3800
rect 447416 3748 447468 3800
rect 542360 3748 542412 3800
rect 557356 3748 557408 3800
rect 572904 3748 572956 3800
rect 376484 3680 376536 3732
rect 392584 3680 392636 3732
rect 443828 3680 443880 3732
rect 541072 3680 541124 3732
rect 553768 3680 553820 3732
rect 571340 3680 571392 3732
rect 15936 3544 15988 3596
rect 195244 3612 195296 3664
rect 319720 3612 319772 3664
rect 340144 3612 340196 3664
rect 351644 3612 351696 3664
rect 364984 3612 365036 3664
rect 365812 3612 365864 3664
rect 378784 3612 378836 3664
rect 390652 3612 390704 3664
rect 405004 3612 405056 3664
rect 408408 3612 408460 3664
rect 425796 3612 425848 3664
rect 440332 3612 440384 3664
rect 539692 3612 539744 3664
rect 550272 3612 550324 3664
rect 570052 3612 570104 3664
rect 4068 3476 4120 3528
rect 4804 3476 4856 3528
rect 8760 3476 8812 3528
rect 10324 3476 10376 3528
rect 13544 3476 13596 3528
rect 14464 3476 14516 3528
rect 14740 3476 14792 3528
rect 15844 3476 15896 3528
rect 193864 3544 193916 3596
rect 226340 3544 226392 3596
rect 227536 3544 227588 3596
rect 248788 3544 248840 3596
rect 253204 3544 253256 3596
rect 572 3408 624 3460
rect 3424 3408 3476 3460
rect 5264 3408 5316 3460
rect 11152 3340 11204 3392
rect 193220 3476 193272 3528
rect 194416 3476 194468 3528
rect 218060 3476 218112 3528
rect 219256 3476 219308 3528
rect 242900 3476 242952 3528
rect 244096 3476 244148 3528
rect 255872 3476 255924 3528
rect 262864 3544 262916 3596
rect 284300 3544 284352 3596
rect 285036 3544 285088 3596
rect 309048 3544 309100 3596
rect 331956 3544 332008 3596
rect 344560 3544 344612 3596
rect 360844 3544 360896 3596
rect 259460 3476 259512 3528
rect 260656 3476 260708 3528
rect 299480 3476 299532 3528
rect 300768 3476 300820 3528
rect 301964 3476 302016 3528
rect 329104 3476 329156 3528
rect 333888 3476 333940 3528
rect 198004 3408 198056 3460
rect 238116 3408 238168 3460
rect 242164 3408 242216 3460
rect 262956 3408 263008 3460
rect 302884 3408 302936 3460
rect 312636 3408 312688 3460
rect 338764 3408 338816 3460
rect 349252 3476 349304 3528
rect 350448 3476 350500 3528
rect 362316 3476 362368 3528
rect 378968 3544 379020 3596
rect 390560 3544 390612 3596
rect 391848 3544 391900 3596
rect 397736 3544 397788 3596
rect 418896 3544 418948 3596
rect 436744 3544 436796 3596
rect 539876 3544 539928 3596
rect 546684 3544 546736 3596
rect 570236 3544 570288 3596
rect 374092 3476 374144 3528
rect 375288 3476 375340 3528
rect 379980 3476 380032 3528
rect 403532 3476 403584 3528
rect 404820 3476 404872 3528
rect 429936 3476 429988 3528
rect 433248 3476 433300 3528
rect 538312 3476 538364 3528
rect 543188 3476 543240 3528
rect 568764 3476 568816 3528
rect 575112 3476 575164 3528
rect 576952 3476 577004 3528
rect 353944 3408 353996 3460
rect 355232 3408 355284 3460
rect 376024 3408 376076 3460
rect 383568 3408 383620 3460
rect 410616 3408 410668 3460
rect 415400 3408 415452 3460
rect 416688 3408 416740 3460
rect 422576 3408 422628 3460
rect 535460 3408 535512 3460
rect 539600 3408 539652 3460
rect 567200 3408 567252 3460
rect 574744 3408 574796 3460
rect 576308 3408 576360 3460
rect 117596 3340 117648 3392
rect 191104 3340 191156 3392
rect 259460 3340 259512 3392
rect 267004 3340 267056 3392
rect 316040 3340 316092 3392
rect 317328 3340 317380 3392
rect 440240 3340 440292 3392
rect 441528 3340 441580 3392
rect 472256 3340 472308 3392
rect 549536 3340 549588 3392
rect 568028 3340 568080 3392
rect 575756 3340 575808 3392
rect 121092 3272 121144 3324
rect 192484 3272 192536 3324
rect 252376 3272 252428 3324
rect 255964 3272 256016 3324
rect 475752 3272 475804 3324
rect 549352 3272 549404 3324
rect 580264 3272 580316 3324
rect 581000 3272 581052 3324
rect 124680 3204 124732 3256
rect 194048 3204 194100 3256
rect 479340 3204 479392 3256
rect 550732 3204 550784 3256
rect 143540 3136 143592 3188
rect 144736 3136 144788 3188
rect 536104 3136 536156 3188
rect 565912 3136 565964 3188
rect 571524 3000 571576 3052
rect 575572 3000 575624 3052
rect 2872 2864 2924 2916
rect 4896 2864 4948 2916
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 181626 50824 181682 50833
rect 181626 50759 181682 50768
rect 449162 50824 449218 50833
rect 449162 50759 449218 50768
rect 162122 50688 162178 50697
rect 99668 50632 100004 50660
rect 99378 50280 99434 50289
rect 99378 50215 99434 50224
rect 97998 49872 98054 49881
rect 97998 49807 98054 49816
rect 98012 49774 98040 49807
rect 3424 49768 3476 49774
rect 3424 49710 3476 49716
rect 98000 49768 98052 49774
rect 98000 49710 98052 49716
rect 98642 49736 98698 49745
rect 1400 47592 1452 47598
rect 1400 47534 1452 47540
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 542 -960 654 480
rect 1412 354 1440 47534
rect 3436 3466 3464 49710
rect 98642 49671 98698 49680
rect 78680 49156 78732 49162
rect 78680 49098 78732 49104
rect 6920 49020 6972 49026
rect 6920 48962 6972 48968
rect 4804 29640 4856 29646
rect 4804 29582 4856 29588
rect 4816 3534 4844 29582
rect 4896 18624 4948 18630
rect 4896 18566 4948 18572
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 3424 3460 3476 3466
rect 3424 3402 3476 3408
rect 2872 2916 2924 2922
rect 2872 2858 2924 2864
rect 2884 480 2912 2858
rect 4080 480 4108 3470
rect 4908 2922 4936 18566
rect 6932 16574 6960 48962
rect 46940 46300 46992 46306
rect 46940 46242 46992 46248
rect 34520 42084 34572 42090
rect 34520 42026 34572 42032
rect 27620 40724 27672 40730
rect 27620 40666 27672 40672
rect 22100 39364 22152 39370
rect 22100 39306 22152 39312
rect 17960 37936 18012 37942
rect 17960 37878 18012 37884
rect 16580 36576 16632 36582
rect 16580 36518 16632 36524
rect 10324 28348 10376 28354
rect 10324 28290 10376 28296
rect 6932 16546 7696 16574
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 4896 2916 4948 2922
rect 4896 2858 4948 2864
rect 5276 480 5304 3402
rect 6458 3360 6514 3369
rect 6458 3295 6514 3304
rect 6472 480 6500 3295
rect 7668 480 7696 16546
rect 9956 7608 10008 7614
rect 9956 7550 10008 7556
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 8772 480 8800 3470
rect 9968 480 9996 7550
rect 10336 3534 10364 28290
rect 14464 19984 14516 19990
rect 14464 19926 14516 19932
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 11164 480 11192 3334
rect 12360 480 12388 4762
rect 14476 3534 14504 19926
rect 16592 16574 16620 36518
rect 16592 16546 17080 16574
rect 15844 15904 15896 15910
rect 15844 15846 15896 15852
rect 15856 3534 15884 15846
rect 15936 3596 15988 3602
rect 15936 3538 15988 3544
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 13556 480 13584 3470
rect 14752 480 14780 3470
rect 15948 480 15976 3538
rect 17052 480 17080 16546
rect 1646 354 1758 480
rect 1412 326 1758 354
rect 1646 -960 1758 326
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 37878
rect 20720 35216 20772 35222
rect 20720 35158 20772 35164
rect 20732 16574 20760 35158
rect 22112 16574 22140 39306
rect 26240 24132 26292 24138
rect 26240 24074 26292 24080
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 19432 8968 19484 8974
rect 19432 8910 19484 8916
rect 19444 480 19472 8910
rect 20628 3664 20680 3670
rect 20628 3606 20680 3612
rect 20640 480 20668 3606
rect 21836 480 21864 16546
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 24216 9172 24268 9178
rect 24216 9114 24268 9120
rect 24228 480 24256 9114
rect 25320 3732 25372 3738
rect 25320 3674 25372 3680
rect 25332 480 25360 3674
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 24074
rect 27632 16574 27660 40666
rect 29000 33856 29052 33862
rect 29000 33798 29052 33804
rect 29012 16574 29040 33798
rect 33140 21412 33192 21418
rect 33140 21354 33192 21360
rect 33152 16574 33180 21354
rect 27632 16546 27752 16574
rect 29012 16546 30144 16574
rect 33152 16546 33640 16574
rect 27724 480 27752 16546
rect 28908 3800 28960 3806
rect 28908 3742 28960 3748
rect 28920 480 28948 3742
rect 30116 480 30144 16546
rect 30840 10328 30892 10334
rect 30840 10270 30892 10276
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 354 30880 10270
rect 32404 3868 32456 3874
rect 32404 3810 32456 3816
rect 32416 480 32444 3810
rect 33612 480 33640 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31270 -960 31382 326
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34532 354 34560 42026
rect 40040 32428 40092 32434
rect 40040 32370 40092 32376
rect 35900 25560 35952 25566
rect 35900 25502 35952 25508
rect 35912 16574 35940 25502
rect 40052 16574 40080 32370
rect 44180 31068 44232 31074
rect 44180 31010 44232 31016
rect 44192 16574 44220 31010
rect 46952 16574 46980 46242
rect 53840 44940 53892 44946
rect 53840 44882 53892 44888
rect 49700 29708 49752 29714
rect 49700 29650 49752 29656
rect 48320 26988 48372 26994
rect 48320 26930 48372 26936
rect 48332 16574 48360 26930
rect 49712 16574 49740 29650
rect 52460 22772 52512 22778
rect 52460 22714 52512 22720
rect 52472 16574 52500 22714
rect 53852 16574 53880 44882
rect 60740 43512 60792 43518
rect 60740 43454 60792 43460
rect 56600 33788 56652 33794
rect 56600 33730 56652 33736
rect 55220 17332 55272 17338
rect 55220 17274 55272 17280
rect 55232 16574 55260 17274
rect 56612 16574 56640 33730
rect 60752 16574 60780 43454
rect 67640 43444 67692 43450
rect 67640 43386 67692 43392
rect 64880 42220 64932 42226
rect 64880 42162 64932 42168
rect 64892 16574 64920 42162
rect 35912 16546 36768 16574
rect 40052 16546 40264 16574
rect 44192 16546 44312 16574
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 52472 16546 52592 16574
rect 53852 16546 54984 16574
rect 55232 16546 56088 16574
rect 56612 16546 56824 16574
rect 60752 16546 61608 16574
rect 64892 16546 65104 16574
rect 35992 3936 36044 3942
rect 35992 3878 36044 3884
rect 36004 480 36032 3878
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 38384 8016 38436 8022
rect 38384 7958 38436 7964
rect 38396 480 38424 7958
rect 39580 4004 39632 4010
rect 39580 3946 39632 3952
rect 39592 480 39620 3946
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40236 354 40264 16546
rect 41880 13184 41932 13190
rect 41880 13126 41932 13132
rect 41892 480 41920 13126
rect 43076 4072 43128 4078
rect 43076 4014 43128 4020
rect 43088 480 43116 4014
rect 44284 480 44312 16546
rect 45468 8084 45520 8090
rect 45468 8026 45520 8032
rect 45480 480 45508 8026
rect 46664 4140 46716 4146
rect 46664 4082 46716 4088
rect 46676 480 46704 4082
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 51080 11756 51132 11762
rect 51080 11698 51132 11704
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51092 354 51120 11698
rect 52564 480 52592 16546
rect 53748 7676 53800 7682
rect 53748 7618 53800 7624
rect 53760 480 53788 7618
rect 54956 480 54984 16546
rect 56060 480 56088 16546
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58440 13116 58492 13122
rect 58440 13058 58492 13064
rect 58452 480 58480 13058
rect 60832 7744 60884 7750
rect 60832 7686 60884 7692
rect 59636 6248 59688 6254
rect 59636 6190 59688 6196
rect 59648 480 59676 6190
rect 60844 480 60872 7686
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61580 354 61608 16546
rect 64328 7812 64380 7818
rect 64328 7754 64380 7760
rect 63224 6316 63276 6322
rect 63224 6258 63276 6264
rect 63236 480 63264 6258
rect 64340 480 64368 7754
rect 61998 354 62110 480
rect 61580 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66720 6384 66772 6390
rect 66720 6326 66772 6332
rect 66732 480 66760 6326
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 43386
rect 75920 40860 75972 40866
rect 75920 40802 75972 40808
rect 74540 26920 74592 26926
rect 74540 26862 74592 26868
rect 74552 16574 74580 26862
rect 74552 16546 75040 16574
rect 72608 14544 72660 14550
rect 72608 14486 72660 14492
rect 69112 10396 69164 10402
rect 69112 10338 69164 10344
rect 69124 480 69152 10338
rect 71504 7880 71556 7886
rect 71504 7822 71556 7828
rect 70308 6520 70360 6526
rect 70308 6462 70360 6468
rect 70320 480 70348 6462
rect 71516 480 71544 7822
rect 72620 480 72648 14486
rect 73804 6588 73856 6594
rect 73804 6530 73856 6536
rect 73816 480 73844 6530
rect 75012 480 75040 16546
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 75932 354 75960 40802
rect 77300 36712 77352 36718
rect 77300 36654 77352 36660
rect 77312 16574 77340 36654
rect 78692 16574 78720 49098
rect 92480 49088 92532 49094
rect 92480 49030 92532 49036
rect 80060 46232 80112 46238
rect 80060 46174 80112 46180
rect 80072 16574 80100 46174
rect 85580 39432 85632 39438
rect 85580 39374 85632 39380
rect 81440 32496 81492 32502
rect 81440 32438 81492 32444
rect 81452 16574 81480 32438
rect 85592 16574 85620 39374
rect 89720 38004 89772 38010
rect 89720 37946 89772 37952
rect 86960 35284 87012 35290
rect 86960 35226 87012 35232
rect 86972 16574 87000 35226
rect 89732 16574 89760 37946
rect 91100 31136 91152 31142
rect 91100 31078 91152 31084
rect 91112 16574 91140 31078
rect 77312 16546 77432 16574
rect 78692 16546 79272 16574
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 85592 16546 86448 16574
rect 86972 16546 87552 16574
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 77404 480 77432 16546
rect 78588 7948 78640 7954
rect 78588 7890 78640 7896
rect 78600 480 78628 7890
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83280 16040 83332 16046
rect 83280 15982 83332 15988
rect 83292 480 83320 15982
rect 84200 14476 84252 14482
rect 84200 14418 84252 14424
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 14418
rect 85672 8152 85724 8158
rect 85672 8094 85724 8100
rect 85684 480 85712 8094
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 16546
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 16546
rect 89168 8220 89220 8226
rect 89168 8162 89220 8168
rect 89180 480 89208 8162
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 49030
rect 93860 47660 93912 47666
rect 93860 47602 93912 47608
rect 93872 6914 93900 47602
rect 93952 44872 94004 44878
rect 93952 44814 94004 44820
rect 93964 16574 93992 44814
rect 98656 18630 98684 49671
rect 99392 49026 99420 50215
rect 99380 49020 99432 49026
rect 99380 48962 99432 48968
rect 99668 47598 99696 50632
rect 162122 50623 162178 50632
rect 178682 50688 178738 50697
rect 178682 50623 178738 50632
rect 180706 50688 180762 50697
rect 180706 50623 180762 50632
rect 181442 50688 181498 50697
rect 181442 50623 181498 50632
rect 102782 50552 102838 50561
rect 102782 50487 102838 50496
rect 109038 50552 109094 50561
rect 109038 50487 109094 50496
rect 113822 50552 113878 50561
rect 113822 50487 113878 50496
rect 133142 50552 133198 50561
rect 133142 50487 133198 50496
rect 142802 50552 142858 50561
rect 142802 50487 142858 50496
rect 152462 50552 152518 50561
rect 152462 50487 152518 50496
rect 160742 50552 160798 50561
rect 160742 50487 160798 50496
rect 101586 50416 101642 50425
rect 101586 50351 101642 50360
rect 101402 49600 101458 49609
rect 101402 49535 101458 49544
rect 99656 47592 99708 47598
rect 99656 47534 99708 47540
rect 99380 36644 99432 36650
rect 99380 36586 99432 36592
rect 98644 18624 98696 18630
rect 98644 18566 98696 18572
rect 96620 17264 96672 17270
rect 96620 17206 96672 17212
rect 96632 16574 96660 17206
rect 99392 16574 99420 36586
rect 100760 18692 100812 18698
rect 100760 18634 100812 18640
rect 93964 16546 94728 16574
rect 96632 16546 97488 16574
rect 99392 16546 99880 16574
rect 93872 6886 93992 6914
rect 93964 480 93992 6886
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94700 354 94728 16546
rect 96252 9240 96304 9246
rect 96252 9182 96304 9188
rect 96264 480 96292 9182
rect 97460 480 97488 16546
rect 98644 5024 98696 5030
rect 98644 4966 98696 4972
rect 98656 480 98684 4966
rect 99852 480 99880 16546
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95118 -960 95230 326
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 100772 354 100800 18634
rect 101416 4826 101444 49535
rect 101600 36582 101628 50351
rect 101588 36576 101640 36582
rect 101588 36518 101640 36524
rect 102796 35222 102824 50487
rect 105910 50416 105966 50425
rect 105648 50374 105910 50402
rect 104162 49872 104218 49881
rect 104162 49807 104218 49816
rect 102784 35216 102836 35222
rect 102784 35158 102836 35164
rect 104176 24138 104204 49807
rect 105648 45554 105676 50374
rect 105910 50351 105966 50360
rect 108118 50416 108174 50425
rect 108118 50351 108174 50360
rect 108302 50416 108358 50425
rect 108302 50351 108358 50360
rect 106922 50280 106978 50289
rect 106922 50215 106978 50224
rect 105726 49736 105782 49745
rect 105726 49671 105782 49680
rect 105556 45526 105676 45554
rect 104164 24132 104216 24138
rect 104164 24074 104216 24080
rect 105556 21418 105584 45526
rect 105740 33862 105768 49671
rect 106280 42152 106332 42158
rect 106280 42094 106332 42100
rect 105728 33856 105780 33862
rect 105728 33798 105780 33804
rect 105544 21412 105596 21418
rect 105544 21354 105596 21360
rect 103520 20052 103572 20058
rect 103520 19994 103572 20000
rect 103532 16574 103560 19994
rect 106292 16574 106320 42094
rect 106936 25566 106964 50215
rect 108132 50153 108160 50351
rect 108118 50144 108174 50153
rect 108118 50079 108174 50088
rect 108316 31074 108344 50351
rect 108486 49736 108542 49745
rect 108486 49671 108542 49680
rect 108500 32434 108528 49671
rect 109052 46306 109080 50487
rect 112442 50416 112498 50425
rect 112442 50351 112498 50360
rect 111062 49872 111118 49881
rect 111062 49807 111118 49816
rect 109040 46300 109092 46306
rect 109040 46242 109092 46248
rect 108488 32428 108540 32434
rect 108488 32370 108540 32376
rect 108304 31068 108356 31074
rect 108304 31010 108356 31016
rect 106924 25560 106976 25566
rect 106924 25502 106976 25508
rect 109040 18624 109092 18630
rect 109040 18566 109092 18572
rect 103532 16546 104112 16574
rect 106292 16546 106504 16574
rect 102232 15972 102284 15978
rect 102232 15914 102284 15920
rect 101404 4820 101456 4826
rect 101404 4762 101456 4768
rect 102244 480 102272 15914
rect 103336 6180 103388 6186
rect 103336 6122 103388 6128
rect 103348 480 103376 6122
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105728 6656 105780 6662
rect 105728 6598 105780 6604
rect 105740 480 105768 6598
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108120 11824 108172 11830
rect 108120 11766 108172 11772
rect 108132 480 108160 11766
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109052 354 109080 18566
rect 111076 11762 111104 49807
rect 112456 13122 112484 50351
rect 112626 49736 112682 49745
rect 112626 49671 112682 49680
rect 112640 44946 112668 49671
rect 112628 44940 112680 44946
rect 112628 44882 112680 44888
rect 113836 43518 113864 50487
rect 119342 50416 119398 50425
rect 119342 50351 119398 50360
rect 123482 50416 123538 50425
rect 123482 50351 123538 50360
rect 131762 50416 131818 50425
rect 131762 50351 131818 50360
rect 116674 50280 116730 50289
rect 116596 50238 116674 50266
rect 115202 49872 115258 49881
rect 115202 49807 115258 49816
rect 113824 43512 113876 43518
rect 113824 43454 113876 43460
rect 113180 40792 113232 40798
rect 113180 40734 113232 40740
rect 113192 16574 113220 40734
rect 113192 16546 114048 16574
rect 112444 13116 112496 13122
rect 112444 13058 112496 13064
rect 111064 11756 111116 11762
rect 111064 11698 111116 11704
rect 110512 6452 110564 6458
rect 110512 6394 110564 6400
rect 110524 480 110552 6394
rect 112812 5092 112864 5098
rect 112812 5034 112864 5040
rect 111616 4820 111668 4826
rect 111616 4762 111668 4768
rect 111628 480 111656 4762
rect 112824 480 112852 5034
rect 114020 480 114048 16546
rect 115216 10402 115244 49807
rect 115386 49736 115442 49745
rect 115386 49671 115442 49680
rect 115400 42226 115428 49671
rect 115388 42220 115440 42226
rect 115388 42162 115440 42168
rect 116596 14550 116624 50238
rect 116674 50215 116730 50224
rect 116674 50008 116730 50017
rect 116674 49943 116730 49952
rect 116688 49745 116716 49943
rect 118606 49872 118662 49881
rect 118606 49807 118662 49816
rect 116674 49736 116730 49745
rect 116674 49671 116730 49680
rect 117962 49736 118018 49745
rect 117962 49671 118018 49680
rect 117976 40866 118004 49671
rect 118620 49162 118648 49807
rect 118608 49156 118660 49162
rect 118608 49098 118660 49104
rect 117964 40860 118016 40866
rect 117964 40802 118016 40808
rect 119356 16046 119384 50351
rect 122470 50280 122526 50289
rect 122470 50215 122526 50224
rect 120722 49872 120778 49881
rect 120722 49807 120778 49816
rect 120736 39438 120764 49807
rect 122102 49736 122158 49745
rect 122102 49671 122158 49680
rect 120724 39432 120776 39438
rect 120724 39374 120776 39380
rect 122116 38010 122144 49671
rect 122484 47666 122512 50215
rect 122472 47660 122524 47666
rect 122472 47602 122524 47608
rect 122104 38004 122156 38010
rect 122104 37946 122156 37952
rect 123496 17270 123524 50351
rect 126426 50280 126482 50289
rect 129278 50280 129334 50289
rect 126426 50215 126482 50224
rect 129200 50238 129278 50266
rect 125046 49872 125102 49881
rect 125046 49807 125102 49816
rect 124862 49736 124918 49745
rect 124862 49671 124918 49680
rect 124876 18698 124904 49671
rect 125060 20058 125088 49807
rect 126440 45554 126468 50215
rect 126518 50008 126574 50017
rect 126518 49943 126574 49952
rect 126532 49745 126560 49943
rect 127622 49872 127678 49881
rect 127622 49807 127678 49816
rect 126518 49736 126574 49745
rect 126518 49671 126574 49680
rect 126256 45526 126468 45554
rect 125048 20052 125100 20058
rect 125048 19994 125100 20000
rect 124864 18692 124916 18698
rect 124864 18634 124916 18640
rect 123484 17264 123536 17270
rect 123484 17206 123536 17212
rect 119344 16040 119396 16046
rect 119344 15982 119396 15988
rect 116584 14544 116636 14550
rect 116584 14486 116636 14492
rect 126256 11830 126284 45526
rect 126980 20052 127032 20058
rect 126980 19994 127032 20000
rect 126244 11824 126296 11830
rect 126244 11766 126296 11772
rect 115204 10396 115256 10402
rect 115204 10338 115256 10344
rect 125600 10396 125652 10402
rect 125600 10338 125652 10344
rect 122288 5364 122340 5370
rect 122288 5306 122340 5312
rect 119896 5228 119948 5234
rect 119896 5170 119948 5176
rect 116400 5160 116452 5166
rect 116400 5102 116452 5108
rect 115204 4888 115256 4894
rect 115204 4830 115256 4836
rect 115216 480 115244 4830
rect 116412 480 116440 5102
rect 118792 4956 118844 4962
rect 118792 4898 118844 4904
rect 117596 3392 117648 3398
rect 117596 3334 117648 3340
rect 117608 480 117636 3334
rect 118804 480 118832 4898
rect 119908 480 119936 5170
rect 121092 3324 121144 3330
rect 121092 3266 121144 3272
rect 121104 480 121132 3266
rect 122300 480 122328 5306
rect 123484 5296 123536 5302
rect 123484 5238 123536 5244
rect 123496 480 123524 5238
rect 124680 3256 124732 3262
rect 124680 3198 124732 3204
rect 124692 480 124720 3198
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125612 354 125640 10338
rect 126992 480 127020 19994
rect 127532 13116 127584 13122
rect 127532 13058 127584 13064
rect 127544 3482 127572 13058
rect 127636 4826 127664 49807
rect 129002 49736 129058 49745
rect 129002 49671 129058 49680
rect 128360 21412 128412 21418
rect 128360 21354 128412 21360
rect 128372 16574 128400 21354
rect 128372 16546 128952 16574
rect 127624 4820 127676 4826
rect 127624 4762 127676 4768
rect 127544 3454 128216 3482
rect 128188 480 128216 3454
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 129016 4894 129044 49671
rect 129200 4962 129228 50238
rect 129278 50215 129334 50224
rect 130382 49600 130438 49609
rect 130382 49535 130438 49544
rect 129740 43580 129792 43586
rect 129740 43522 129792 43528
rect 129752 16574 129780 43522
rect 129752 16546 130332 16574
rect 129188 4956 129240 4962
rect 129188 4898 129240 4904
rect 129004 4888 129056 4894
rect 129004 4830 129056 4836
rect 130304 3482 130332 16546
rect 130396 5370 130424 49535
rect 131776 28354 131804 50351
rect 131946 49736 132002 49745
rect 131946 49671 132002 49680
rect 131960 29646 131988 49671
rect 131948 29640 132000 29646
rect 131948 29582 132000 29588
rect 131764 28348 131816 28354
rect 131764 28290 131816 28296
rect 131120 28280 131172 28286
rect 131120 28222 131172 28228
rect 131132 16574 131160 28222
rect 132500 22908 132552 22914
rect 132500 22850 132552 22856
rect 132512 16574 132540 22850
rect 133156 19990 133184 50487
rect 138662 50416 138718 50425
rect 138662 50351 138718 50360
rect 141606 50416 141662 50425
rect 141606 50351 141662 50360
rect 136086 50280 136142 50289
rect 136086 50215 136142 50224
rect 134706 49872 134762 49881
rect 134706 49807 134762 49816
rect 134522 49736 134578 49745
rect 134522 49671 134578 49680
rect 134536 37942 134564 49671
rect 134720 39370 134748 49807
rect 136100 45554 136128 50215
rect 136178 50008 136234 50017
rect 136178 49943 136234 49952
rect 136192 49745 136220 49943
rect 137282 49872 137338 49881
rect 137282 49807 137338 49816
rect 136178 49736 136234 49745
rect 136178 49671 136234 49680
rect 135916 45526 136128 45554
rect 135916 40730 135944 45526
rect 135904 40724 135956 40730
rect 135904 40666 135956 40672
rect 134708 39364 134760 39370
rect 134708 39306 134760 39312
rect 134524 37936 134576 37942
rect 134524 37878 134576 37884
rect 133880 33924 133932 33930
rect 133880 33866 133932 33872
rect 133144 19984 133196 19990
rect 133144 19926 133196 19932
rect 131132 16546 131344 16574
rect 132512 16546 133000 16574
rect 130384 5364 130436 5370
rect 130384 5306 130436 5312
rect 130304 3454 130608 3482
rect 130580 480 130608 3454
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 132972 480 133000 16546
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 133892 354 133920 33866
rect 135260 32428 135312 32434
rect 135260 32370 135312 32376
rect 135272 480 135300 32370
rect 135352 24200 135404 24206
rect 135352 24142 135404 24148
rect 135364 16574 135392 24142
rect 135364 16546 136496 16574
rect 136468 480 136496 16546
rect 137192 11824 137244 11830
rect 137192 11766 137244 11772
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 11766
rect 137296 10334 137324 49807
rect 138020 47592 138072 47598
rect 138020 47534 138072 47540
rect 137284 10328 137336 10334
rect 137284 10270 137336 10276
rect 138032 6914 138060 47534
rect 138676 8022 138704 50351
rect 140042 50280 140098 50289
rect 140042 50215 140098 50224
rect 138846 49736 138902 49745
rect 138846 49671 138902 49680
rect 138860 42090 138888 49671
rect 138848 42084 138900 42090
rect 138848 42026 138900 42032
rect 140056 13190 140084 50215
rect 141422 49736 141478 49745
rect 141422 49671 141478 49680
rect 140780 25696 140832 25702
rect 140780 25638 140832 25644
rect 140792 16574 140820 25638
rect 140792 16546 141280 16574
rect 140044 13184 140096 13190
rect 140044 13126 140096 13132
rect 138664 8016 138716 8022
rect 138664 7958 138716 7964
rect 138032 6886 138888 6914
rect 138860 480 138888 6886
rect 140044 4820 140096 4826
rect 140044 4762 140096 4768
rect 140056 480 140084 4762
rect 141252 480 141280 16546
rect 141436 8090 141464 49671
rect 141620 26994 141648 50351
rect 141608 26988 141660 26994
rect 141608 26930 141660 26936
rect 142816 22778 142844 50487
rect 148506 50416 148562 50425
rect 148506 50351 148562 50360
rect 151082 50416 151138 50425
rect 151082 50351 151138 50360
rect 145838 50280 145894 50289
rect 145838 50215 145894 50224
rect 148322 50280 148378 50289
rect 148322 50215 148378 50224
rect 144182 49872 144238 49881
rect 144182 49807 144238 49816
rect 142804 22772 142856 22778
rect 142804 22714 142856 22720
rect 142160 17264 142212 17270
rect 142160 17206 142212 17212
rect 141424 8084 141476 8090
rect 141424 8026 141476 8032
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142172 354 142200 17206
rect 143540 13388 143592 13394
rect 143540 13330 143592 13336
rect 143552 3194 143580 13330
rect 144196 6254 144224 49807
rect 144366 49736 144422 49745
rect 144366 49671 144422 49680
rect 144380 17338 144408 49671
rect 145852 45554 145880 50215
rect 145930 50008 145986 50017
rect 145930 49943 145986 49952
rect 145944 49745 145972 49943
rect 145930 49736 145986 49745
rect 145930 49671 145986 49680
rect 146942 49736 146998 49745
rect 146942 49671 146998 49680
rect 145576 45526 145880 45554
rect 144368 17332 144420 17338
rect 144368 17274 144420 17280
rect 144920 17332 144972 17338
rect 144920 17274 144972 17280
rect 144932 16574 144960 17274
rect 144932 16546 145512 16574
rect 144184 6248 144236 6254
rect 144184 6190 144236 6196
rect 143632 4888 143684 4894
rect 143632 4830 143684 4836
rect 143540 3188 143592 3194
rect 143540 3130 143592 3136
rect 143644 2530 143672 4830
rect 144736 3188 144788 3194
rect 144736 3130 144788 3136
rect 143552 2502 143672 2530
rect 143552 480 143580 2502
rect 144748 480 144776 3130
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 145576 6322 145604 45526
rect 146956 6390 146984 49671
rect 147864 13456 147916 13462
rect 147864 13398 147916 13404
rect 146944 6384 146996 6390
rect 146944 6326 146996 6332
rect 145564 6316 145616 6322
rect 145564 6258 145616 6264
rect 147128 4956 147180 4962
rect 147128 4898 147180 4904
rect 147140 480 147168 4898
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 13398
rect 148336 6526 148364 50215
rect 148520 6594 148548 50351
rect 150530 49872 150586 49881
rect 150530 49807 150586 49816
rect 149794 49736 149850 49745
rect 149794 49671 149850 49680
rect 149808 45554 149836 49671
rect 150440 49224 150492 49230
rect 150440 49166 150492 49172
rect 149716 45526 149836 45554
rect 149716 36718 149744 45526
rect 149704 36712 149756 36718
rect 149704 36654 149756 36660
rect 149060 24132 149112 24138
rect 149060 24074 149112 24080
rect 149072 16574 149100 24074
rect 150452 16574 150480 49166
rect 150544 46238 150572 49807
rect 150532 46232 150584 46238
rect 150532 46174 150584 46180
rect 149072 16546 149560 16574
rect 150452 16546 150664 16574
rect 148508 6588 148560 6594
rect 148508 6530 148560 6536
rect 148324 6520 148376 6526
rect 148324 6462 148376 6468
rect 149532 480 149560 16546
rect 150636 480 150664 16546
rect 151096 14482 151124 50351
rect 151726 50280 151782 50289
rect 151726 50215 151782 50224
rect 151740 49745 151768 50215
rect 151726 49736 151782 49745
rect 151726 49671 151782 49680
rect 152476 35290 152504 50487
rect 155590 50416 155646 50425
rect 155328 50374 155590 50402
rect 153842 49872 153898 49881
rect 153842 49807 153898 49816
rect 152464 35284 152516 35290
rect 152464 35226 152516 35232
rect 153856 31142 153884 49807
rect 155328 45554 155356 50374
rect 155590 50351 155646 50360
rect 157798 50416 157854 50425
rect 157798 50351 157854 50360
rect 156602 50280 156658 50289
rect 156602 50215 156658 50224
rect 155406 49736 155462 49745
rect 155406 49671 155462 49680
rect 155236 45526 155356 45554
rect 154580 44940 154632 44946
rect 154580 44882 154632 44888
rect 153844 31136 153896 31142
rect 153844 31078 153896 31084
rect 153200 25628 153252 25634
rect 153200 25570 153252 25576
rect 151820 17400 151872 17406
rect 151820 17342 151872 17348
rect 151084 14476 151136 14482
rect 151084 14418 151136 14424
rect 151832 9674 151860 17342
rect 153212 16574 153240 25570
rect 154592 16574 154620 44882
rect 153212 16546 153792 16574
rect 154592 16546 155172 16574
rect 151912 13524 151964 13530
rect 151912 13466 151964 13472
rect 151740 9654 151860 9674
rect 151728 9648 151860 9654
rect 151780 9646 151860 9648
rect 151728 9590 151780 9596
rect 151924 6914 151952 13466
rect 153016 9648 153068 9654
rect 153016 9590 153068 9596
rect 151832 6886 151952 6914
rect 151832 480 151860 6886
rect 153028 480 153056 9590
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16546
rect 155144 3482 155172 16546
rect 155236 5030 155264 45526
rect 155420 44878 155448 49671
rect 155408 44872 155460 44878
rect 155408 44814 155460 44820
rect 155960 17468 156012 17474
rect 155960 17410 156012 17416
rect 155972 16574 156000 17410
rect 155972 16546 156184 16574
rect 155224 5024 155276 5030
rect 155224 4966 155276 4972
rect 155144 3454 155448 3482
rect 155420 480 155448 3454
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 156616 15978 156644 50215
rect 157812 50153 157840 50351
rect 159454 50280 159510 50289
rect 159454 50215 159510 50224
rect 157798 50144 157854 50153
rect 157798 50079 157854 50088
rect 158166 49872 158222 49881
rect 158166 49807 158222 49816
rect 157982 49736 158038 49745
rect 157982 49671 158038 49680
rect 156604 15972 156656 15978
rect 156604 15914 156656 15920
rect 157996 6662 158024 49671
rect 158180 18630 158208 49807
rect 159468 45554 159496 50215
rect 159546 50008 159602 50017
rect 159546 49943 159602 49952
rect 159560 49745 159588 49943
rect 159546 49736 159602 49745
rect 159546 49671 159602 49680
rect 159376 45526 159496 45554
rect 158720 22840 158772 22846
rect 158720 22782 158772 22788
rect 158168 18624 158220 18630
rect 158168 18566 158220 18572
rect 158732 16574 158760 22782
rect 158732 16546 158944 16574
rect 157984 6656 158036 6662
rect 157984 6598 158036 6604
rect 157800 6248 157852 6254
rect 157800 6190 157852 6196
rect 157812 480 157840 6190
rect 158916 480 158944 16546
rect 159376 5098 159404 45526
rect 160100 17536 160152 17542
rect 160100 17478 160152 17484
rect 159364 5092 159416 5098
rect 159364 5034 159416 5040
rect 160112 480 160140 17478
rect 160652 15972 160704 15978
rect 160652 15914 160704 15920
rect 160664 3482 160692 15914
rect 160756 5234 160784 50487
rect 160926 49736 160982 49745
rect 160926 49671 160982 49680
rect 160744 5228 160796 5234
rect 160744 5170 160796 5176
rect 160940 5166 160968 49671
rect 162136 5302 162164 50623
rect 170402 50552 170458 50561
rect 170402 50487 170458 50496
rect 165342 50416 165398 50425
rect 164896 50374 165342 50402
rect 163502 49872 163558 49881
rect 163502 49807 163558 49816
rect 162492 9036 162544 9042
rect 162492 8978 162544 8984
rect 162124 5296 162176 5302
rect 162124 5238 162176 5244
rect 160928 5160 160980 5166
rect 160928 5102 160980 5108
rect 160664 3454 161336 3482
rect 161308 480 161336 3454
rect 162504 480 162532 8978
rect 163516 7614 163544 49807
rect 164424 14612 164476 14618
rect 164424 14554 164476 14560
rect 163688 13184 163740 13190
rect 163688 13126 163740 13132
rect 163504 7608 163556 7614
rect 163504 7550 163556 7556
rect 163700 480 163728 13126
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164436 354 164464 14554
rect 164896 8974 164924 50374
rect 165342 50351 165398 50360
rect 167642 50416 167698 50425
rect 167826 50416 167882 50425
rect 167698 50374 167776 50402
rect 167642 50351 167698 50360
rect 166262 50280 166318 50289
rect 166262 50215 166318 50224
rect 167642 50280 167698 50289
rect 167642 50215 167698 50224
rect 165066 49736 165122 49745
rect 165066 49671 165122 49680
rect 165080 15910 165108 49671
rect 165068 15904 165120 15910
rect 165068 15846 165120 15852
rect 166276 9178 166304 50215
rect 167000 29640 167052 29646
rect 167000 29582 167052 29588
rect 167012 16574 167040 29582
rect 167012 16546 167224 16574
rect 166264 9172 166316 9178
rect 166264 9114 166316 9120
rect 166080 9104 166132 9110
rect 166080 9046 166132 9052
rect 164884 8968 164936 8974
rect 164884 8910 164936 8916
rect 166092 480 166120 9046
rect 167196 480 167224 16546
rect 167656 3806 167684 50215
rect 167748 50153 167776 50374
rect 167826 50351 167882 50360
rect 167734 50144 167790 50153
rect 167734 50079 167790 50088
rect 167840 3874 167868 50351
rect 169022 49872 169078 49881
rect 169022 49807 169078 49816
rect 168380 44872 168432 44878
rect 168380 44814 168432 44820
rect 167828 3868 167880 3874
rect 167828 3810 167880 3816
rect 167644 3800 167696 3806
rect 167644 3742 167696 3748
rect 168392 480 168420 44814
rect 169036 3942 169064 49807
rect 170312 13252 170364 13258
rect 170312 13194 170364 13200
rect 169576 9172 169628 9178
rect 169576 9114 169628 9120
rect 169024 3936 169076 3942
rect 169024 3878 169076 3884
rect 169588 480 169616 9114
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 13194
rect 170416 4010 170444 50487
rect 174726 50416 174782 50425
rect 174726 50351 174782 50360
rect 177118 50416 177174 50425
rect 177118 50351 177174 50360
rect 177486 50416 177542 50425
rect 177486 50351 177542 50360
rect 173162 50280 173218 50289
rect 173162 50215 173218 50224
rect 172150 49872 172206 49881
rect 172150 49807 172206 49816
rect 171782 49736 171838 49745
rect 171782 49671 171838 49680
rect 171692 10464 171744 10470
rect 171692 10406 171744 10412
rect 170404 4004 170456 4010
rect 170404 3946 170456 3952
rect 171704 3482 171732 10406
rect 171796 4078 171824 49671
rect 172164 45554 172192 49807
rect 171980 45526 172192 45554
rect 171980 16574 172008 45526
rect 172520 31204 172572 31210
rect 172520 31146 172572 31152
rect 172532 16574 172560 31146
rect 173176 29714 173204 50215
rect 173254 50008 173310 50017
rect 173254 49943 173310 49952
rect 173268 49745 173296 49943
rect 173254 49736 173310 49745
rect 173254 49671 173310 49680
rect 174542 49736 174598 49745
rect 174542 49671 174598 49680
rect 173164 29708 173216 29714
rect 173164 29650 173216 29656
rect 171980 16546 172100 16574
rect 172532 16546 172744 16574
rect 172072 4146 172100 16546
rect 172060 4140 172112 4146
rect 172060 4082 172112 4088
rect 171784 4072 171836 4078
rect 171784 4014 171836 4020
rect 171704 3454 172008 3482
rect 171980 480 172008 3454
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 173900 13320 173952 13326
rect 173900 13262 173952 13268
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173912 354 173940 13262
rect 174556 7682 174584 49671
rect 174740 33794 174768 50351
rect 176014 50280 176070 50289
rect 175936 50238 176014 50266
rect 175280 46232 175332 46238
rect 175280 46174 175332 46180
rect 174728 33788 174780 33794
rect 174728 33730 174780 33736
rect 175292 16574 175320 46174
rect 175292 16546 175504 16574
rect 174544 7676 174596 7682
rect 174544 7618 174596 7624
rect 175476 480 175504 16546
rect 175936 7750 175964 50238
rect 176014 50215 176070 50224
rect 177132 50153 177160 50351
rect 177118 50144 177174 50153
rect 177118 50079 177174 50088
rect 177302 49736 177358 49745
rect 177302 49671 177358 49680
rect 176660 36576 176712 36582
rect 176660 36518 176712 36524
rect 176672 11762 176700 36518
rect 176752 29776 176804 29782
rect 176752 29718 176804 29724
rect 176660 11756 176712 11762
rect 176660 11698 176712 11704
rect 175924 7744 175976 7750
rect 175924 7686 175976 7692
rect 176764 6914 176792 29718
rect 177316 7818 177344 49671
rect 177500 43450 177528 50351
rect 177488 43444 177540 43450
rect 177488 43386 177540 43392
rect 178040 18624 178092 18630
rect 178040 18566 178092 18572
rect 178052 16574 178080 18566
rect 178052 16546 178632 16574
rect 177856 11756 177908 11762
rect 177856 11698 177908 11704
rect 177304 7812 177356 7818
rect 177304 7754 177356 7760
rect 176672 6886 176792 6914
rect 176672 480 176700 6886
rect 177868 480 177896 11698
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 173134 -960 173246 326
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 178696 7886 178724 50623
rect 180062 50552 180118 50561
rect 180062 50487 180118 50496
rect 180076 26926 180104 50487
rect 180720 50425 180748 50623
rect 180706 50416 180762 50425
rect 180706 50351 180762 50360
rect 180800 35216 180852 35222
rect 180800 35158 180852 35164
rect 180064 26920 180116 26926
rect 180064 26862 180116 26868
rect 179420 21616 179472 21622
rect 179420 21558 179472 21564
rect 179432 16574 179460 21558
rect 180812 16574 180840 35158
rect 179432 16546 180288 16574
rect 180812 16546 181024 16574
rect 178684 7880 178736 7886
rect 178684 7822 178736 7828
rect 180260 480 180288 16546
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181456 7954 181484 50623
rect 181640 32502 181668 50759
rect 200762 50688 200818 50697
rect 200762 50623 200818 50632
rect 278686 50688 278742 50697
rect 278686 50623 278742 50632
rect 288346 50688 288402 50697
rect 288346 50623 288402 50632
rect 363050 50688 363106 50697
rect 363050 50623 363106 50632
rect 410522 50688 410578 50697
rect 410522 50623 410578 50632
rect 421746 50688 421802 50697
rect 421746 50623 421802 50632
rect 424506 50688 424562 50697
rect 424506 50623 424562 50632
rect 431314 50688 431370 50697
rect 431314 50623 431370 50632
rect 434626 50688 434682 50697
rect 434626 50623 434682 50632
rect 185582 50552 185638 50561
rect 185582 50487 185638 50496
rect 195242 50552 195298 50561
rect 195242 50487 195298 50496
rect 199382 50552 199438 50561
rect 199382 50487 199438 50496
rect 184846 50416 184902 50425
rect 184846 50351 184902 50360
rect 182822 49872 182878 49881
rect 182822 49807 182878 49816
rect 181628 32496 181680 32502
rect 181628 32438 181680 32444
rect 182836 8158 182864 49807
rect 184202 49736 184258 49745
rect 184202 49671 184258 49680
rect 183560 18828 183612 18834
rect 183560 18770 183612 18776
rect 183572 16574 183600 18770
rect 183572 16546 183784 16574
rect 182824 8152 182876 8158
rect 182824 8094 182876 8100
rect 181444 7948 181496 7954
rect 181444 7890 181496 7896
rect 182548 7608 182600 7614
rect 182548 7550 182600 7556
rect 182560 480 182588 7550
rect 183756 480 183784 16546
rect 184216 8226 184244 49671
rect 184860 49094 184888 50351
rect 184848 49088 184900 49094
rect 184848 49030 184900 49036
rect 184940 33788 184992 33794
rect 184940 33730 184992 33736
rect 184204 8220 184256 8226
rect 184204 8162 184256 8168
rect 184952 480 184980 33730
rect 185032 19984 185084 19990
rect 185032 19926 185084 19932
rect 185044 6914 185072 19926
rect 185596 9246 185624 50487
rect 188526 50416 188582 50425
rect 188526 50351 188582 50360
rect 190918 50416 190974 50425
rect 190918 50351 190974 50360
rect 193862 50416 193918 50425
rect 193862 50351 193918 50360
rect 186962 49736 187018 49745
rect 186962 49671 187018 49680
rect 186320 39568 186372 39574
rect 186320 39510 186372 39516
rect 186332 16574 186360 39510
rect 186976 36650 187004 49671
rect 188342 49600 188398 49609
rect 188342 49535 188398 49544
rect 186964 36644 187016 36650
rect 186964 36586 187016 36592
rect 187700 31068 187752 31074
rect 187700 31010 187752 31016
rect 187712 16574 187740 31010
rect 186332 16546 186912 16574
rect 187712 16546 188292 16574
rect 185584 9240 185636 9246
rect 185584 9182 185636 9188
rect 185044 6886 186176 6914
rect 186148 480 186176 6886
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 181414 -960 181526 326
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 188264 3482 188292 16546
rect 188356 6186 188384 49535
rect 188540 42158 188568 50351
rect 189722 50280 189778 50289
rect 189722 50215 189778 50224
rect 188528 42152 188580 42158
rect 188528 42094 188580 42100
rect 189736 6458 189764 50215
rect 190932 50153 190960 50351
rect 192574 50280 192630 50289
rect 192496 50238 192574 50266
rect 190918 50144 190974 50153
rect 190918 50079 190974 50088
rect 191102 49872 191158 49881
rect 191102 49807 191158 49816
rect 190460 47728 190512 47734
rect 190460 47670 190512 47676
rect 189724 6452 189776 6458
rect 189724 6394 189776 6400
rect 188344 6180 188396 6186
rect 188344 6122 188396 6128
rect 189724 5024 189776 5030
rect 189724 4966 189776 4972
rect 188264 3454 188568 3482
rect 188540 480 188568 3454
rect 189736 480 189764 4966
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190472 354 190500 47670
rect 191116 3398 191144 49807
rect 191286 49736 191342 49745
rect 191286 49671 191342 49680
rect 191300 40798 191328 49671
rect 191288 40792 191340 40798
rect 191288 40734 191340 40740
rect 191840 39364 191892 39370
rect 191840 39306 191892 39312
rect 191852 16574 191880 39306
rect 191852 16546 192064 16574
rect 191104 3392 191156 3398
rect 191104 3334 191156 3340
rect 192036 480 192064 16546
rect 192496 3330 192524 50238
rect 192574 50215 192630 50224
rect 192574 50008 192630 50017
rect 192574 49943 192630 49952
rect 192588 49745 192616 49943
rect 192574 49736 192630 49745
rect 192574 49671 192630 49680
rect 193220 38072 193272 38078
rect 193220 38014 193272 38020
rect 193232 3534 193260 38014
rect 193312 5092 193364 5098
rect 193312 5034 193364 5040
rect 193220 3528 193272 3534
rect 193220 3470 193272 3476
rect 192484 3324 192536 3330
rect 192484 3266 192536 3272
rect 193324 2530 193352 5034
rect 193876 3602 193904 50351
rect 194046 49736 194102 49745
rect 194046 49671 194102 49680
rect 193864 3596 193916 3602
rect 193864 3538 193916 3544
rect 194060 3262 194088 49671
rect 194600 42084 194652 42090
rect 194600 42026 194652 42032
rect 194612 16574 194640 42026
rect 194612 16546 195192 16574
rect 194416 3528 194468 3534
rect 194416 3470 194468 3476
rect 194048 3256 194100 3262
rect 194048 3198 194100 3204
rect 193232 2502 193352 2530
rect 193232 480 193260 2502
rect 194428 480 194456 3470
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 195256 3670 195284 50487
rect 198462 50416 198518 50425
rect 198016 50374 198462 50402
rect 196622 49736 196678 49745
rect 196622 49671 196678 49680
rect 196636 3738 196664 49671
rect 197360 49156 197412 49162
rect 197360 49098 197412 49104
rect 197372 16574 197400 49098
rect 197372 16546 197952 16574
rect 196808 5160 196860 5166
rect 196808 5102 196860 5108
rect 196624 3732 196676 3738
rect 196624 3674 196676 3680
rect 195244 3664 195296 3670
rect 195244 3606 195296 3612
rect 196820 480 196848 5102
rect 197924 480 197952 16546
rect 198016 3466 198044 50374
rect 198462 50351 198518 50360
rect 198186 49600 198242 49609
rect 198186 49535 198242 49544
rect 198200 3806 198228 49535
rect 198740 49020 198792 49026
rect 198740 48962 198792 48968
rect 198188 3800 198240 3806
rect 198188 3742 198240 3748
rect 198004 3460 198056 3466
rect 198004 3402 198056 3408
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 48962
rect 199396 3369 199424 50487
rect 200120 47660 200172 47666
rect 200120 47602 200172 47608
rect 200132 16574 200160 47602
rect 200132 16546 200344 16574
rect 199382 3360 199438 3369
rect 199382 3295 199438 3304
rect 200316 480 200344 16546
rect 200776 10402 200804 50623
rect 214562 50552 214618 50561
rect 214562 50487 214618 50496
rect 221462 50552 221518 50561
rect 221462 50487 221518 50496
rect 225602 50552 225658 50561
rect 225602 50487 225658 50496
rect 227718 50552 227774 50561
rect 227718 50487 227774 50496
rect 250994 50552 251050 50561
rect 250994 50487 251050 50496
rect 259366 50552 259422 50561
rect 259366 50487 259422 50496
rect 269026 50552 269082 50561
rect 269026 50487 269082 50496
rect 277306 50552 277362 50561
rect 277306 50487 277362 50496
rect 211802 50416 211858 50425
rect 211802 50351 211858 50360
rect 203522 50280 203578 50289
rect 203522 50215 203578 50224
rect 206282 50280 206338 50289
rect 206282 50215 206338 50224
rect 209134 50280 209190 50289
rect 209134 50215 209190 50224
rect 202142 49872 202198 49881
rect 202142 49807 202198 49816
rect 200946 49736 201002 49745
rect 200946 49671 201002 49680
rect 200960 21418 200988 49671
rect 201500 46368 201552 46374
rect 201500 46310 201552 46316
rect 200948 21412 201000 21418
rect 200948 21354 201000 21360
rect 200764 10396 200816 10402
rect 200764 10338 200816 10344
rect 201512 480 201540 46310
rect 201592 25560 201644 25566
rect 201592 25502 201644 25508
rect 201604 16574 201632 25502
rect 202156 22914 202184 49807
rect 203536 24206 203564 50215
rect 204258 50008 204314 50017
rect 204258 49943 204314 49952
rect 203890 49872 203946 49881
rect 204272 49858 204300 49943
rect 203946 49830 204300 49858
rect 204902 49872 204958 49881
rect 203890 49807 203946 49816
rect 204902 49807 204958 49816
rect 204260 42288 204312 42294
rect 204260 42230 204312 42236
rect 203524 24200 203576 24206
rect 203524 24142 203576 24148
rect 202144 22908 202196 22914
rect 202144 22850 202196 22856
rect 204272 16574 204300 42230
rect 201604 16546 202736 16574
rect 204272 16546 204852 16574
rect 202708 480 202736 16546
rect 203892 6180 203944 6186
rect 203892 6122 203944 6128
rect 203904 480 203932 6122
rect 204824 3482 204852 16546
rect 204916 4826 204944 49807
rect 205086 49736 205142 49745
rect 205086 49671 205142 49680
rect 205100 16574 205128 49671
rect 205100 16546 205220 16574
rect 205192 4894 205220 16546
rect 206192 14476 206244 14482
rect 206192 14418 206244 14424
rect 205180 4888 205232 4894
rect 205180 4830 205232 4836
rect 204904 4820 204956 4826
rect 204904 4762 204956 4768
rect 204824 3454 205128 3482
rect 205100 480 205128 3454
rect 206204 480 206232 14418
rect 206296 4962 206324 50215
rect 208122 49872 208178 49881
rect 208122 49807 208178 49816
rect 207662 49600 207718 49609
rect 207662 49535 207718 49544
rect 207676 25634 207704 49535
rect 208136 49230 208164 49807
rect 208124 49224 208176 49230
rect 208124 49166 208176 49172
rect 209148 45554 209176 50215
rect 211066 49872 211122 49881
rect 210528 49830 211066 49858
rect 210528 45554 210556 49830
rect 211066 49807 211122 49816
rect 210606 49736 210662 49745
rect 210606 49671 210662 49680
rect 209056 45526 209176 45554
rect 210436 45526 210556 45554
rect 207664 25628 207716 25634
rect 207664 25570 207716 25576
rect 208584 10328 208636 10334
rect 208584 10270 208636 10276
rect 206284 4956 206336 4962
rect 206284 4898 206336 4904
rect 207388 4820 207440 4826
rect 207388 4762 207440 4768
rect 207400 480 207428 4762
rect 208596 480 208624 10270
rect 209056 6254 209084 45526
rect 209780 15904 209832 15910
rect 209780 15846 209832 15852
rect 209792 9674 209820 15846
rect 210436 14618 210464 45526
rect 210620 15978 210648 49671
rect 211816 44878 211844 50351
rect 213182 49736 213238 49745
rect 213182 49671 213238 49680
rect 211804 44872 211856 44878
rect 211804 44814 211856 44820
rect 210608 15972 210660 15978
rect 210608 15914 210660 15920
rect 210424 14612 210476 14618
rect 210424 14554 210476 14560
rect 209872 14544 209924 14550
rect 209872 14486 209924 14492
rect 209700 9654 209820 9674
rect 209688 9648 209820 9654
rect 209740 9646 209820 9648
rect 209688 9590 209740 9596
rect 209884 6914 209912 14486
rect 213196 10470 213224 49671
rect 214576 18630 214604 50487
rect 218702 50416 218758 50425
rect 218702 50351 218758 50360
rect 214930 50280 214986 50289
rect 214930 50215 214986 50224
rect 214944 46238 214972 50215
rect 217322 49872 217378 49881
rect 217322 49807 217378 49816
rect 215942 49736 215998 49745
rect 215942 49671 215998 49680
rect 214932 46232 214984 46238
rect 214932 46174 214984 46180
rect 215300 40928 215352 40934
rect 215300 40870 215352 40876
rect 214564 18624 214616 18630
rect 214564 18566 214616 18572
rect 213368 14612 213420 14618
rect 213368 14554 213420 14560
rect 213184 10464 213236 10470
rect 213184 10406 213236 10412
rect 211712 10396 211764 10402
rect 211712 10338 211764 10344
rect 210976 9648 211028 9654
rect 210976 9590 211028 9596
rect 209792 6886 209912 6914
rect 209044 6248 209096 6254
rect 209044 6190 209096 6196
rect 209792 480 209820 6886
rect 210988 480 211016 9590
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 10338
rect 213380 480 213408 14554
rect 214472 4752 214524 4758
rect 214472 4694 214524 4700
rect 214484 480 214512 4694
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 40870
rect 215956 7614 215984 49671
rect 216864 14680 216916 14686
rect 216864 14622 216916 14628
rect 215944 7608 215996 7614
rect 215944 7550 215996 7556
rect 216876 480 216904 14622
rect 217336 5030 217364 49807
rect 217506 49600 217562 49609
rect 217506 49535 217562 49544
rect 217520 19990 217548 49535
rect 218060 20256 218112 20262
rect 218060 20198 218112 20204
rect 217508 19984 217560 19990
rect 217508 19926 217560 19932
rect 217324 5024 217376 5030
rect 217324 4966 217376 4972
rect 218072 3534 218100 20198
rect 218716 5098 218744 50351
rect 220082 49736 220138 49745
rect 220082 49671 220138 49680
rect 219440 43444 219492 43450
rect 219440 43386 219492 43392
rect 219452 16574 219480 43386
rect 219452 16546 220032 16574
rect 218704 5092 218756 5098
rect 218704 5034 218756 5040
rect 218152 4956 218204 4962
rect 218152 4898 218204 4904
rect 218060 3528 218112 3534
rect 218060 3470 218112 3476
rect 218164 2530 218192 4898
rect 219256 3528 219308 3534
rect 219256 3470 219308 3476
rect 218072 2502 218192 2530
rect 218072 480 218100 2502
rect 219268 480 219296 3470
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 220096 5166 220124 49671
rect 221476 6186 221504 50487
rect 221830 50280 221886 50289
rect 224682 50280 224738 50289
rect 221830 50215 221886 50224
rect 224328 50238 224682 50266
rect 221844 47666 221872 50215
rect 222842 49872 222898 49881
rect 222842 49807 222898 49816
rect 221832 47660 221884 47666
rect 221832 47602 221884 47608
rect 222752 10464 222804 10470
rect 222752 10406 222804 10412
rect 221464 6180 221516 6186
rect 221464 6122 221516 6128
rect 221556 5568 221608 5574
rect 221556 5510 221608 5516
rect 220084 5160 220136 5166
rect 220084 5102 220136 5108
rect 221568 480 221596 5510
rect 222764 480 222792 10406
rect 222856 4826 222884 49807
rect 224328 45554 224356 50238
rect 224682 50215 224738 50224
rect 224406 49736 224462 49745
rect 224406 49671 224462 49680
rect 224236 45526 224356 45554
rect 223580 18624 223632 18630
rect 223580 18566 223632 18572
rect 222844 4820 222896 4826
rect 222844 4762 222896 4768
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 220422 -960 220534 326
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223592 354 223620 18566
rect 224236 4758 224264 45526
rect 224420 15910 224448 49671
rect 224408 15904 224460 15910
rect 224408 15846 224460 15852
rect 225616 4962 225644 50487
rect 226982 49872 227038 49881
rect 226982 49807 227038 49816
rect 226340 14748 226392 14754
rect 226340 14690 226392 14696
rect 225604 4956 225656 4962
rect 225604 4898 225656 4904
rect 224224 4752 224276 4758
rect 224224 4694 224276 4700
rect 225144 4208 225196 4214
rect 225144 4150 225196 4156
rect 225156 480 225184 4150
rect 226352 3602 226380 14690
rect 226432 7744 226484 7750
rect 226432 7686 226484 7692
rect 226340 3596 226392 3602
rect 226340 3538 226392 3544
rect 226444 3482 226472 7686
rect 226996 4214 227024 49807
rect 227166 49736 227222 49745
rect 227166 49671 227222 49680
rect 227180 5574 227208 49671
rect 227732 16574 227760 50487
rect 233146 50416 233202 50425
rect 233146 50351 233202 50360
rect 234434 50416 234490 50425
rect 234434 50351 234490 50360
rect 249706 50416 249762 50425
rect 249706 50351 249762 50360
rect 231490 50280 231546 50289
rect 231490 50215 231546 50224
rect 230386 49872 230442 49881
rect 230386 49807 230442 49816
rect 227732 16546 228312 16574
rect 227168 5568 227220 5574
rect 227168 5510 227220 5516
rect 226984 4208 227036 4214
rect 226984 4150 227036 4156
rect 227536 3596 227588 3602
rect 227536 3538 227588 3544
rect 226352 3454 226472 3482
rect 226352 480 226380 3454
rect 227548 480 227576 3538
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16546
rect 229376 10532 229428 10538
rect 229376 10474 229428 10480
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 10474
rect 230400 4214 230428 49807
rect 231032 14816 231084 14822
rect 231032 14758 231084 14764
rect 230388 4208 230440 4214
rect 230388 4150 230440 4156
rect 231044 480 231072 14758
rect 231504 4826 231532 50215
rect 231674 49736 231730 49745
rect 231674 49671 231730 49680
rect 231492 4820 231544 4826
rect 231492 4762 231544 4768
rect 231688 4282 231716 49671
rect 233160 6254 233188 50351
rect 234448 45554 234476 50351
rect 235906 50280 235962 50289
rect 235906 50215 235962 50224
rect 238482 50280 238538 50289
rect 238482 50215 238538 50224
rect 241426 50280 241482 50289
rect 241426 50215 241482 50224
rect 248050 50280 248106 50289
rect 248050 50215 248106 50224
rect 234526 49872 234582 49881
rect 234526 49807 234582 49816
rect 234356 45526 234476 45554
rect 233240 18896 233292 18902
rect 233240 18838 233292 18844
rect 233252 16574 233280 18838
rect 233252 16546 233464 16574
rect 233148 6248 233200 6254
rect 233148 6190 233200 6196
rect 231676 4276 231728 4282
rect 231676 4218 231728 4224
rect 232228 4208 232280 4214
rect 232228 4150 232280 4156
rect 232240 480 232268 4150
rect 233436 480 233464 16546
rect 234356 7818 234384 45526
rect 234344 7812 234396 7818
rect 234344 7754 234396 7760
rect 234540 6186 234568 49807
rect 235920 15910 235948 50215
rect 237286 49736 237342 49745
rect 237286 49671 237342 49680
rect 236000 21684 236052 21690
rect 236000 21626 236052 21632
rect 236012 16574 236040 21626
rect 236012 16546 236592 16574
rect 235908 15904 235960 15910
rect 235908 15846 235960 15852
rect 234620 14884 234672 14890
rect 234620 14826 234672 14832
rect 234528 6180 234580 6186
rect 234528 6122 234580 6128
rect 234632 480 234660 14826
rect 235816 4276 235868 4282
rect 235816 4218 235868 4224
rect 235828 480 235856 4218
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 237300 7682 237328 49671
rect 238496 19990 238524 50215
rect 241242 49872 241298 49881
rect 241242 49807 241298 49816
rect 238666 49736 238722 49745
rect 238666 49671 238722 49680
rect 238484 19984 238536 19990
rect 238484 19926 238536 19932
rect 238680 18698 238708 49671
rect 240140 36848 240192 36854
rect 240140 36790 240192 36796
rect 238668 18692 238720 18698
rect 238668 18634 238720 18640
rect 237288 7676 237340 7682
rect 237288 7618 237340 7624
rect 239312 4820 239364 4826
rect 239312 4762 239364 4768
rect 238116 3460 238168 3466
rect 238116 3402 238168 3408
rect 238128 480 238156 3402
rect 239324 480 239352 4762
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 236982 -960 237094 326
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240152 354 240180 36790
rect 241256 21418 241284 49807
rect 241244 21412 241296 21418
rect 241244 21354 241296 21360
rect 241440 7614 241468 50215
rect 242714 50008 242770 50017
rect 242714 49943 242770 49952
rect 246762 50008 246818 50017
rect 246762 49943 246818 49952
rect 242728 47666 242756 49943
rect 242806 49736 242862 49745
rect 242806 49671 242862 49680
rect 245566 49736 245622 49745
rect 245566 49671 245622 49680
rect 242716 47660 242768 47666
rect 242716 47602 242768 47608
rect 241520 40724 241572 40730
rect 241520 40666 241572 40672
rect 241532 16574 241560 40666
rect 242820 22914 242848 49671
rect 244280 37936 244332 37942
rect 244280 37878 244332 37884
rect 242900 28484 242952 28490
rect 242900 28426 242952 28432
rect 242808 22908 242860 22914
rect 242808 22850 242860 22856
rect 242164 21480 242216 21486
rect 242164 21422 242216 21428
rect 241532 16546 241744 16574
rect 241428 7608 241480 7614
rect 241428 7550 241480 7556
rect 241716 480 241744 16546
rect 242176 3466 242204 21422
rect 242912 3534 242940 28426
rect 244292 16574 244320 37878
rect 244292 16546 245240 16574
rect 242992 6248 243044 6254
rect 242992 6190 243044 6196
rect 242900 3528 242952 3534
rect 242900 3470 242952 3476
rect 242164 3460 242216 3466
rect 242164 3402 242216 3408
rect 243004 3210 243032 6190
rect 244096 3528 244148 3534
rect 244096 3470 244148 3476
rect 242912 3182 243032 3210
rect 242912 480 242940 3182
rect 244108 480 244136 3470
rect 245212 480 245240 16546
rect 245580 4962 245608 49671
rect 246776 46306 246804 49943
rect 246946 49872 247002 49881
rect 246946 49807 247002 49816
rect 246854 49600 246910 49609
rect 246854 49535 246910 49544
rect 246764 46300 246816 46306
rect 246764 46242 246816 46248
rect 246868 45554 246896 49535
rect 246960 49094 246988 49807
rect 246948 49088 247000 49094
rect 246948 49030 247000 49036
rect 246868 45526 246988 45554
rect 246396 7812 246448 7818
rect 246396 7754 246448 7760
rect 245568 4956 245620 4962
rect 245568 4898 245620 4904
rect 246408 480 246436 7754
rect 246960 5166 246988 45526
rect 248064 39438 248092 50215
rect 248234 49736 248290 49745
rect 248234 49671 248290 49680
rect 248248 44878 248276 49671
rect 248236 44872 248288 44878
rect 248236 44814 248288 44820
rect 248052 39432 248104 39438
rect 248052 39374 248104 39380
rect 247040 32632 247092 32638
rect 247040 32574 247092 32580
rect 247052 16574 247080 32574
rect 247052 16546 247632 16574
rect 246948 5160 247000 5166
rect 246948 5102 247000 5108
rect 247604 480 247632 16546
rect 249720 5098 249748 50351
rect 250810 49872 250866 49881
rect 250810 49807 250866 49816
rect 249984 6180 250036 6186
rect 249984 6122 250036 6128
rect 249708 5092 249760 5098
rect 249708 5034 249760 5040
rect 248788 3596 248840 3602
rect 248788 3538 248840 3544
rect 248800 480 248828 3538
rect 249996 480 250024 6122
rect 250824 4894 250852 49807
rect 251008 5030 251036 50487
rect 253754 50416 253810 50425
rect 253754 50351 253810 50360
rect 253570 50280 253626 50289
rect 253570 50215 253626 50224
rect 252466 49736 252522 49745
rect 252466 49671 252522 49680
rect 251180 35488 251232 35494
rect 251180 35430 251232 35436
rect 250996 5024 251048 5030
rect 250996 4966 251048 4972
rect 250812 4888 250864 4894
rect 250812 4830 250864 4836
rect 251192 480 251220 35430
rect 252480 4758 252508 49671
rect 253204 46232 253256 46238
rect 253204 46174 253256 46180
rect 253112 15904 253164 15910
rect 253112 15846 253164 15852
rect 252468 4752 252520 4758
rect 252468 4694 252520 4700
rect 253124 3482 253152 15846
rect 253216 3602 253244 46174
rect 253584 38010 253612 50215
rect 253768 42158 253796 50351
rect 257894 50280 257950 50289
rect 257894 50215 257950 50224
rect 257802 49872 257858 49881
rect 256608 49836 256660 49842
rect 257802 49807 257804 49816
rect 256608 49778 256660 49784
rect 257856 49807 257858 49816
rect 257804 49778 257856 49784
rect 255226 49736 255282 49745
rect 255226 49671 255282 49680
rect 253756 42152 253808 42158
rect 253756 42094 253808 42100
rect 253572 38004 253624 38010
rect 253572 37946 253624 37952
rect 253940 31408 253992 31414
rect 253940 31350 253992 31356
rect 253952 16574 253980 31350
rect 253952 16546 254256 16574
rect 253204 3596 253256 3602
rect 253204 3538 253256 3544
rect 253124 3454 253520 3482
rect 252376 3324 252428 3330
rect 252376 3266 252428 3272
rect 252388 480 252416 3266
rect 253492 480 253520 3454
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 255240 6730 255268 49671
rect 255964 11756 256016 11762
rect 255964 11698 256016 11704
rect 255228 6724 255280 6730
rect 255228 6666 255280 6672
rect 255872 3528 255924 3534
rect 255872 3470 255924 3476
rect 255884 480 255912 3470
rect 255976 3330 256004 11698
rect 256620 6662 256648 49778
rect 257802 49736 257858 49745
rect 257802 49671 257858 49680
rect 257816 45554 257844 49671
rect 257724 45526 257844 45554
rect 257068 7676 257120 7682
rect 257068 7618 257120 7624
rect 256608 6656 256660 6662
rect 256608 6598 256660 6604
rect 255964 3324 256016 3330
rect 255964 3266 256016 3272
rect 257080 480 257108 7618
rect 257724 6594 257752 45526
rect 257712 6588 257764 6594
rect 257712 6530 257764 6536
rect 257908 6526 257936 50215
rect 258080 29980 258132 29986
rect 258080 29922 258132 29928
rect 258092 16574 258120 29922
rect 258092 16546 258304 16574
rect 257896 6520 257948 6526
rect 257896 6462 257948 6468
rect 258276 480 258304 16546
rect 259380 6458 259408 50487
rect 266266 50416 266322 50425
rect 266266 50351 266322 50360
rect 262126 50280 262182 50289
rect 262126 50215 262182 50224
rect 264794 50280 264850 50289
rect 264794 50215 264850 50224
rect 260654 49872 260710 49881
rect 260654 49807 260710 49816
rect 260470 49736 260526 49745
rect 260470 49671 260526 49680
rect 259460 18692 259512 18698
rect 259460 18634 259512 18640
rect 259368 6452 259420 6458
rect 259368 6394 259420 6400
rect 259472 3534 259500 18634
rect 260484 6390 260512 49671
rect 260472 6384 260524 6390
rect 260472 6326 260524 6332
rect 260668 6322 260696 49807
rect 262140 43722 262168 50215
rect 262678 50008 262734 50017
rect 262678 49943 262734 49952
rect 262310 49872 262366 49881
rect 262692 49858 262720 49943
rect 262366 49830 262720 49858
rect 263506 49872 263562 49881
rect 262310 49807 262366 49816
rect 263506 49807 263562 49816
rect 262128 43716 262180 43722
rect 262128 43658 262180 43664
rect 260840 27192 260892 27198
rect 260840 27134 260892 27140
rect 260852 16574 260880 27134
rect 262864 22772 262916 22778
rect 262864 22714 262916 22720
rect 260852 16546 261800 16574
rect 260656 6316 260708 6322
rect 260656 6258 260708 6264
rect 259460 3528 259512 3534
rect 259460 3470 259512 3476
rect 260656 3528 260708 3534
rect 260656 3470 260708 3476
rect 259460 3392 259512 3398
rect 259460 3334 259512 3340
rect 259472 480 259500 3334
rect 260668 480 260696 3470
rect 261772 480 261800 16546
rect 262876 3602 262904 22714
rect 263520 6254 263548 49807
rect 264610 49736 264666 49745
rect 264610 49671 264666 49680
rect 263600 19984 263652 19990
rect 263600 19926 263652 19932
rect 263612 16574 263640 19926
rect 263612 16546 264192 16574
rect 263508 6248 263560 6254
rect 263508 6190 263560 6196
rect 262864 3596 262916 3602
rect 262864 3538 262916 3544
rect 262956 3460 263008 3466
rect 262956 3402 263008 3408
rect 262968 480 262996 3402
rect 264164 480 264192 16546
rect 264624 6186 264652 49671
rect 264808 41002 264836 50215
rect 264796 40996 264848 41002
rect 264796 40938 264848 40944
rect 266280 36922 266308 50351
rect 267554 49872 267610 49881
rect 267554 49807 267610 49816
rect 267370 49736 267426 49745
rect 267370 49671 267426 49680
rect 266268 36916 266320 36922
rect 266268 36858 266320 36864
rect 266360 26920 266412 26926
rect 266360 26862 266412 26868
rect 264980 24404 265032 24410
rect 264980 24346 265032 24352
rect 264612 6180 264664 6186
rect 264612 6122 264664 6128
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 264992 354 265020 24346
rect 266372 16574 266400 26862
rect 267384 24478 267412 49671
rect 267568 35562 267596 49807
rect 267740 47660 267792 47666
rect 267740 47602 267792 47608
rect 267556 35556 267608 35562
rect 267556 35498 267608 35504
rect 267372 24472 267424 24478
rect 267372 24414 267424 24420
rect 267004 24200 267056 24206
rect 267004 24142 267056 24148
rect 266372 16546 266584 16574
rect 266556 480 266584 16546
rect 267016 3398 267044 24142
rect 267004 3392 267056 3398
rect 267004 3334 267056 3340
rect 267752 480 267780 47602
rect 269040 25838 269068 50487
rect 271786 50280 271842 50289
rect 271786 50215 271842 50224
rect 274362 50280 274418 50289
rect 274362 50215 274418 50224
rect 270406 49872 270462 49881
rect 270406 49807 270462 49816
rect 270222 49736 270278 49745
rect 270222 49671 270278 49680
rect 270236 32706 270264 49671
rect 270224 32700 270276 32706
rect 270224 32642 270276 32648
rect 270420 27130 270448 49807
rect 270408 27124 270460 27130
rect 270408 27066 270460 27072
rect 269028 25832 269080 25838
rect 269028 25774 269080 25780
rect 271800 23050 271828 50215
rect 272430 50008 272486 50017
rect 272430 49943 272486 49952
rect 272062 49872 272118 49881
rect 272444 49858 272472 49943
rect 272118 49830 272472 49858
rect 273166 49872 273222 49881
rect 272062 49807 272118 49816
rect 273166 49807 273222 49816
rect 273180 34066 273208 49807
rect 273168 34060 273220 34066
rect 273168 34002 273220 34008
rect 274376 29918 274404 50215
rect 274546 49736 274602 49745
rect 274546 49671 274602 49680
rect 277214 49736 277270 49745
rect 277214 49671 277270 49680
rect 274364 29912 274416 29918
rect 274364 29854 274416 29860
rect 274560 28558 274588 49671
rect 275926 49600 275982 49609
rect 275926 49535 275982 49544
rect 275940 31346 275968 49535
rect 276020 47864 276072 47870
rect 276020 47806 276072 47812
rect 275928 31340 275980 31346
rect 275928 31282 275980 31288
rect 274548 28552 274600 28558
rect 274548 28494 274600 28500
rect 271788 23044 271840 23050
rect 271788 22986 271840 22992
rect 270500 21412 270552 21418
rect 270500 21354 270552 21360
rect 270512 16574 270540 21354
rect 271880 20324 271932 20330
rect 271880 20266 271932 20272
rect 271892 16574 271920 20266
rect 270512 16546 270816 16574
rect 271892 16546 272472 16574
rect 270040 15904 270092 15910
rect 270040 15846 270092 15852
rect 268384 11892 268436 11898
rect 268384 11834 268436 11840
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 11834
rect 270052 480 270080 15846
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 270788 354 270816 16546
rect 272444 480 272472 16546
rect 273260 15972 273312 15978
rect 273260 15914 273312 15920
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273272 354 273300 15914
rect 274824 7608 274876 7614
rect 274824 7550 274876 7556
rect 274836 480 274864 7550
rect 276032 480 276060 47806
rect 277228 45554 277256 49671
rect 277320 46442 277348 50487
rect 277308 46436 277360 46442
rect 277308 46378 277360 46384
rect 277228 45526 277348 45554
rect 277320 39642 277348 45526
rect 278700 45150 278728 50623
rect 286690 50552 286746 50561
rect 286690 50487 286746 50496
rect 281170 50416 281226 50425
rect 281170 50351 281226 50360
rect 285586 50416 285642 50425
rect 285586 50351 285642 50360
rect 278688 45144 278740 45150
rect 278688 45086 278740 45092
rect 277308 39636 277360 39642
rect 277308 39578 277360 39584
rect 277400 22908 277452 22914
rect 277400 22850 277452 22856
rect 277412 16574 277440 22850
rect 277412 16546 278360 16574
rect 276664 16040 276716 16046
rect 276664 15982 276716 15988
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276676 354 276704 15982
rect 278332 480 278360 16546
rect 280712 16108 280764 16114
rect 280712 16050 280764 16056
rect 279056 11960 279108 11966
rect 279056 11902 279108 11908
rect 277094 354 277206 480
rect 276676 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 11902
rect 280724 480 280752 16050
rect 281184 7682 281212 50351
rect 282734 49872 282790 49881
rect 283102 49872 283158 49881
rect 282734 49807 282790 49816
rect 282840 49830 283102 49858
rect 281354 49736 281410 49745
rect 281354 49671 281410 49680
rect 281368 38146 281396 49671
rect 282748 49230 282776 49807
rect 282736 49224 282788 49230
rect 282736 49166 282788 49172
rect 281540 49088 281592 49094
rect 281540 49030 281592 49036
rect 281356 38140 281408 38146
rect 281356 38082 281408 38088
rect 281172 7676 281224 7682
rect 281172 7618 281224 7624
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281552 354 281580 49030
rect 282840 7614 282868 49830
rect 283102 49807 283158 49816
rect 284022 49736 284078 49745
rect 284022 49671 284078 49680
rect 282920 46504 282972 46510
rect 282920 46446 282972 46452
rect 282932 16574 282960 46446
rect 284036 42362 284064 49671
rect 284300 46300 284352 46306
rect 284300 46242 284352 46248
rect 284024 42356 284076 42362
rect 284024 42298 284076 42304
rect 282932 16546 283144 16574
rect 282828 7608 282880 7614
rect 282828 7550 282880 7556
rect 283116 480 283144 16546
rect 284312 3602 284340 46242
rect 285600 24342 285628 50351
rect 286322 49872 286378 49881
rect 286322 49807 286378 49816
rect 286336 47802 286364 49807
rect 286324 47796 286376 47802
rect 286324 47738 286376 47744
rect 286704 25770 286732 50487
rect 286966 49872 287022 49881
rect 286966 49807 287022 49816
rect 286980 45554 287008 49807
rect 286888 45526 287008 45554
rect 286888 43654 286916 45526
rect 286876 43648 286928 43654
rect 286876 43590 286928 43596
rect 286692 25764 286744 25770
rect 286692 25706 286744 25712
rect 285588 24336 285640 24342
rect 285588 24278 285640 24284
rect 288360 22982 288388 50623
rect 292486 50552 292542 50561
rect 292486 50487 292542 50496
rect 315946 50552 316002 50561
rect 315946 50487 316002 50496
rect 330482 50552 330538 50561
rect 330482 50487 330538 50496
rect 336002 50552 336058 50561
rect 336002 50487 336058 50496
rect 343638 50552 343694 50561
rect 343638 50487 343694 50496
rect 354678 50552 354734 50561
rect 354678 50487 354734 50496
rect 290922 50416 290978 50425
rect 290844 50374 290922 50402
rect 289726 49736 289782 49745
rect 289726 49671 289782 49680
rect 289740 40866 289768 49671
rect 289728 40860 289780 40866
rect 289728 40802 289780 40808
rect 290844 35358 290872 50374
rect 290922 50351 290978 50360
rect 291014 49736 291070 49745
rect 291014 49671 291070 49680
rect 291028 36718 291056 49671
rect 291016 36712 291068 36718
rect 291016 36654 291068 36660
rect 290832 35352 290884 35358
rect 290832 35294 290884 35300
rect 292500 32570 292528 50487
rect 297730 50416 297786 50425
rect 297730 50351 297786 50360
rect 304814 50416 304870 50425
rect 304814 50351 304870 50360
rect 307482 50416 307538 50425
rect 307482 50351 307538 50360
rect 314290 50416 314346 50425
rect 314290 50351 314346 50360
rect 295246 50280 295302 50289
rect 295246 50215 295302 50224
rect 293590 49872 293646 49881
rect 293590 49807 293646 49816
rect 292580 39704 292632 39710
rect 292580 39646 292632 39652
rect 292488 32564 292540 32570
rect 292488 32506 292540 32512
rect 288348 22976 288400 22982
rect 288348 22918 288400 22924
rect 292592 16574 292620 39646
rect 293604 27062 293632 49807
rect 293774 49736 293830 49745
rect 293774 49671 293830 49680
rect 293788 33998 293816 49671
rect 293776 33992 293828 33998
rect 293776 33934 293828 33940
rect 293592 27056 293644 27062
rect 293592 26998 293644 27004
rect 292592 16546 293264 16574
rect 291384 16312 291436 16318
rect 291384 16254 291436 16260
rect 287336 16244 287388 16250
rect 287336 16186 287388 16192
rect 284392 16176 284444 16182
rect 284392 16118 284444 16124
rect 284300 3596 284352 3602
rect 284300 3538 284352 3544
rect 284404 3482 284432 16118
rect 286600 12028 286652 12034
rect 286600 11970 286652 11976
rect 285036 3596 285088 3602
rect 285036 3538 285088 3544
rect 284312 3454 284432 3482
rect 284312 480 284340 3454
rect 281878 354 281990 480
rect 281552 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285048 354 285076 3538
rect 286612 480 286640 11970
rect 285374 354 285486 480
rect 285048 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287348 354 287376 16186
rect 288992 4956 289044 4962
rect 288992 4898 289044 4904
rect 290188 4956 290240 4962
rect 290188 4898 290240 4904
rect 289004 480 289032 4898
rect 290200 480 290228 4898
rect 291396 480 291424 16254
rect 292580 5160 292632 5166
rect 292580 5102 292632 5108
rect 292592 480 292620 5102
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 294880 16380 294932 16386
rect 294880 16322 294932 16328
rect 294892 480 294920 16322
rect 295260 8974 295288 50215
rect 296626 49600 296682 49609
rect 296626 49535 296682 49544
rect 295340 44872 295392 44878
rect 295340 44814 295392 44820
rect 295352 16574 295380 44814
rect 296640 28422 296668 49535
rect 296628 28416 296680 28422
rect 296628 28358 296680 28364
rect 297744 18766 297772 50351
rect 297914 50280 297970 50289
rect 297914 50215 297970 50224
rect 300674 50280 300730 50289
rect 303526 50280 303582 50289
rect 300674 50215 300730 50224
rect 303448 50238 303526 50266
rect 297928 45014 297956 50215
rect 299386 49872 299442 49881
rect 299386 49807 299442 49816
rect 297916 45008 297968 45014
rect 297916 44950 297968 44956
rect 299400 20194 299428 49807
rect 300490 49736 300546 49745
rect 300490 49671 300546 49680
rect 299480 49292 299532 49298
rect 299480 49234 299532 49240
rect 299388 20188 299440 20194
rect 299388 20130 299440 20136
rect 297732 18760 297784 18766
rect 297732 18702 297784 18708
rect 295352 16546 295656 16574
rect 295248 8968 295300 8974
rect 295248 8910 295300 8916
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 295628 354 295656 16546
rect 298100 16448 298152 16454
rect 298100 16390 298152 16396
rect 297272 9240 297324 9246
rect 297272 9182 297324 9188
rect 297284 480 297312 9182
rect 296046 354 296158 480
rect 295628 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298112 354 298140 16390
rect 299492 3534 299520 49234
rect 299572 39432 299624 39438
rect 299572 39374 299624 39380
rect 299584 16574 299612 39374
rect 300504 21554 300532 49671
rect 300688 22914 300716 50215
rect 303448 45554 303476 50238
rect 303526 50215 303582 50224
rect 303526 49736 303582 49745
rect 303526 49671 303582 49680
rect 303356 45526 303476 45554
rect 303356 25634 303384 45526
rect 303344 25628 303396 25634
rect 303344 25570 303396 25576
rect 303540 24274 303568 49671
rect 304828 45554 304856 50351
rect 304906 49872 304962 49881
rect 304906 49807 304962 49816
rect 304920 47666 304948 49807
rect 306286 49736 306342 49745
rect 306286 49671 306342 49680
rect 304908 47660 304960 47666
rect 304908 47602 304960 47608
rect 304828 45526 304948 45554
rect 303620 38208 303672 38214
rect 303620 38150 303672 38156
rect 303528 24268 303580 24274
rect 303528 24210 303580 24216
rect 300676 22908 300728 22914
rect 300676 22850 300728 22856
rect 300492 21548 300544 21554
rect 300492 21490 300544 21496
rect 302884 20120 302936 20126
rect 302884 20062 302936 20068
rect 299584 16546 299704 16574
rect 299480 3528 299532 3534
rect 299480 3470 299532 3476
rect 299676 480 299704 16546
rect 300768 3528 300820 3534
rect 300768 3470 300820 3476
rect 301964 3528 302016 3534
rect 301964 3470 302016 3476
rect 300780 480 300808 3470
rect 301976 480 302004 3470
rect 302896 3466 302924 20062
rect 303632 16574 303660 38150
rect 304920 26994 304948 45526
rect 306300 28354 306328 49671
rect 307496 31142 307524 50351
rect 307666 50280 307722 50289
rect 307666 50215 307722 50224
rect 310426 50280 310482 50289
rect 310426 50215 310482 50224
rect 311806 50280 311862 50289
rect 311806 50215 311862 50224
rect 307484 31136 307536 31142
rect 307484 31078 307536 31084
rect 307680 29714 307708 50215
rect 310242 49872 310298 49881
rect 310242 49807 310298 49816
rect 307760 42424 307812 42430
rect 307760 42366 307812 42372
rect 307668 29708 307720 29714
rect 307668 29650 307720 29656
rect 306288 28348 306340 28354
rect 306288 28290 306340 28296
rect 304908 26988 304960 26994
rect 304908 26930 304960 26936
rect 305000 17604 305052 17610
rect 305000 17546 305052 17552
rect 305012 16574 305040 17546
rect 307772 16574 307800 42366
rect 310256 33862 310284 49807
rect 310244 33856 310296 33862
rect 310244 33798 310296 33804
rect 310440 32502 310468 50215
rect 311714 50008 311770 50017
rect 311714 49943 311770 49952
rect 311728 49094 311756 49943
rect 311716 49088 311768 49094
rect 311716 49030 311768 49036
rect 310520 43784 310572 43790
rect 310520 43726 310572 43732
rect 310428 32496 310480 32502
rect 310428 32438 310480 32444
rect 310532 16574 310560 43726
rect 311820 35290 311848 50215
rect 313186 49736 313242 49745
rect 313186 49671 313242 49680
rect 313200 36650 313228 49671
rect 313188 36644 313240 36650
rect 313188 36586 313240 36592
rect 311808 35284 311860 35290
rect 311808 35226 311860 35232
rect 303632 16546 303936 16574
rect 305012 16546 305592 16574
rect 307772 16546 307984 16574
rect 310532 16546 311480 16574
rect 303160 5092 303212 5098
rect 303160 5034 303212 5040
rect 302884 3460 302936 3466
rect 302884 3402 302936 3408
rect 303172 480 303200 5034
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305564 480 305592 16546
rect 306748 5024 306800 5030
rect 306748 4966 306800 4972
rect 306760 480 306788 4966
rect 307956 480 307984 16546
rect 310244 4888 310296 4894
rect 310244 4830 310296 4836
rect 309048 3596 309100 3602
rect 309048 3538 309100 3544
rect 309060 480 309088 3538
rect 310256 480 310284 4830
rect 311452 480 311480 16546
rect 313832 4820 313884 4826
rect 313832 4762 313884 4768
rect 312636 3460 312688 3466
rect 312636 3402 312688 3408
rect 312648 480 312676 3402
rect 313844 480 313872 4762
rect 314304 4758 314332 50351
rect 314474 49600 314530 49609
rect 314474 49535 314530 49544
rect 314488 4826 314516 49535
rect 315960 46306 315988 50487
rect 324134 50416 324190 50425
rect 324134 50351 324190 50360
rect 326158 50416 326214 50425
rect 326158 50351 326214 50360
rect 327722 50416 327778 50425
rect 327722 50351 327778 50360
rect 318706 50280 318762 50289
rect 318706 50215 318762 50224
rect 321466 50280 321522 50289
rect 321466 50215 321522 50224
rect 318154 50008 318210 50017
rect 318154 49943 318210 49952
rect 317142 49872 317198 49881
rect 317142 49807 317198 49816
rect 315948 46300 316000 46306
rect 315948 46242 316000 46248
rect 317156 39438 317184 49807
rect 318168 49745 318196 49943
rect 317326 49736 317382 49745
rect 317326 49671 317382 49680
rect 318154 49736 318210 49745
rect 318154 49671 318210 49680
rect 317144 39432 317196 39438
rect 317144 39374 317196 39380
rect 317340 38010 317368 49671
rect 318720 40798 318748 50215
rect 321098 50008 321154 50017
rect 321098 49943 321154 49952
rect 320086 49872 320142 49881
rect 319916 49830 320086 49858
rect 319916 45554 319944 49830
rect 320086 49807 320142 49816
rect 321112 49745 321140 49943
rect 319994 49736 320050 49745
rect 319994 49671 320050 49680
rect 321098 49736 321154 49745
rect 321098 49671 321154 49680
rect 319824 45526 319944 45554
rect 319824 43518 319852 45526
rect 320008 44878 320036 49671
rect 319996 44872 320048 44878
rect 319996 44814 320048 44820
rect 319812 43512 319864 43518
rect 319812 43454 319864 43460
rect 321480 42158 321508 50215
rect 322846 49736 322902 49745
rect 322846 49671 322902 49680
rect 321560 45212 321612 45218
rect 321560 45154 321612 45160
rect 320180 42152 320232 42158
rect 320180 42094 320232 42100
rect 321468 42152 321520 42158
rect 321468 42094 321520 42100
rect 318708 40792 318760 40798
rect 318708 40734 318760 40740
rect 316040 38004 316092 38010
rect 316040 37946 316092 37952
rect 317328 38004 317380 38010
rect 317328 37946 317380 37952
rect 315028 5024 315080 5030
rect 315028 4966 315080 4972
rect 314476 4820 314528 4826
rect 314476 4762 314528 4768
rect 314292 4752 314344 4758
rect 314292 4694 314344 4700
rect 315040 480 315068 4966
rect 316052 3398 316080 37946
rect 316132 17672 316184 17678
rect 316132 17614 316184 17620
rect 316144 16574 316172 17614
rect 320192 16574 320220 42094
rect 321572 16574 321600 45154
rect 322860 18698 322888 49671
rect 323950 49600 324006 49609
rect 323950 49535 324006 49544
rect 323964 19990 323992 49535
rect 324148 21418 324176 50351
rect 324962 50280 325018 50289
rect 324962 50215 325018 50224
rect 324136 21412 324188 21418
rect 324136 21354 324188 21360
rect 324976 20058 325004 50215
rect 326172 50153 326200 50351
rect 326158 50144 326214 50153
rect 326158 50079 326214 50088
rect 326342 49872 326398 49881
rect 326342 49807 326398 49816
rect 326356 33930 326384 49807
rect 326526 49736 326582 49745
rect 326526 49671 326582 49680
rect 326540 43586 326568 49671
rect 326528 43580 326580 43586
rect 326528 43522 326580 43528
rect 326344 33924 326396 33930
rect 326344 33866 326396 33872
rect 324964 20052 325016 20058
rect 324964 19994 325016 20000
rect 323952 19984 324004 19990
rect 323952 19926 324004 19932
rect 322848 18692 322900 18698
rect 322848 18634 322900 18640
rect 322940 17740 322992 17746
rect 322940 17682 322992 17688
rect 316144 16546 316264 16574
rect 320192 16546 320496 16574
rect 321572 16546 322152 16574
rect 316040 3392 316092 3398
rect 316040 3334 316092 3340
rect 316236 480 316264 16546
rect 318064 10600 318116 10606
rect 318064 10542 318116 10548
rect 317328 3392 317380 3398
rect 317328 3334 317380 3340
rect 317340 480 317368 3334
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 10542
rect 319720 3664 319772 3670
rect 319720 3606 319772 3612
rect 319732 480 319760 3606
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 322124 480 322152 16546
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 322952 354 322980 17682
rect 327736 11830 327764 50351
rect 329194 49872 329250 49881
rect 329194 49807 329250 49816
rect 329104 45076 329156 45082
rect 329104 45018 329156 45024
rect 327724 11824 327776 11830
rect 327724 11766 327776 11772
rect 325608 6792 325660 6798
rect 325608 6734 325660 6740
rect 324412 6724 324464 6730
rect 324412 6666 324464 6672
rect 324424 480 324452 6666
rect 325620 480 325648 6734
rect 328000 6656 328052 6662
rect 328000 6598 328052 6604
rect 326804 3800 326856 3806
rect 326804 3742 326856 3748
rect 326816 480 326844 3742
rect 328012 480 328040 6598
rect 329116 3534 329144 45018
rect 329208 25702 329236 49807
rect 329196 25696 329248 25702
rect 329196 25638 329248 25644
rect 330496 13462 330524 50487
rect 333702 50416 333758 50425
rect 333256 50374 333702 50402
rect 331862 50280 331918 50289
rect 331862 50215 331918 50224
rect 330666 49736 330722 49745
rect 330666 49671 330722 49680
rect 330484 13456 330536 13462
rect 330484 13398 330536 13404
rect 330680 13394 330708 49671
rect 331876 13530 331904 50215
rect 331956 39500 332008 39506
rect 331956 39442 332008 39448
rect 331864 13524 331916 13530
rect 331864 13466 331916 13472
rect 330668 13388 330720 13394
rect 330668 13330 330720 13336
rect 329196 6656 329248 6662
rect 329196 6598 329248 6604
rect 329104 3528 329156 3534
rect 329104 3470 329156 3476
rect 329208 480 329236 6598
rect 331588 6588 331640 6594
rect 331588 6530 331640 6536
rect 330392 3732 330444 3738
rect 330392 3674 330444 3680
rect 330404 480 330432 3674
rect 331600 480 331628 6530
rect 331968 3602 331996 39442
rect 333256 22846 333284 50374
rect 333702 50351 333758 50360
rect 334714 50280 334770 50289
rect 334714 50215 334770 50224
rect 333426 49736 333482 49745
rect 333426 49671 333482 49680
rect 333440 44946 333468 49671
rect 334728 45554 334756 50215
rect 334636 45526 334756 45554
rect 333428 44940 333480 44946
rect 333428 44882 333480 44888
rect 333244 22840 333296 22846
rect 333244 22782 333296 22788
rect 334636 9042 334664 45526
rect 336016 9178 336044 50487
rect 336186 49736 336242 49745
rect 336186 49671 336242 49680
rect 342258 49736 342314 49745
rect 342258 49671 342314 49680
rect 336004 9172 336056 9178
rect 336004 9114 336056 9120
rect 336200 9110 336228 49671
rect 340144 31272 340196 31278
rect 340144 31214 340196 31220
rect 338764 29844 338816 29850
rect 338764 29786 338816 29792
rect 336188 9104 336240 9110
rect 336188 9046 336240 9052
rect 334624 9036 334676 9042
rect 334624 8978 334676 8984
rect 332692 6588 332744 6594
rect 332692 6530 332744 6536
rect 331956 3596 332008 3602
rect 331956 3538 332008 3544
rect 332704 480 332732 6530
rect 335084 6520 335136 6526
rect 335084 6462 335136 6468
rect 336280 6520 336332 6526
rect 336280 6462 336332 6468
rect 333888 3528 333940 3534
rect 333888 3470 333940 3476
rect 333900 480 333928 3470
rect 335096 480 335124 6462
rect 336292 480 336320 6462
rect 338672 6452 338724 6458
rect 338672 6394 338724 6400
rect 337476 3868 337528 3874
rect 337476 3810 337528 3816
rect 337488 480 337516 3810
rect 338684 480 338712 6394
rect 338776 3466 338804 29786
rect 339868 6452 339920 6458
rect 339868 6394 339920 6400
rect 338764 3460 338816 3466
rect 338764 3402 338816 3408
rect 339880 480 339908 6394
rect 340156 3670 340184 31214
rect 342272 31210 342300 49671
rect 342904 42220 342956 42226
rect 342904 42162 342956 42168
rect 342260 31204 342312 31210
rect 342260 31146 342312 31152
rect 340972 11824 341024 11830
rect 340972 11766 341024 11772
rect 340144 3664 340196 3670
rect 340144 3606 340196 3612
rect 340984 480 341012 11766
rect 342168 6384 342220 6390
rect 342168 6326 342220 6332
rect 342180 480 342208 6326
rect 342916 3806 342944 42162
rect 343652 29782 343680 50487
rect 345202 50416 345258 50425
rect 345202 50351 345258 50360
rect 345018 50008 345074 50017
rect 345018 49943 345074 49952
rect 345032 47734 345060 49943
rect 345110 49736 345166 49745
rect 345110 49671 345166 49680
rect 345020 47728 345072 47734
rect 345020 47670 345072 47676
rect 345124 45554 345152 49671
rect 345032 45526 345152 45554
rect 343640 29776 343692 29782
rect 343640 29718 343692 29724
rect 345032 18834 345060 45526
rect 345216 21622 345244 50351
rect 346490 50280 346546 50289
rect 346490 50215 346546 50224
rect 351918 50280 351974 50289
rect 351974 50238 352052 50266
rect 351918 50215 351974 50224
rect 346398 49872 346454 49881
rect 346398 49807 346454 49816
rect 346412 49162 346440 49807
rect 346400 49156 346452 49162
rect 346400 49098 346452 49104
rect 346400 47932 346452 47938
rect 346400 47874 346452 47880
rect 345204 21616 345256 21622
rect 345204 21558 345256 21564
rect 345020 18828 345072 18834
rect 345020 18770 345072 18776
rect 345664 18828 345716 18834
rect 345664 18770 345716 18776
rect 343364 6384 343416 6390
rect 343364 6326 343416 6332
rect 342904 3800 342956 3806
rect 342904 3742 342956 3748
rect 343376 480 343404 6326
rect 345676 3874 345704 18770
rect 346412 16574 346440 47874
rect 346504 39574 346532 50215
rect 351826 49872 351882 49881
rect 351826 49807 351828 49816
rect 351880 49807 351882 49816
rect 351828 49778 351880 49784
rect 347962 49736 348018 49745
rect 347962 49671 348018 49680
rect 348146 49736 348202 49745
rect 348146 49671 348202 49680
rect 346492 39568 346544 39574
rect 346492 39510 346544 39516
rect 347976 38078 348004 49671
rect 348160 46374 348188 49671
rect 348148 46368 348200 46374
rect 348148 46310 348200 46316
rect 349160 43716 349212 43722
rect 349160 43658 349212 43664
rect 348424 43580 348476 43586
rect 348424 43522 348476 43528
rect 347964 38072 348016 38078
rect 347964 38014 348016 38020
rect 346412 16546 346992 16574
rect 345756 6316 345808 6322
rect 345756 6258 345808 6264
rect 345664 3868 345716 3874
rect 345664 3810 345716 3816
rect 344560 3596 344612 3602
rect 344560 3538 344612 3544
rect 344572 480 344600 3538
rect 345768 480 345796 6258
rect 346964 480 346992 16546
rect 348056 4140 348108 4146
rect 348056 4082 348108 4088
rect 348068 480 348096 4082
rect 348436 3738 348464 43522
rect 348424 3732 348476 3738
rect 348424 3674 348476 3680
rect 349172 3346 349200 43658
rect 352024 42294 352052 50238
rect 353300 49836 353352 49842
rect 353300 49778 353352 49784
rect 352194 49736 352250 49745
rect 352194 49671 352250 49680
rect 352012 42288 352064 42294
rect 352012 42230 352064 42236
rect 349252 41064 349304 41070
rect 349252 41006 349304 41012
rect 349264 3534 349292 41006
rect 352208 10334 352236 49671
rect 353312 10402 353340 49778
rect 353944 36780 353996 36786
rect 353944 36722 353996 36728
rect 353300 10396 353352 10402
rect 353300 10338 353352 10344
rect 352196 10328 352248 10334
rect 352196 10270 352248 10276
rect 352840 6248 352892 6254
rect 352840 6190 352892 6196
rect 351644 3664 351696 3670
rect 351644 3606 351696 3612
rect 349252 3528 349304 3534
rect 349252 3470 349304 3476
rect 350448 3528 350500 3534
rect 350448 3470 350500 3476
rect 349172 3318 349292 3346
rect 349264 480 349292 3318
rect 350460 480 350488 3470
rect 351656 480 351684 3606
rect 352852 480 352880 6190
rect 353956 3466 353984 36722
rect 354692 20262 354720 50487
rect 356058 50416 356114 50425
rect 356058 50351 356114 50360
rect 354862 49872 354918 49881
rect 354862 49807 354918 49816
rect 354876 40934 354904 49807
rect 354864 40928 354916 40934
rect 354864 40870 354916 40876
rect 354680 20256 354732 20262
rect 354680 20198 354732 20204
rect 356072 10470 356100 50351
rect 357714 50280 357770 50289
rect 357714 50215 357770 50224
rect 360198 50280 360254 50289
rect 360198 50215 360254 50224
rect 357530 49736 357586 49745
rect 357530 49671 357586 49680
rect 356704 21616 356756 21622
rect 356704 21558 356756 21564
rect 356060 10464 356112 10470
rect 356060 10406 356112 10412
rect 354036 6248 354088 6254
rect 354036 6190 354088 6196
rect 353944 3460 353996 3466
rect 353944 3402 353996 3408
rect 354048 480 354076 6190
rect 356336 6180 356388 6186
rect 356336 6122 356388 6128
rect 355232 3460 355284 3466
rect 355232 3402 355284 3408
rect 355244 480 355272 3402
rect 356348 480 356376 6122
rect 356716 4146 356744 21558
rect 357544 10538 357572 49671
rect 357532 10532 357584 10538
rect 357532 10474 357584 10480
rect 357728 7750 357756 50215
rect 358910 49872 358966 49881
rect 358910 49807 358966 49816
rect 358820 40996 358872 41002
rect 358820 40938 358872 40944
rect 358832 16574 358860 40938
rect 358924 18902 358952 49807
rect 360212 21690 360240 50215
rect 360658 50008 360714 50017
rect 360658 49943 360714 49952
rect 360672 49745 360700 49943
rect 361578 49872 361634 49881
rect 361634 49830 361712 49858
rect 361578 49807 361634 49816
rect 360658 49736 360714 49745
rect 360658 49671 360714 49680
rect 361578 49736 361634 49745
rect 361578 49671 361634 49680
rect 360844 35420 360896 35426
rect 360844 35362 360896 35368
rect 360200 21684 360252 21690
rect 360200 21626 360252 21632
rect 358912 18896 358964 18902
rect 358912 18838 358964 18844
rect 358832 16546 359504 16574
rect 357716 7744 357768 7750
rect 357716 7686 357768 7692
rect 357532 6180 357584 6186
rect 357532 6122 357584 6128
rect 356704 4140 356756 4146
rect 356704 4082 356756 4088
rect 357544 480 357572 6122
rect 358728 3732 358780 3738
rect 358728 3674 358780 3680
rect 358740 480 358768 3674
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 16546
rect 360856 3602 360884 35362
rect 361592 28490 361620 49671
rect 361684 45554 361712 49830
rect 361684 45526 361804 45554
rect 361776 36854 361804 45526
rect 362960 36916 363012 36922
rect 362960 36858 363012 36864
rect 361764 36848 361816 36854
rect 361764 36790 361816 36796
rect 361580 28484 361632 28490
rect 361580 28426 361632 28432
rect 362972 16574 363000 36858
rect 363064 32638 363092 50623
rect 364614 50552 364670 50561
rect 364614 50487 364670 50496
rect 382278 50552 382334 50561
rect 382278 50487 382334 50496
rect 398930 50552 398986 50561
rect 398930 50487 398986 50496
rect 364430 49872 364486 49881
rect 364430 49807 364486 49816
rect 364444 35494 364472 49807
rect 364432 35488 364484 35494
rect 364432 35430 364484 35436
rect 363052 32632 363104 32638
rect 363052 32574 363104 32580
rect 364628 31414 364656 50487
rect 365718 50416 365774 50425
rect 365718 50351 365774 50360
rect 374366 50416 374422 50425
rect 374366 50351 374422 50360
rect 364616 31408 364668 31414
rect 364616 31350 364668 31356
rect 365732 29986 365760 50351
rect 367282 50280 367338 50289
rect 367282 50215 367338 50224
rect 369950 50280 370006 50289
rect 369950 50215 370006 50224
rect 367098 49736 367154 49745
rect 367098 49671 367154 49680
rect 365720 29980 365772 29986
rect 365720 29922 365772 29928
rect 364984 28484 365036 28490
rect 364984 28426 365036 28432
rect 362972 16546 363552 16574
rect 361120 7744 361172 7750
rect 361120 7686 361172 7692
rect 360844 3596 360896 3602
rect 360844 3538 360896 3544
rect 361132 480 361160 7686
rect 362224 5092 362276 5098
rect 362224 5034 362276 5040
rect 362236 4962 362264 5034
rect 362224 4956 362276 4962
rect 362224 4898 362276 4904
rect 362316 3528 362368 3534
rect 362316 3470 362368 3476
rect 362328 480 362356 3470
rect 363524 480 363552 16546
rect 364616 7812 364668 7818
rect 364616 7754 364668 7760
rect 364628 480 364656 7754
rect 364996 3670 365024 28426
rect 365720 24472 365772 24478
rect 365720 24414 365772 24420
rect 365732 7546 365760 24414
rect 367112 24410 367140 49671
rect 367296 27198 367324 50215
rect 368754 50076 368810 50085
rect 368754 50011 368810 50020
rect 368478 49872 368534 49881
rect 368478 49807 368534 49816
rect 367284 27192 367336 27198
rect 367284 27134 367336 27140
rect 367100 24404 367152 24410
rect 367100 24346 367152 24352
rect 368492 11898 368520 49807
rect 368768 47870 368796 50011
rect 369858 49872 369914 49881
rect 369858 49807 369914 49816
rect 368756 47864 368808 47870
rect 368756 47806 368808 47812
rect 369872 46510 369900 49807
rect 369860 46504 369912 46510
rect 369860 46446 369912 46452
rect 369860 35556 369912 35562
rect 369860 35498 369912 35504
rect 369872 16574 369900 35498
rect 369964 20330 369992 50215
rect 371422 49736 371478 49745
rect 371422 49671 371478 49680
rect 374182 49736 374238 49745
rect 374182 49671 374238 49680
rect 371240 46368 371292 46374
rect 371240 46310 371292 46316
rect 369952 20324 370004 20330
rect 369952 20266 370004 20272
rect 369872 16546 370176 16574
rect 368480 11892 368532 11898
rect 368480 11834 368532 11840
rect 369400 10328 369452 10334
rect 369400 10270 369452 10276
rect 368204 7880 368256 7886
rect 368204 7822 368256 7828
rect 365720 7540 365772 7546
rect 365720 7482 365772 7488
rect 367008 7540 367060 7546
rect 367008 7482 367060 7488
rect 364984 3664 365036 3670
rect 364984 3606 365036 3612
rect 365812 3664 365864 3670
rect 365812 3606 365864 3612
rect 365824 480 365852 3606
rect 367020 480 367048 7482
rect 368216 480 368244 7822
rect 369412 480 369440 10270
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370148 354 370176 16546
rect 370504 11892 370556 11898
rect 370504 11834 370556 11840
rect 370516 3738 370544 11834
rect 370504 3732 370556 3738
rect 370504 3674 370556 3680
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 371252 354 371280 46310
rect 371436 11966 371464 49671
rect 374000 25832 374052 25838
rect 374000 25774 374052 25780
rect 371424 11960 371476 11966
rect 371424 11902 371476 11908
rect 372896 3732 372948 3738
rect 372896 3674 372948 3680
rect 372908 480 372936 3674
rect 374012 3346 374040 25774
rect 374092 12164 374144 12170
rect 374092 12106 374144 12112
rect 374104 3534 374132 12106
rect 374196 5098 374224 49671
rect 374380 12034 374408 50351
rect 376850 50280 376906 50289
rect 376850 50215 376906 50224
rect 379518 50280 379574 50289
rect 379518 50215 379574 50224
rect 375194 49872 375250 49881
rect 375250 49830 375512 49858
rect 375194 49807 375250 49816
rect 375378 49736 375434 49745
rect 375378 49671 375434 49680
rect 375392 49298 375420 49671
rect 375380 49292 375432 49298
rect 375380 49234 375432 49240
rect 375484 45554 375512 49830
rect 375392 45526 375512 45554
rect 375392 39710 375420 45526
rect 376024 40928 376076 40934
rect 376024 40870 376076 40876
rect 375380 39704 375432 39710
rect 375380 39646 375432 39652
rect 374368 12028 374420 12034
rect 374368 11970 374420 11976
rect 374184 5092 374236 5098
rect 374184 5034 374236 5040
rect 374092 3528 374144 3534
rect 374092 3470 374144 3476
rect 375288 3528 375340 3534
rect 375288 3470 375340 3476
rect 374012 3318 374132 3346
rect 374104 480 374132 3318
rect 375300 480 375328 3470
rect 376036 3466 376064 40870
rect 376760 32700 376812 32706
rect 376760 32642 376812 32648
rect 376772 6914 376800 32642
rect 376864 9246 376892 50215
rect 378322 49736 378378 49745
rect 378322 49671 378378 49680
rect 378336 38214 378364 49671
rect 378784 49156 378836 49162
rect 378784 49098 378836 49104
rect 378324 38208 378376 38214
rect 378324 38150 378376 38156
rect 376852 9240 376904 9246
rect 376852 9182 376904 9188
rect 376772 6886 377720 6914
rect 376484 3732 376536 3738
rect 376484 3674 376536 3680
rect 376024 3460 376076 3466
rect 376024 3402 376076 3408
rect 376496 480 376524 3674
rect 377692 480 377720 6886
rect 378796 3670 378824 49098
rect 379532 42430 379560 50215
rect 380070 50008 380126 50017
rect 380070 49943 380126 49952
rect 380084 49745 380112 49943
rect 380898 49872 380954 49881
rect 380898 49807 380954 49816
rect 380070 49736 380126 49745
rect 380070 49671 380126 49680
rect 380912 43790 380940 49807
rect 381082 49736 381138 49745
rect 381082 49671 381138 49680
rect 380900 43784 380952 43790
rect 380900 43726 380952 43732
rect 379520 42424 379572 42430
rect 379520 42366 379572 42372
rect 378876 33924 378928 33930
rect 378876 33866 378928 33872
rect 378888 16574 378916 33866
rect 380900 27124 380952 27130
rect 380900 27066 380952 27072
rect 380912 16574 380940 27066
rect 378888 16546 379008 16574
rect 380912 16546 381032 16574
rect 378876 7948 378928 7954
rect 378876 7890 378928 7896
rect 378784 3664 378836 3670
rect 378784 3606 378836 3612
rect 378888 480 378916 7890
rect 378980 3602 379008 16546
rect 378968 3596 379020 3602
rect 378968 3538 379020 3544
rect 379980 3528 380032 3534
rect 379980 3470 380032 3476
rect 381004 3482 381032 16546
rect 381096 5030 381124 49671
rect 382292 10606 382320 50487
rect 383750 50416 383806 50425
rect 383750 50351 383806 50360
rect 385038 50416 385094 50425
rect 385038 50351 385094 50360
rect 387982 50416 388038 50425
rect 387982 50351 388038 50360
rect 393410 50416 393466 50425
rect 393410 50351 393466 50360
rect 395066 50416 395122 50425
rect 395066 50351 395122 50360
rect 382924 47728 382976 47734
rect 382924 47670 382976 47676
rect 382280 10600 382332 10606
rect 382280 10542 382332 10548
rect 382372 8016 382424 8022
rect 382372 7958 382424 7964
rect 381084 5024 381136 5030
rect 381084 4966 381136 4972
rect 379992 480 380020 3470
rect 381004 3454 381216 3482
rect 381188 480 381216 3454
rect 382384 480 382412 7958
rect 382936 3806 382964 47670
rect 383660 23044 383712 23050
rect 383660 22986 383712 22992
rect 382924 3800 382976 3806
rect 382924 3742 382976 3748
rect 383568 3460 383620 3466
rect 383568 3402 383620 3408
rect 383580 480 383608 3402
rect 383672 626 383700 22986
rect 383764 6798 383792 50351
rect 383934 49872 383990 49881
rect 383934 49807 383990 49816
rect 383948 45218 383976 49807
rect 383936 45212 383988 45218
rect 383936 45154 383988 45160
rect 383752 6792 383804 6798
rect 383752 6734 383804 6740
rect 385052 6662 385080 50351
rect 386510 50280 386566 50289
rect 386510 50215 386566 50224
rect 386420 10396 386472 10402
rect 386420 10338 386472 10344
rect 385040 6656 385092 6662
rect 385040 6598 385092 6604
rect 385960 6316 386012 6322
rect 385960 6258 386012 6264
rect 383672 598 384344 626
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 598
rect 385972 480 386000 6258
rect 386432 490 386460 10338
rect 386524 6594 386552 50215
rect 387798 50008 387854 50017
rect 387798 49943 387854 49952
rect 387812 47938 387840 49943
rect 387800 47932 387852 47938
rect 387800 47874 387852 47880
rect 387800 34060 387852 34066
rect 387800 34002 387852 34008
rect 386512 6588 386564 6594
rect 386512 6530 386564 6536
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 386432 462 386736 490
rect 386708 354 386736 462
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 34002
rect 387996 6458 388024 50351
rect 389178 50280 389234 50289
rect 389178 50215 389234 50224
rect 388166 49872 388222 49881
rect 388166 49807 388222 49816
rect 388180 6526 388208 49807
rect 388168 6520 388220 6526
rect 388168 6462 388220 6468
rect 387984 6452 388036 6458
rect 387984 6394 388036 6400
rect 389192 6390 389220 50215
rect 391938 49872 391994 49881
rect 391938 49807 391994 49816
rect 390742 49736 390798 49745
rect 390742 49671 390798 49680
rect 390756 41070 390784 49671
rect 390744 41064 390796 41070
rect 390744 41006 390796 41012
rect 390560 28552 390612 28558
rect 390560 28494 390612 28500
rect 389456 6520 389508 6526
rect 389456 6462 389508 6468
rect 389180 6384 389232 6390
rect 389180 6326 389232 6332
rect 389468 480 389496 6462
rect 390572 3602 390600 28494
rect 391952 6254 391980 49807
rect 392584 38072 392636 38078
rect 392584 38014 392636 38020
rect 391940 6248 391992 6254
rect 391940 6190 391992 6196
rect 392596 3738 392624 38014
rect 393320 10464 393372 10470
rect 393320 10406 393372 10412
rect 393044 6384 393096 6390
rect 393044 6326 393096 6332
rect 392584 3732 392636 3738
rect 392584 3674 392636 3680
rect 390652 3664 390704 3670
rect 390652 3606 390704 3612
rect 390560 3596 390612 3602
rect 390560 3538 390612 3544
rect 390664 480 390692 3606
rect 391848 3596 391900 3602
rect 391848 3538 391900 3544
rect 391860 480 391888 3538
rect 393056 480 393084 6326
rect 393332 3482 393360 10406
rect 393424 6186 393452 50351
rect 394698 49872 394754 49881
rect 394754 49830 394832 49858
rect 394698 49807 394754 49816
rect 394698 49736 394754 49745
rect 394698 49671 394754 49680
rect 394712 46374 394740 49671
rect 394700 46368 394752 46374
rect 394700 46310 394752 46316
rect 394804 45554 394832 49830
rect 394804 45526 394924 45554
rect 394700 29912 394752 29918
rect 394700 29854 394752 29860
rect 394712 6914 394740 29854
rect 394896 7818 394924 45526
rect 394884 7812 394936 7818
rect 394884 7754 394936 7760
rect 395080 7750 395108 50351
rect 396170 50280 396226 50289
rect 396170 50215 396226 50224
rect 396080 46980 396132 46986
rect 396080 46922 396132 46928
rect 395068 7744 395120 7750
rect 395068 7686 395120 7692
rect 394712 6886 395384 6914
rect 393412 6180 393464 6186
rect 393412 6122 393464 6128
rect 393332 3454 394280 3482
rect 394252 480 394280 3454
rect 395356 480 395384 6886
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 46922
rect 396184 7886 396212 50215
rect 397458 49736 397514 49745
rect 397458 49671 397514 49680
rect 397472 12170 397500 49671
rect 398840 31340 398892 31346
rect 398840 31282 398892 31288
rect 397460 12164 397512 12170
rect 397460 12106 397512 12112
rect 396172 7880 396224 7886
rect 396172 7822 396224 7828
rect 398852 6914 398880 31282
rect 398944 7954 398972 50487
rect 400494 50416 400550 50425
rect 400494 50351 400550 50360
rect 400310 49736 400366 49745
rect 400310 49671 400366 49680
rect 400220 10532 400272 10538
rect 400220 10474 400272 10480
rect 400128 8356 400180 8362
rect 400128 8298 400180 8304
rect 398932 7948 398984 7954
rect 398932 7890 398984 7896
rect 398852 6886 398972 6914
rect 397736 3596 397788 3602
rect 397736 3538 397788 3544
rect 397748 480 397776 3538
rect 398944 480 398972 6886
rect 400140 480 400168 8298
rect 400232 1578 400260 10474
rect 400324 6322 400352 49671
rect 400508 8022 400536 50351
rect 403070 50280 403126 50289
rect 403070 50215 403126 50224
rect 404542 50280 404598 50289
rect 404542 50215 404598 50224
rect 407762 50280 407818 50289
rect 407762 50215 407818 50224
rect 402978 49872 403034 49881
rect 402978 49807 403034 49816
rect 401690 49736 401746 49745
rect 401690 49671 401746 49680
rect 401600 39636 401652 39642
rect 401600 39578 401652 39584
rect 400496 8016 400548 8022
rect 400496 7958 400548 7964
rect 400312 6316 400364 6322
rect 400312 6258 400364 6264
rect 401612 3482 401640 39578
rect 401704 6526 401732 49671
rect 402992 46986 403020 49807
rect 402980 46980 403032 46986
rect 402980 46922 403032 46928
rect 403084 45554 403112 50215
rect 402992 45526 403112 45554
rect 401692 6520 401744 6526
rect 401692 6462 401744 6468
rect 402992 6390 403020 45526
rect 403624 39568 403676 39574
rect 403624 39510 403676 39516
rect 403636 6914 403664 39510
rect 404556 8362 404584 50215
rect 407118 49872 407174 49881
rect 407118 49807 407174 49816
rect 405830 49736 405886 49745
rect 405830 49671 405886 49680
rect 405740 46436 405792 46442
rect 405740 46378 405792 46384
rect 405004 20052 405056 20058
rect 405004 19994 405056 20000
rect 404544 8356 404596 8362
rect 404544 8298 404596 8304
rect 403544 6886 403664 6914
rect 402980 6384 403032 6390
rect 402980 6326 403032 6332
rect 403544 3534 403572 6886
rect 403624 5568 403676 5574
rect 403624 5510 403676 5516
rect 403532 3528 403584 3534
rect 401612 3454 402560 3482
rect 403532 3470 403584 3476
rect 400232 1550 400904 1578
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 1550
rect 402532 480 402560 3454
rect 403636 480 403664 5510
rect 405016 3670 405044 19994
rect 405004 3664 405056 3670
rect 405004 3606 405056 3612
rect 404820 3528 404872 3534
rect 404820 3470 404872 3476
rect 405752 3482 405780 46378
rect 405844 5574 405872 49671
rect 407132 16574 407160 49807
rect 407132 16546 407252 16574
rect 405832 5568 405884 5574
rect 405832 5510 405884 5516
rect 404832 480 404860 3470
rect 405752 3454 406056 3482
rect 406028 480 406056 3454
rect 407224 480 407252 16546
rect 407776 5574 407804 50215
rect 409142 49872 409198 49881
rect 409142 49807 409198 49816
rect 408500 45144 408552 45150
rect 408500 45086 408552 45092
rect 408512 6914 408540 45086
rect 409156 16574 409184 49807
rect 409156 16546 409276 16574
rect 408512 6886 409184 6914
rect 407764 5568 407816 5574
rect 407764 5510 407816 5516
rect 408408 3664 408460 3670
rect 408408 3606 408460 3612
rect 408420 480 408448 3606
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 6886
rect 409248 5642 409276 16546
rect 410536 6526 410564 50623
rect 412086 50552 412142 50561
rect 412086 50487 412142 50496
rect 411902 49736 411958 49745
rect 411902 49671 411958 49680
rect 410616 25696 410668 25702
rect 410616 25638 410668 25644
rect 410524 6520 410576 6526
rect 410524 6462 410576 6468
rect 409236 5636 409288 5642
rect 409236 5578 409288 5584
rect 410628 3466 410656 25638
rect 411260 22840 411312 22846
rect 411260 22782 411312 22788
rect 411272 6914 411300 22782
rect 411916 16574 411944 49671
rect 411916 16546 412036 16574
rect 411272 6886 411944 6914
rect 410800 5568 410852 5574
rect 410800 5510 410852 5516
rect 410616 3460 410668 3466
rect 410616 3402 410668 3408
rect 410812 480 410840 5510
rect 411916 480 411944 6886
rect 412008 6390 412036 16546
rect 412100 6458 412128 50487
rect 416686 50416 416742 50425
rect 416686 50351 416742 50360
rect 420182 50416 420238 50425
rect 420182 50351 420238 50360
rect 413282 50280 413338 50289
rect 413282 50215 413338 50224
rect 412546 50008 412602 50017
rect 412546 49943 412602 49952
rect 412560 49745 412588 49943
rect 412546 49736 412602 49745
rect 412546 49671 412602 49680
rect 412640 49224 412692 49230
rect 412640 49166 412692 49172
rect 412088 6452 412140 6458
rect 412088 6394 412140 6400
rect 411996 6384 412048 6390
rect 411996 6326 412048 6332
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 49166
rect 413296 6322 413324 50215
rect 414846 49872 414902 49881
rect 414846 49807 414902 49816
rect 414662 49736 414718 49745
rect 414662 49671 414718 49680
rect 413284 6316 413336 6322
rect 413284 6258 413336 6264
rect 414676 6186 414704 49671
rect 414860 6254 414888 49807
rect 416700 46374 416728 50351
rect 417422 50280 417478 50289
rect 417422 50215 417478 50224
rect 416688 46368 416740 46374
rect 416688 46310 416740 46316
rect 415400 38140 415452 38146
rect 415400 38082 415452 38088
rect 414848 6248 414900 6254
rect 414848 6190 414900 6196
rect 414664 6180 414716 6186
rect 414664 6122 414716 6128
rect 414296 5636 414348 5642
rect 414296 5578 414348 5584
rect 414308 480 414336 5578
rect 415412 3466 415440 38082
rect 417436 7886 417464 50215
rect 418802 49872 418858 49881
rect 418802 49807 418858 49816
rect 417606 49736 417662 49745
rect 417606 49671 417662 49680
rect 417424 7880 417476 7886
rect 417424 7822 417476 7828
rect 417620 7818 417648 49671
rect 418528 10600 418580 10606
rect 418528 10542 418580 10548
rect 417608 7812 417660 7818
rect 417608 7754 417660 7760
rect 417884 6520 417936 6526
rect 417884 6462 417936 6468
rect 415492 3800 415544 3806
rect 415492 3742 415544 3748
rect 415400 3460 415452 3466
rect 415400 3402 415452 3408
rect 415504 480 415532 3742
rect 416688 3460 416740 3466
rect 416688 3402 416740 3408
rect 416700 480 416728 3402
rect 417896 480 417924 6462
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418540 354 418568 10542
rect 418816 7750 418844 49807
rect 418896 44940 418948 44946
rect 418896 44882 418948 44888
rect 418804 7744 418856 7750
rect 418804 7686 418856 7692
rect 418908 3602 418936 44882
rect 420196 16574 420224 50351
rect 421760 50153 421788 50623
rect 422942 50280 422998 50289
rect 422942 50215 422998 50224
rect 421746 50144 421802 50153
rect 421746 50079 421802 50088
rect 421562 49872 421618 49881
rect 421562 49807 421618 49816
rect 420196 16546 420316 16574
rect 420288 7682 420316 16546
rect 421576 8158 421604 49807
rect 421746 49736 421802 49745
rect 421746 49671 421802 49680
rect 421760 9382 421788 49671
rect 421748 9376 421800 9382
rect 421748 9318 421800 9324
rect 422956 9314 422984 50215
rect 424322 49600 424378 49609
rect 424322 49535 424378 49544
rect 422944 9308 422996 9314
rect 422944 9250 422996 9256
rect 424336 9178 424364 49535
rect 424520 9246 424548 50623
rect 427082 50552 427138 50561
rect 427082 50487 427138 50496
rect 425702 49736 425758 49745
rect 425702 49671 425758 49680
rect 425520 10668 425572 10674
rect 425520 10610 425572 10616
rect 424508 9240 424560 9246
rect 424508 9182 424560 9188
rect 424324 9172 424376 9178
rect 424324 9114 424376 9120
rect 421564 8152 421616 8158
rect 421564 8094 421616 8100
rect 420184 7676 420236 7682
rect 420184 7618 420236 7624
rect 420276 7676 420328 7682
rect 420276 7618 420328 7624
rect 418896 3596 418948 3602
rect 418896 3538 418948 3544
rect 420196 480 420224 7618
rect 423772 7608 423824 7614
rect 423772 7550 423824 7556
rect 421380 6452 421432 6458
rect 421380 6394 421432 6400
rect 421392 480 421420 6394
rect 422576 3460 422628 3466
rect 422576 3402 422628 3408
rect 422588 480 422616 3402
rect 423784 480 423812 7550
rect 424968 6384 425020 6390
rect 424968 6326 425020 6332
rect 424980 480 425008 6326
rect 425532 490 425560 10610
rect 425716 6914 425744 49671
rect 426440 47796 426492 47802
rect 426440 47738 426492 47744
rect 425796 32632 425848 32638
rect 425796 32574 425848 32580
rect 425624 6886 425744 6914
rect 425624 4962 425652 6886
rect 425612 4956 425664 4962
rect 425612 4898 425664 4904
rect 425808 3670 425836 32574
rect 426452 16574 426480 47738
rect 426452 16546 426848 16574
rect 425796 3664 425848 3670
rect 425796 3606 425848 3612
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425532 462 425744 490
rect 425716 354 425744 462
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 16546
rect 427096 9110 427124 50487
rect 428462 50416 428518 50425
rect 428462 50351 428518 50360
rect 427084 9104 427136 9110
rect 427084 9046 427136 9052
rect 428476 6594 428504 50351
rect 429750 50280 429806 50289
rect 429750 50215 429806 50224
rect 429658 50008 429714 50017
rect 429658 49943 429714 49952
rect 429672 49745 429700 49943
rect 428646 49736 428702 49745
rect 428646 49671 428702 49680
rect 429658 49736 429714 49745
rect 429658 49671 429714 49680
rect 428464 6588 428516 6594
rect 428464 6530 428516 6536
rect 428660 6526 428688 49671
rect 429764 45554 429792 50215
rect 431328 50153 431356 50623
rect 432602 50416 432658 50425
rect 432602 50351 432658 50360
rect 431314 50144 431370 50153
rect 431314 50079 431370 50088
rect 431406 49872 431462 49881
rect 431406 49807 431462 49816
rect 431222 49736 431278 49745
rect 431222 49671 431278 49680
rect 429764 45526 429884 45554
rect 428648 6520 428700 6526
rect 428648 6462 428700 6468
rect 429856 6458 429884 45526
rect 430580 42356 430632 42362
rect 430580 42298 430632 42304
rect 429936 42288 429988 42294
rect 429936 42230 429988 42236
rect 429844 6452 429896 6458
rect 429844 6394 429896 6400
rect 428464 6316 428516 6322
rect 428464 6258 428516 6264
rect 428476 480 428504 6258
rect 429948 3534 429976 42230
rect 430592 16574 430620 42298
rect 430592 16546 430896 16574
rect 429936 3528 429988 3534
rect 429936 3470 429988 3476
rect 429658 3360 429714 3369
rect 429658 3295 429714 3304
rect 429672 480 429700 3295
rect 430868 480 430896 16546
rect 431236 6322 431264 49671
rect 431420 6390 431448 49807
rect 431408 6384 431460 6390
rect 431408 6326 431460 6332
rect 431224 6316 431276 6322
rect 431224 6258 431276 6264
rect 432616 6254 432644 50351
rect 433982 50280 434038 50289
rect 433982 50215 434038 50224
rect 433996 24342 434024 50215
rect 434640 47802 434668 50623
rect 441066 50416 441122 50425
rect 441066 50351 441122 50360
rect 445666 50416 445722 50425
rect 445666 50351 445722 50360
rect 438122 50280 438178 50289
rect 438122 50215 438178 50224
rect 436466 50008 436522 50017
rect 436466 49943 436522 49952
rect 435362 49736 435418 49745
rect 435362 49671 435418 49680
rect 434628 47796 434680 47802
rect 434628 47738 434680 47744
rect 433340 24336 433392 24342
rect 433340 24278 433392 24284
rect 433984 24336 434036 24342
rect 433984 24278 434036 24284
rect 433352 16574 433380 24278
rect 433352 16546 434024 16574
rect 432052 6248 432104 6254
rect 432052 6190 432104 6196
rect 432604 6248 432656 6254
rect 432604 6190 432656 6196
rect 432064 480 432092 6190
rect 433248 3528 433300 3534
rect 433248 3470 433300 3476
rect 433260 480 433288 3470
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 435376 11966 435404 49671
rect 436480 49298 436508 49943
rect 436558 49872 436614 49881
rect 436558 49807 436614 49816
rect 436468 49292 436520 49298
rect 436468 49234 436520 49240
rect 436572 45554 436600 49807
rect 436572 45526 436784 45554
rect 435364 11960 435416 11966
rect 435364 11902 435416 11908
rect 436756 6186 436784 45526
rect 438136 25770 438164 50215
rect 440422 49872 440478 49881
rect 440422 49807 440478 49816
rect 439502 49736 439558 49745
rect 439502 49671 439558 49680
rect 438860 46368 438912 46374
rect 438860 46310 438912 46316
rect 437480 25764 437532 25770
rect 437480 25706 437532 25712
rect 438124 25764 438176 25770
rect 438124 25706 438176 25712
rect 435548 6180 435600 6186
rect 435548 6122 435600 6128
rect 436744 6180 436796 6186
rect 436744 6122 436796 6128
rect 435560 480 435588 6122
rect 436744 3596 436796 3602
rect 436744 3538 436796 3544
rect 436756 480 436784 3538
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 434414 -960 434526 326
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437492 354 437520 25706
rect 438872 16574 438900 46310
rect 439516 23050 439544 49671
rect 440436 45554 440464 49807
rect 440436 45526 440924 45554
rect 440240 43648 440292 43654
rect 440240 43590 440292 43596
rect 439504 23044 439556 23050
rect 439504 22986 439556 22992
rect 438872 16546 439176 16574
rect 439148 480 439176 16546
rect 440252 3398 440280 43590
rect 440896 29782 440924 45526
rect 441080 31210 441108 50351
rect 442262 49872 442318 49881
rect 442262 49807 442318 49816
rect 441068 31204 441120 31210
rect 441068 31146 441120 31152
rect 440884 29776 440936 29782
rect 440884 29718 440936 29724
rect 442276 27130 442304 49807
rect 445022 49736 445078 49745
rect 445022 49671 445078 49680
rect 443734 49600 443790 49609
rect 443734 49535 443790 49544
rect 443644 43648 443696 43654
rect 443644 43590 443696 43596
rect 442264 27124 442316 27130
rect 442264 27066 442316 27072
rect 442632 7880 442684 7886
rect 442632 7822 442684 7828
rect 440332 3664 440384 3670
rect 440332 3606 440384 3612
rect 440240 3392 440292 3398
rect 440240 3334 440292 3340
rect 440344 480 440372 3606
rect 441528 3392 441580 3398
rect 441528 3334 441580 3340
rect 441540 480 441568 3334
rect 442644 480 442672 7822
rect 443656 3806 443684 43590
rect 443748 38146 443776 49535
rect 443736 38140 443788 38146
rect 443736 38082 443788 38088
rect 445036 32706 445064 49671
rect 445680 46374 445708 50351
rect 446310 50280 446366 50289
rect 446310 50215 446366 50224
rect 446218 50008 446274 50017
rect 446218 49943 446274 49952
rect 446232 49745 446260 49943
rect 446218 49736 446274 49745
rect 446218 49671 446274 49680
rect 445668 46368 445720 46374
rect 445668 46310 445720 46316
rect 446324 45554 446352 50215
rect 447966 49872 448022 49881
rect 447966 49807 448022 49816
rect 447782 49736 447838 49745
rect 447782 49671 447838 49680
rect 446324 45526 446444 45554
rect 445024 32700 445076 32706
rect 445024 32642 445076 32648
rect 444380 22976 444432 22982
rect 444380 22918 444432 22924
rect 444392 16574 444420 22918
rect 444392 16546 445064 16574
rect 443644 3800 443696 3806
rect 443644 3742 443696 3748
rect 443828 3732 443880 3738
rect 443828 3674 443880 3680
rect 443840 480 443868 3674
rect 445036 480 445064 16546
rect 446416 8090 446444 45526
rect 446404 8084 446456 8090
rect 446404 8026 446456 8032
rect 447796 7954 447824 49671
rect 447980 8022 448008 49807
rect 448520 40860 448572 40866
rect 448520 40802 448572 40808
rect 448532 16574 448560 40802
rect 448532 16546 448652 16574
rect 447968 8016 448020 8022
rect 447968 7958 448020 7964
rect 447784 7948 447836 7954
rect 447784 7890 447836 7896
rect 446220 7812 446272 7818
rect 446220 7754 446272 7760
rect 446232 480 446260 7754
rect 447416 3800 447468 3806
rect 447416 3742 447468 3748
rect 447428 480 447456 3742
rect 448624 480 448652 16546
rect 449176 13394 449204 50759
rect 450542 50688 450598 50697
rect 450542 50623 450598 50632
rect 461030 50688 461086 50697
rect 461030 50623 461086 50632
rect 498290 50688 498346 50697
rect 498290 50623 498346 50632
rect 545210 50688 545266 50697
rect 545210 50623 545266 50632
rect 449164 13388 449216 13394
rect 449164 13330 449216 13336
rect 450556 7886 450584 50623
rect 453302 50552 453358 50561
rect 453302 50487 453358 50496
rect 451922 49872 451978 49881
rect 451922 49807 451978 49816
rect 450726 49736 450782 49745
rect 450726 49671 450782 49680
rect 450544 7880 450596 7886
rect 450544 7822 450596 7828
rect 450740 7818 450768 49671
rect 451280 36712 451332 36718
rect 451280 36654 451332 36660
rect 451292 16574 451320 36654
rect 451292 16546 451688 16574
rect 450912 9036 450964 9042
rect 450912 8978 450964 8984
rect 450728 7812 450780 7818
rect 450728 7754 450780 7760
rect 449808 7744 449860 7750
rect 449808 7686 449860 7692
rect 449820 480 449848 7686
rect 450924 480 450952 8978
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 451936 7750 451964 49807
rect 453316 16574 453344 50487
rect 454682 50416 454738 50425
rect 454682 50351 454738 50360
rect 454406 50008 454462 50017
rect 454406 49943 454462 49952
rect 454038 49736 454094 49745
rect 454038 49671 454094 49680
rect 453316 16546 453436 16574
rect 451924 7744 451976 7750
rect 451924 7686 451976 7692
rect 453408 7682 453436 16546
rect 454052 13122 454080 49671
rect 454420 47598 454448 49943
rect 454408 47592 454460 47598
rect 454408 47534 454460 47540
rect 454040 13116 454092 13122
rect 454040 13058 454092 13064
rect 453304 7676 453356 7682
rect 453304 7618 453356 7624
rect 453396 7676 453448 7682
rect 453396 7618 453448 7624
rect 453316 480 453344 7618
rect 454696 7614 454724 50351
rect 456982 50280 457038 50289
rect 456982 50215 457038 50224
rect 455510 49872 455566 49881
rect 455510 49807 455566 49816
rect 455420 35352 455472 35358
rect 455420 35294 455472 35300
rect 455432 16574 455460 35294
rect 455524 28286 455552 49807
rect 456996 32434 457024 50215
rect 458270 49736 458326 49745
rect 458270 49671 458326 49680
rect 459558 49736 459614 49745
rect 459558 49671 459614 49680
rect 458180 32564 458232 32570
rect 458180 32506 458232 32512
rect 456984 32428 457036 32434
rect 456984 32370 457036 32376
rect 455512 28280 455564 28286
rect 455512 28222 455564 28228
rect 458192 16574 458220 32506
rect 458284 17270 458312 49671
rect 459572 17338 459600 49671
rect 461044 24138 461072 50623
rect 462410 50552 462466 50561
rect 462410 50487 462466 50496
rect 491298 50552 491354 50561
rect 491298 50487 491354 50496
rect 461214 49872 461270 49881
rect 461214 49807 461270 49816
rect 461032 24132 461084 24138
rect 461032 24074 461084 24080
rect 461228 17406 461256 49807
rect 462320 27056 462372 27062
rect 462320 26998 462372 27004
rect 461216 17400 461268 17406
rect 461216 17342 461268 17348
rect 459560 17332 459612 17338
rect 459560 17274 459612 17280
rect 458272 17264 458324 17270
rect 458272 17206 458324 17212
rect 455432 16546 455736 16574
rect 458192 16546 459232 16574
rect 454684 7608 454736 7614
rect 454684 7550 454736 7556
rect 454500 3868 454552 3874
rect 454500 3810 454552 3816
rect 454512 480 454540 3810
rect 455708 480 455736 16546
rect 456892 8152 456944 8158
rect 456892 8094 456944 8100
rect 456904 480 456932 8094
rect 458088 3936 458140 3942
rect 458088 3878 458140 3884
rect 458100 480 458128 3878
rect 459204 480 459232 16546
rect 460388 9376 460440 9382
rect 460388 9318 460440 9324
rect 460400 480 460428 9318
rect 461584 4004 461636 4010
rect 461584 3946 461636 3952
rect 461596 480 461624 3946
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462332 354 462360 26998
rect 462424 17474 462452 50487
rect 463790 50416 463846 50425
rect 463790 50351 463846 50360
rect 466550 50416 466606 50425
rect 466550 50351 466606 50360
rect 470690 50416 470746 50425
rect 470690 50351 470746 50360
rect 470966 50416 471022 50425
rect 470966 50351 471022 50360
rect 473358 50416 473414 50425
rect 473358 50351 473414 50360
rect 476486 50416 476542 50425
rect 476486 50351 476542 50360
rect 478878 50416 478934 50425
rect 478878 50351 478934 50360
rect 483294 50416 483350 50425
rect 483294 50351 483350 50360
rect 488538 50416 488594 50425
rect 488538 50351 488594 50360
rect 463804 17542 463832 50351
rect 465170 50280 465226 50289
rect 465170 50215 465226 50224
rect 463974 49736 464030 49745
rect 463974 49671 464030 49680
rect 463792 17536 463844 17542
rect 463792 17478 463844 17484
rect 462412 17468 462464 17474
rect 462412 17410 462464 17416
rect 463988 13190 464016 49671
rect 465080 33992 465132 33998
rect 465080 33934 465132 33940
rect 465092 16574 465120 33934
rect 465184 29646 465212 50215
rect 465172 29640 465224 29646
rect 465172 29582 465224 29588
rect 465092 16546 465856 16574
rect 463976 13184 464028 13190
rect 463976 13126 464028 13132
rect 463976 9308 464028 9314
rect 463976 9250 464028 9256
rect 463988 480 464016 9250
rect 465172 4072 465224 4078
rect 465172 4014 465224 4020
rect 465184 480 465212 4014
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 354 465856 16546
rect 466564 13326 466592 50351
rect 467654 50280 467710 50289
rect 467710 50238 467880 50266
rect 467654 50215 467710 50224
rect 466734 49872 466790 49881
rect 466734 49807 466790 49816
rect 466552 13320 466604 13326
rect 466552 13262 466604 13268
rect 466748 13258 466776 49807
rect 467852 36582 467880 50238
rect 469218 49736 469274 49745
rect 469218 49671 469274 49680
rect 470598 49736 470654 49745
rect 470598 49671 470654 49680
rect 467840 36576 467892 36582
rect 467840 36518 467892 36524
rect 469232 35222 469260 49671
rect 470612 49026 470640 49671
rect 470600 49020 470652 49026
rect 470600 48962 470652 48968
rect 469220 35216 469272 35222
rect 469220 35158 469272 35164
rect 470704 33794 470732 50351
rect 470980 50153 471008 50351
rect 471978 50280 472034 50289
rect 471978 50215 472034 50224
rect 470966 50144 471022 50153
rect 470966 50079 471022 50088
rect 470874 49872 470930 49881
rect 470874 49807 470930 49816
rect 470692 33788 470744 33794
rect 470692 33730 470744 33736
rect 470888 31074 470916 49807
rect 471992 39370 472020 50215
rect 473372 42090 473400 50351
rect 474462 49736 474518 49745
rect 476302 49736 476358 49745
rect 474518 49694 474780 49722
rect 474462 49671 474518 49680
rect 473360 42084 473412 42090
rect 473360 42026 473412 42032
rect 471980 39364 472032 39370
rect 471980 39306 472032 39312
rect 470876 31068 470928 31074
rect 470876 31010 470928 31016
rect 473360 28416 473412 28422
rect 473360 28358 473412 28364
rect 473372 16574 473400 28358
rect 474752 25566 474780 49694
rect 476302 49671 476358 49680
rect 476120 45008 476172 45014
rect 476120 44950 476172 44956
rect 474740 25560 474792 25566
rect 474740 25502 474792 25508
rect 473372 16546 473492 16574
rect 466736 13252 466788 13258
rect 466736 13194 466788 13200
rect 467472 9240 467524 9246
rect 467472 9182 467524 9188
rect 467484 480 467512 9182
rect 471060 9172 471112 9178
rect 471060 9114 471112 9120
rect 469864 8968 469916 8974
rect 469864 8910 469916 8916
rect 468668 4140 468720 4146
rect 468668 4082 468720 4088
rect 468680 480 468708 4082
rect 469876 480 469904 8910
rect 471072 480 471100 9114
rect 472256 3392 472308 3398
rect 472256 3334 472308 3340
rect 472268 480 472296 3334
rect 473464 480 473492 16546
rect 476132 6914 476160 44950
rect 476316 14550 476344 49671
rect 476304 14544 476356 14550
rect 476304 14486 476356 14492
rect 476500 14482 476528 50351
rect 477498 49736 477554 49745
rect 477498 49671 477554 49680
rect 477512 14618 477540 49671
rect 478892 14686 478920 50351
rect 480350 50280 480406 50289
rect 480406 50238 480484 50266
rect 480350 50215 480406 50224
rect 480258 50008 480314 50017
rect 480258 49943 480314 49952
rect 480272 49745 480300 49943
rect 480350 49872 480406 49881
rect 480350 49807 480406 49816
rect 480258 49736 480314 49745
rect 480258 49671 480314 49680
rect 480364 43450 480392 49807
rect 480456 45554 480484 50238
rect 481362 49736 481418 49745
rect 483110 49736 483166 49745
rect 481418 49694 481680 49722
rect 481362 49671 481418 49680
rect 480456 45526 480576 45554
rect 480352 43444 480404 43450
rect 480352 43386 480404 43392
rect 480260 18760 480312 18766
rect 480260 18702 480312 18708
rect 480272 16574 480300 18702
rect 480548 18630 480576 45526
rect 480536 18624 480588 18630
rect 480536 18566 480588 18572
rect 480272 16546 480576 16574
rect 478880 14680 478932 14686
rect 478880 14622 478932 14628
rect 477500 14612 477552 14618
rect 477500 14554 477552 14560
rect 476488 14476 476540 14482
rect 476488 14418 476540 14424
rect 478144 9104 478196 9110
rect 478144 9046 478196 9052
rect 476132 6886 476528 6914
rect 474556 4956 474608 4962
rect 474556 4898 474608 4904
rect 474568 480 474596 4898
rect 475752 3324 475804 3330
rect 475752 3266 475804 3272
rect 475764 480 475792 3266
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476500 354 476528 6886
rect 478156 480 478184 9046
rect 479340 3256 479392 3262
rect 479340 3198 479392 3204
rect 479352 480 479380 3198
rect 480548 480 480576 16546
rect 481652 14754 481680 49694
rect 483110 49671 483166 49680
rect 483020 20188 483072 20194
rect 483020 20130 483072 20136
rect 481640 14748 481692 14754
rect 481640 14690 481692 14696
rect 483032 6914 483060 20130
rect 483124 14890 483152 49671
rect 483112 14884 483164 14890
rect 483112 14826 483164 14832
rect 483308 14822 483336 50351
rect 484306 50280 484362 50289
rect 484362 50238 484440 50266
rect 484306 50215 484362 50224
rect 484412 21486 484440 50238
rect 484582 50008 484638 50017
rect 484582 49943 484638 49952
rect 484596 46238 484624 49943
rect 487434 49872 487490 49881
rect 487434 49807 487490 49816
rect 485778 49736 485834 49745
rect 485778 49671 485834 49680
rect 484584 46232 484636 46238
rect 484584 46174 484636 46180
rect 485792 40730 485820 49671
rect 485780 40724 485832 40730
rect 485780 40666 485832 40672
rect 487448 37942 487476 49807
rect 487436 37936 487488 37942
rect 487436 37878 487488 37884
rect 487160 21548 487212 21554
rect 487160 21490 487212 21496
rect 484400 21480 484452 21486
rect 484400 21422 484452 21428
rect 483296 14816 483348 14822
rect 483296 14758 483348 14764
rect 483032 6886 484072 6914
rect 481732 6588 481784 6594
rect 481732 6530 481784 6536
rect 481744 480 481772 6530
rect 482836 4956 482888 4962
rect 482836 4898 482888 4904
rect 482848 480 482876 4898
rect 484044 480 484072 6886
rect 485228 6520 485280 6526
rect 485228 6462 485280 6468
rect 485240 480 485268 6462
rect 486424 5024 486476 5030
rect 486424 4966 486476 4972
rect 486436 480 486464 4966
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487172 354 487200 21490
rect 488552 11762 488580 50351
rect 490194 49872 490250 49881
rect 490194 49807 490250 49816
rect 490010 49736 490066 49745
rect 490010 49671 490066 49680
rect 490024 24206 490052 49671
rect 490012 24200 490064 24206
rect 490012 24142 490064 24148
rect 489920 22908 489972 22914
rect 489920 22850 489972 22856
rect 489932 16574 489960 22850
rect 490208 22778 490236 49807
rect 490196 22772 490248 22778
rect 490196 22714 490248 22720
rect 491312 20126 491340 50487
rect 492862 50280 492918 50289
rect 492862 50215 492918 50224
rect 495438 50280 495494 50289
rect 495438 50215 495494 50224
rect 492678 49736 492734 49745
rect 492678 49671 492734 49680
rect 491300 20120 491352 20126
rect 491300 20062 491352 20068
rect 489932 16546 490696 16574
rect 488540 11756 488592 11762
rect 488540 11698 488592 11704
rect 488816 6452 488868 6458
rect 488816 6394 488868 6400
rect 488828 480 488856 6394
rect 489920 5092 489972 5098
rect 489920 5034 489972 5040
rect 489932 480 489960 5034
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490668 354 490696 16546
rect 492692 15910 492720 49671
rect 492876 26926 492904 50215
rect 494150 49736 494206 49745
rect 494150 49671 494206 49680
rect 494060 47660 494112 47666
rect 494060 47602 494112 47608
rect 492864 26920 492916 26926
rect 492864 26862 492916 26868
rect 492680 15904 492732 15910
rect 492680 15846 492732 15852
rect 494072 6914 494100 47602
rect 494164 15978 494192 49671
rect 495452 16046 495480 50215
rect 495898 50008 495954 50017
rect 495898 49943 495954 49952
rect 495912 49745 495940 49943
rect 496910 49872 496966 49881
rect 496910 49807 496966 49816
rect 495898 49736 495954 49745
rect 495898 49671 495954 49680
rect 496924 16114 496952 49807
rect 497094 49736 497150 49745
rect 497094 49671 497150 49680
rect 497108 16182 497136 49671
rect 498200 24268 498252 24274
rect 498200 24210 498252 24216
rect 497096 16176 497148 16182
rect 497096 16118 497148 16124
rect 496912 16108 496964 16114
rect 496912 16050 496964 16056
rect 495440 16040 495492 16046
rect 495440 15982 495492 15988
rect 494152 15972 494204 15978
rect 494152 15914 494204 15920
rect 494072 6886 494744 6914
rect 492312 6384 492364 6390
rect 492312 6326 492364 6332
rect 492324 480 492352 6326
rect 493508 5160 493560 5166
rect 493508 5102 493560 5108
rect 493520 480 493548 5102
rect 494716 480 494744 6886
rect 495900 6316 495952 6322
rect 495900 6258 495952 6264
rect 495912 480 495940 6258
rect 497096 5228 497148 5234
rect 497096 5170 497148 5176
rect 497108 480 497136 5170
rect 498212 480 498240 24210
rect 498304 16250 498332 50623
rect 499670 50552 499726 50561
rect 499670 50487 499726 50496
rect 501050 50552 501106 50561
rect 501050 50487 501106 50496
rect 507950 50552 508006 50561
rect 507950 50487 508006 50496
rect 514850 50552 514906 50561
rect 514850 50487 514906 50496
rect 530030 50552 530086 50561
rect 530030 50487 530086 50496
rect 499684 16386 499712 50487
rect 499854 49872 499910 49881
rect 499854 49807 499910 49816
rect 499672 16380 499724 16386
rect 499672 16322 499724 16328
rect 499868 16318 499896 49807
rect 500960 25628 501012 25634
rect 500960 25570 501012 25576
rect 499856 16312 499908 16318
rect 499856 16254 499908 16260
rect 498292 16244 498344 16250
rect 498292 16186 498344 16192
rect 500972 6914 501000 25570
rect 501064 16454 501092 50487
rect 503718 50416 503774 50425
rect 503718 50351 503774 50360
rect 502338 49736 502394 49745
rect 502338 49671 502394 49680
rect 502352 45082 502380 49671
rect 502432 47796 502484 47802
rect 502432 47738 502484 47744
rect 502340 45076 502392 45082
rect 502340 45018 502392 45024
rect 502444 16574 502472 47738
rect 503732 17610 503760 50351
rect 505098 50280 505154 50289
rect 505098 50215 505154 50224
rect 503902 49736 503958 49745
rect 503902 49671 503958 49680
rect 503916 39506 503944 49671
rect 503904 39500 503956 39506
rect 503904 39442 503956 39448
rect 505112 29850 505140 50215
rect 505650 50008 505706 50017
rect 505650 49943 505706 49952
rect 505664 49745 505692 49943
rect 506570 49872 506626 49881
rect 506570 49807 506626 49816
rect 505650 49736 505706 49745
rect 505650 49671 505706 49680
rect 505100 29844 505152 29850
rect 505100 29786 505152 29792
rect 505100 26988 505152 26994
rect 505100 26930 505152 26936
rect 503720 17604 503772 17610
rect 503720 17546 503772 17552
rect 505112 16574 505140 26930
rect 506480 24336 506532 24342
rect 506480 24278 506532 24284
rect 502444 16546 503024 16574
rect 505112 16546 505416 16574
rect 501052 16448 501104 16454
rect 501052 16390 501104 16396
rect 500972 6886 501368 6914
rect 499396 6248 499448 6254
rect 499396 6190 499448 6196
rect 499408 480 499436 6190
rect 500592 5296 500644 5302
rect 500592 5238 500644 5244
rect 500604 480 500632 5238
rect 491086 354 491198 480
rect 490668 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501340 354 501368 6886
rect 502996 480 503024 16546
rect 504180 5364 504232 5370
rect 504180 5306 504232 5312
rect 504192 480 504220 5306
rect 505388 480 505416 16546
rect 506492 480 506520 24278
rect 506584 17678 506612 49807
rect 506754 49736 506810 49745
rect 506754 49671 506810 49680
rect 506768 31278 506796 49671
rect 506756 31272 506808 31278
rect 506756 31214 506808 31220
rect 507860 28348 507912 28354
rect 507860 28290 507912 28296
rect 506572 17672 506624 17678
rect 506572 17614 506624 17620
rect 507872 16574 507900 28290
rect 507964 17746 507992 50487
rect 509514 50416 509570 50425
rect 509514 50351 509570 50360
rect 509330 49736 509386 49745
rect 509330 49671 509386 49680
rect 509344 43586 509372 49671
rect 509332 43580 509384 43586
rect 509332 43522 509384 43528
rect 509528 42226 509556 50351
rect 512090 50280 512146 50289
rect 512090 50215 512146 50224
rect 510710 49736 510766 49745
rect 510710 49671 510766 49680
rect 510620 47592 510672 47598
rect 510620 47534 510672 47540
rect 509516 42220 509568 42226
rect 509516 42162 509568 42168
rect 507952 17740 508004 17746
rect 507952 17682 508004 17688
rect 510632 16574 510660 47534
rect 510724 36786 510752 49671
rect 510712 36780 510764 36786
rect 510712 36722 510764 36728
rect 512000 29708 512052 29714
rect 512000 29650 512052 29656
rect 507872 16546 508912 16574
rect 510632 16546 511304 16574
rect 507216 14476 507268 14482
rect 507216 14418 507268 14424
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 354 507256 14418
rect 508884 480 508912 16546
rect 509608 11960 509660 11966
rect 509608 11902 509660 11908
rect 507646 354 507758 480
rect 507228 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 11902
rect 511276 480 511304 16546
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 29650
rect 512104 18834 512132 50215
rect 512458 50008 512514 50017
rect 512458 49943 512514 49952
rect 512472 49745 512500 49943
rect 513654 49872 513710 49881
rect 513654 49807 513710 49816
rect 512458 49736 512514 49745
rect 512458 49671 512514 49680
rect 513470 49736 513526 49745
rect 513470 49671 513526 49680
rect 513484 35426 513512 49671
rect 513472 35420 513524 35426
rect 513472 35362 513524 35368
rect 512092 18828 512144 18834
rect 512092 18770 512144 18776
rect 513668 11830 513696 49807
rect 514760 31136 514812 31142
rect 514760 31078 514812 31084
rect 514772 16574 514800 31078
rect 514864 21622 514892 50487
rect 516138 50416 516194 50425
rect 516138 50351 516194 50360
rect 518990 50416 519046 50425
rect 518990 50351 519046 50360
rect 516152 28490 516180 50351
rect 517702 50008 517758 50017
rect 517702 49943 517758 49952
rect 517518 49872 517574 49881
rect 517518 49807 517574 49816
rect 516322 49736 516378 49745
rect 516322 49671 516378 49680
rect 516336 40934 516364 49671
rect 516324 40928 516376 40934
rect 516324 40870 516376 40876
rect 516140 28484 516192 28490
rect 516140 28426 516192 28432
rect 516140 25764 516192 25770
rect 516140 25706 516192 25712
rect 514852 21616 514904 21622
rect 514852 21558 514904 21564
rect 516152 16574 516180 25706
rect 514772 16546 515536 16574
rect 516152 16546 517192 16574
rect 513656 11824 513708 11830
rect 513656 11766 513708 11772
rect 513564 6180 513616 6186
rect 513564 6122 513616 6128
rect 514760 6180 514812 6186
rect 514760 6122 514812 6128
rect 513576 480 513604 6122
rect 514772 480 514800 6122
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 512430 -960 512542 326
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515508 354 515536 16546
rect 517164 480 517192 16546
rect 517532 11898 517560 49807
rect 517716 49162 517744 49943
rect 517704 49156 517756 49162
rect 517704 49098 517756 49104
rect 518900 49088 518952 49094
rect 518900 49030 518952 49036
rect 518912 16574 518940 49030
rect 519004 33930 519032 50351
rect 520278 50280 520334 50289
rect 523038 50280 523094 50289
rect 520334 50238 520412 50266
rect 520278 50215 520334 50224
rect 519174 49736 519230 49745
rect 519174 49671 519230 49680
rect 519188 47734 519216 49671
rect 520280 49292 520332 49298
rect 520280 49234 520332 49240
rect 519176 47728 519228 47734
rect 519176 47670 519228 47676
rect 518992 33924 519044 33930
rect 518992 33866 519044 33872
rect 518912 16546 519584 16574
rect 517520 11892 517572 11898
rect 517520 11834 517572 11840
rect 517888 11756 517940 11762
rect 517888 11698 517940 11704
rect 515926 354 516038 480
rect 515508 326 516038 354
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 517900 354 517928 11698
rect 519556 480 519584 16546
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 49234
rect 520384 10334 520412 50238
rect 523038 50215 523094 50224
rect 525890 50280 525946 50289
rect 525890 50215 525946 50224
rect 527086 50280 527142 50289
rect 527142 50238 527220 50266
rect 527086 50215 527142 50224
rect 521752 49020 521804 49026
rect 521752 48962 521804 48968
rect 521764 16574 521792 48962
rect 523052 38078 523080 50215
rect 524142 49872 524198 49881
rect 524198 49830 524460 49858
rect 524142 49807 524198 49816
rect 523222 49736 523278 49745
rect 523222 49671 523278 49680
rect 523236 39574 523264 49671
rect 524432 45554 524460 49830
rect 524432 45526 524552 45554
rect 523224 39568 523276 39574
rect 523224 39510 523276 39516
rect 523040 38072 523092 38078
rect 523040 38014 523092 38020
rect 524420 33788 524472 33794
rect 524420 33730 524472 33736
rect 523040 32496 523092 32502
rect 523040 32438 523092 32444
rect 521764 16546 521884 16574
rect 520372 10328 520424 10334
rect 520372 10270 520424 10276
rect 521856 480 521884 16546
rect 523052 480 523080 32438
rect 523132 23044 523184 23050
rect 523132 22986 523184 22992
rect 523144 16574 523172 22986
rect 524432 16574 524460 33730
rect 524524 25702 524552 45526
rect 525800 33856 525852 33862
rect 525800 33798 525852 33804
rect 524512 25696 524564 25702
rect 524512 25638 524564 25644
rect 523144 16546 523816 16574
rect 524432 16546 525472 16574
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 520710 -960 520822 326
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 523788 354 523816 16546
rect 525444 480 525472 16546
rect 525812 6914 525840 33798
rect 525904 10402 525932 50215
rect 526074 49736 526130 49745
rect 526074 49671 526130 49680
rect 526088 20058 526116 49671
rect 527192 45554 527220 50238
rect 528558 49736 528614 49745
rect 528558 49671 528614 49680
rect 527192 45526 527312 45554
rect 527180 29776 527232 29782
rect 527180 29718 527232 29724
rect 526076 20052 526128 20058
rect 526076 19994 526128 20000
rect 525892 10396 525944 10402
rect 525892 10338 525944 10344
rect 527192 6914 527220 29718
rect 527284 10470 527312 45526
rect 528572 44946 528600 49671
rect 528560 44940 528612 44946
rect 528560 44882 528612 44888
rect 529940 35284 529992 35290
rect 529940 35226 529992 35232
rect 528560 15904 528612 15910
rect 528560 15846 528612 15852
rect 527272 10464 527324 10470
rect 527272 10406 527324 10412
rect 525812 6886 526208 6914
rect 527192 6886 527864 6914
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526180 354 526208 6886
rect 527836 480 527864 6886
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 15846
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 35226
rect 530044 10538 530072 50487
rect 532698 50416 532754 50425
rect 532698 50351 532754 50360
rect 536838 50416 536894 50425
rect 537482 50416 537538 50425
rect 536894 50374 536972 50402
rect 536838 50351 536894 50360
rect 531318 50280 531374 50289
rect 531318 50215 531374 50224
rect 530214 49736 530270 49745
rect 530214 49671 530270 49680
rect 530228 42294 530256 49671
rect 530216 42288 530268 42294
rect 530216 42230 530268 42236
rect 531332 32638 531360 50215
rect 532712 43654 532740 50351
rect 534170 50280 534226 50289
rect 534170 50215 534226 50224
rect 532882 49872 532938 49881
rect 532882 49807 532938 49816
rect 532700 43648 532752 43654
rect 532700 43590 532752 43596
rect 532700 36644 532752 36650
rect 532700 36586 532752 36592
rect 531320 32632 531372 32638
rect 531320 32574 531372 32580
rect 531320 31204 531372 31210
rect 531320 31146 531372 31152
rect 530032 10532 530084 10538
rect 530032 10474 530084 10480
rect 531332 480 531360 31146
rect 532712 16574 532740 36586
rect 532896 22846 532924 49807
rect 534080 27124 534132 27130
rect 534080 27066 534132 27072
rect 532884 22840 532936 22846
rect 532884 22782 532936 22788
rect 532712 16546 533752 16574
rect 532516 8968 532568 8974
rect 532516 8910 532568 8916
rect 532528 480 532556 8910
rect 533724 480 533752 16546
rect 534092 6914 534120 27066
rect 534184 10606 534212 50215
rect 535458 49736 535514 49745
rect 535458 49671 535514 49680
rect 534172 10600 534224 10606
rect 534172 10542 534224 10548
rect 534092 6886 534488 6914
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534460 354 534488 6886
rect 535472 3466 535500 49671
rect 536944 10674 536972 50374
rect 537482 50351 537538 50360
rect 539690 50416 539746 50425
rect 542358 50416 542414 50425
rect 539746 50374 539824 50402
rect 539690 50351 539746 50360
rect 537496 50153 537524 50351
rect 538310 50280 538366 50289
rect 538310 50215 538366 50224
rect 537482 50144 537538 50153
rect 537482 50079 537538 50088
rect 537114 49872 537170 49881
rect 537114 49807 537170 49816
rect 536932 10668 536984 10674
rect 536932 10610 536984 10616
rect 535460 3460 535512 3466
rect 535460 3402 535512 3408
rect 537128 3369 537156 49807
rect 538220 38140 538272 38146
rect 538220 38082 538272 38088
rect 537208 4888 537260 4894
rect 537208 4830 537260 4836
rect 537114 3360 537170 3369
rect 537114 3295 537170 3304
rect 536104 3188 536156 3194
rect 536104 3130 536156 3136
rect 536116 480 536144 3130
rect 537220 480 537248 4830
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 38082
rect 538324 3534 538352 50215
rect 539690 49736 539746 49745
rect 539690 49671 539746 49680
rect 539704 3670 539732 49671
rect 539796 45554 539824 50374
rect 542358 50351 542414 50360
rect 540702 49872 540758 49881
rect 540758 49830 541112 49858
rect 540702 49807 540758 49816
rect 540980 46368 541032 46374
rect 540980 46310 541032 46316
rect 539796 45526 539916 45554
rect 539692 3664 539744 3670
rect 539692 3606 539744 3612
rect 539888 3602 539916 45526
rect 540796 4820 540848 4826
rect 540796 4762 540848 4768
rect 539876 3596 539928 3602
rect 539876 3538 539928 3544
rect 538312 3528 538364 3534
rect 538312 3470 538364 3476
rect 539600 3460 539652 3466
rect 539600 3402 539652 3408
rect 539612 480 539640 3402
rect 540808 480 540836 4762
rect 540992 3482 541020 46310
rect 541084 3738 541112 49830
rect 542372 3806 542400 50351
rect 543830 49872 543886 49881
rect 543830 49807 543886 49816
rect 542542 49736 542598 49745
rect 542542 49671 542598 49680
rect 542556 9042 542584 49671
rect 543740 46300 543792 46306
rect 543740 46242 543792 46248
rect 542544 9036 542596 9042
rect 542544 8978 542596 8984
rect 542360 3800 542412 3806
rect 542360 3742 542412 3748
rect 541072 3732 541124 3738
rect 541072 3674 541124 3680
rect 543188 3528 543240 3534
rect 540992 3454 542032 3482
rect 543188 3470 543240 3476
rect 543752 3482 543780 46242
rect 543844 3874 543872 49807
rect 545120 32700 545172 32706
rect 545120 32642 545172 32648
rect 543832 3868 543884 3874
rect 543832 3810 543884 3816
rect 545132 3482 545160 32642
rect 545224 3942 545252 50623
rect 546774 50552 546830 50561
rect 546774 50487 546830 50496
rect 546590 49736 546646 49745
rect 546590 49671 546646 49680
rect 546604 4078 546632 49671
rect 546592 4072 546644 4078
rect 546592 4014 546644 4020
rect 546788 4010 546816 50487
rect 549534 50416 549590 50425
rect 549534 50351 549590 50360
rect 553490 50416 553546 50425
rect 553490 50351 553546 50360
rect 556158 50416 556214 50425
rect 556158 50351 556214 50360
rect 565910 50416 565966 50425
rect 565910 50351 565966 50360
rect 570234 50416 570290 50425
rect 570234 50351 570290 50360
rect 573086 50416 573142 50425
rect 573086 50351 573142 50360
rect 575570 50416 575626 50425
rect 575570 50351 575626 50360
rect 580262 50416 580318 50425
rect 580262 50351 580318 50360
rect 549350 50280 549406 50289
rect 549350 50215 549406 50224
rect 548062 49872 548118 49881
rect 548062 49807 548118 49816
rect 547880 38004 547932 38010
rect 547880 37946 547932 37952
rect 546776 4004 546828 4010
rect 546776 3946 546828 3952
rect 545212 3936 545264 3942
rect 545212 3878 545264 3884
rect 546684 3596 546736 3602
rect 546684 3538 546736 3544
rect 542004 480 542032 3454
rect 543200 480 543228 3470
rect 543752 3454 544424 3482
rect 545132 3454 545528 3482
rect 544396 480 544424 3454
rect 545500 480 545528 3454
rect 546696 480 546724 3538
rect 547892 480 547920 37946
rect 548076 4146 548104 49807
rect 549076 8084 549128 8090
rect 549076 8026 549128 8032
rect 548064 4140 548116 4146
rect 548064 4082 548116 4088
rect 549088 480 549116 8026
rect 549364 3330 549392 50215
rect 549548 3398 549576 50351
rect 552018 50280 552074 50289
rect 552018 50215 552074 50224
rect 550730 49736 550786 49745
rect 550730 49671 550786 49680
rect 550640 39432 550692 39438
rect 550640 39374 550692 39380
rect 550272 3664 550324 3670
rect 550272 3606 550324 3612
rect 549536 3392 549588 3398
rect 549536 3334 549588 3340
rect 549352 3324 549404 3330
rect 549352 3266 549404 3272
rect 550284 480 550312 3606
rect 550652 490 550680 39374
rect 550744 3262 550772 49671
rect 552032 4962 552060 50215
rect 552664 8016 552716 8022
rect 552664 7958 552716 7964
rect 552020 4956 552072 4962
rect 552020 4898 552072 4904
rect 550732 3256 550784 3262
rect 550732 3198 550784 3204
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 550652 462 551048 490
rect 552676 480 552704 7958
rect 553504 5098 553532 50351
rect 554870 50280 554926 50289
rect 554870 50215 554926 50224
rect 553674 49872 553730 49881
rect 553674 49807 553730 49816
rect 553492 5092 553544 5098
rect 553492 5034 553544 5040
rect 553688 5030 553716 49807
rect 554780 40792 554832 40798
rect 554780 40734 554832 40740
rect 553676 5024 553728 5030
rect 553676 4966 553728 4972
rect 553768 3732 553820 3738
rect 553768 3674 553820 3680
rect 553780 480 553808 3674
rect 551020 354 551048 462
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 40734
rect 554884 5166 554912 50215
rect 556172 45554 556200 50351
rect 557538 50280 557594 50289
rect 557538 50215 557594 50224
rect 559102 50280 559158 50289
rect 559102 50215 559158 50224
rect 561770 50280 561826 50289
rect 561770 50215 561826 50224
rect 564530 50280 564586 50289
rect 564530 50215 564586 50224
rect 556250 49872 556306 49881
rect 556306 49830 556384 49858
rect 556250 49807 556306 49816
rect 556356 45554 556384 49830
rect 557552 45554 557580 50215
rect 557630 50144 557686 50153
rect 557630 50079 557686 50088
rect 557644 47598 557672 50079
rect 557632 47592 557684 47598
rect 557632 47534 557684 47540
rect 556172 45526 556292 45554
rect 556356 45526 556476 45554
rect 557552 45526 557672 45554
rect 556160 7948 556212 7954
rect 556160 7890 556212 7896
rect 554872 5160 554924 5166
rect 554872 5102 554924 5108
rect 556172 480 556200 7890
rect 556264 5302 556292 45526
rect 556252 5296 556304 5302
rect 556252 5238 556304 5244
rect 556448 5234 556476 45526
rect 557540 44872 557592 44878
rect 557540 44814 557592 44820
rect 556436 5228 556488 5234
rect 556436 5170 556488 5176
rect 557356 3800 557408 3806
rect 557356 3742 557408 3748
rect 557368 480 557396 3742
rect 557552 3482 557580 44814
rect 557644 5370 557672 45526
rect 559116 14482 559144 50215
rect 560390 49872 560446 49881
rect 560390 49807 560446 49816
rect 560298 49736 560354 49745
rect 560298 49671 560354 49680
rect 559104 14476 559156 14482
rect 559104 14418 559156 14424
rect 559288 13388 559340 13394
rect 559288 13330 559340 13336
rect 557632 5364 557684 5370
rect 557632 5306 557684 5312
rect 557552 3454 558592 3482
rect 558564 480 558592 3454
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559300 354 559328 13330
rect 560312 6186 560340 49671
rect 560404 49026 560432 49807
rect 560392 49020 560444 49026
rect 560392 48962 560444 48968
rect 561680 43512 561732 43518
rect 561680 43454 561732 43460
rect 561692 6914 561720 43454
rect 561784 11762 561812 50215
rect 563242 49736 563298 49745
rect 563242 49671 563298 49680
rect 563256 33794 563284 49671
rect 564440 42152 564492 42158
rect 564440 42094 564492 42100
rect 563244 33788 563296 33794
rect 563244 33730 563296 33736
rect 561772 11756 561824 11762
rect 561772 11698 561824 11704
rect 563244 7880 563296 7886
rect 563244 7822 563296 7828
rect 561692 6886 562088 6914
rect 560300 6180 560352 6186
rect 560300 6122 560352 6128
rect 560852 3868 560904 3874
rect 560852 3810 560904 3816
rect 560864 480 560892 3810
rect 562060 480 562088 6886
rect 563256 480 563284 7822
rect 564452 6914 564480 42094
rect 564544 15910 564572 50215
rect 564532 15904 564584 15910
rect 564532 15846 564584 15852
rect 564452 6886 565216 6914
rect 564440 3936 564492 3942
rect 564440 3878 564492 3884
rect 564452 480 564480 3878
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 559718 -960 559830 326
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565188 354 565216 6886
rect 565924 3194 565952 50351
rect 567106 50280 567162 50289
rect 567162 50238 567240 50266
rect 567106 50215 567162 50224
rect 566002 49872 566058 49881
rect 566002 49807 566058 49816
rect 566016 45554 566044 49807
rect 566016 45526 566136 45554
rect 566108 8974 566136 45526
rect 566096 8968 566148 8974
rect 566096 8910 566148 8916
rect 566832 7812 566884 7818
rect 566832 7754 566884 7760
rect 565912 3188 565964 3194
rect 565912 3130 565964 3136
rect 566844 480 566872 7754
rect 567212 3466 567240 50238
rect 570050 49872 570106 49881
rect 570050 49807 570106 49816
rect 568670 49736 568726 49745
rect 568670 49671 568726 49680
rect 568580 18692 568632 18698
rect 568580 18634 568632 18640
rect 568592 6914 568620 18634
rect 568684 16574 568712 49671
rect 568684 16546 568804 16574
rect 568592 6886 568712 6914
rect 567200 3460 567252 3466
rect 567200 3402 567252 3408
rect 568028 3392 568080 3398
rect 568028 3334 568080 3340
rect 568040 480 568068 3334
rect 565606 354 565718 480
rect 565188 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 568684 354 568712 6886
rect 568776 3534 568804 16546
rect 570064 3670 570092 49807
rect 570052 3664 570104 3670
rect 570052 3606 570104 3612
rect 570248 3602 570276 50351
rect 571338 50280 571394 50289
rect 571338 50215 571394 50224
rect 570328 7744 570380 7750
rect 570328 7686 570380 7692
rect 570236 3596 570288 3602
rect 570236 3538 570288 3544
rect 568764 3528 568816 3534
rect 568764 3470 568816 3476
rect 570340 480 570368 7686
rect 571352 3738 571380 50215
rect 572810 49872 572866 49881
rect 572810 49807 572866 49816
rect 572824 45554 572852 49807
rect 572824 45526 572944 45554
rect 572720 19984 572772 19990
rect 572720 19926 572772 19932
rect 571340 3732 571392 3738
rect 571340 3674 571392 3680
rect 571524 3052 571576 3058
rect 571524 2994 571576 3000
rect 571536 480 571564 2994
rect 572732 480 572760 19926
rect 572916 3806 572944 45526
rect 573100 3874 573128 50351
rect 574098 50280 574154 50289
rect 574098 50215 574154 50224
rect 573916 7676 573968 7682
rect 573916 7618 573968 7624
rect 573088 3868 573140 3874
rect 573088 3810 573140 3816
rect 572904 3800 572956 3806
rect 572904 3742 572956 3748
rect 573928 480 573956 7618
rect 574112 3942 574140 50215
rect 574744 21412 574796 21418
rect 574744 21354 574796 21360
rect 574100 3936 574152 3942
rect 574100 3878 574152 3884
rect 574756 3466 574784 21354
rect 575112 3528 575164 3534
rect 575112 3470 575164 3476
rect 574744 3460 574796 3466
rect 574744 3402 574796 3408
rect 575124 480 575152 3470
rect 575584 3058 575612 50351
rect 576950 50280 577006 50289
rect 576950 50215 577006 50224
rect 575754 49872 575810 49881
rect 575754 49807 575810 49816
rect 575768 3398 575796 49807
rect 576964 3534 576992 50215
rect 578238 49736 578294 49745
rect 578238 49671 578294 49680
rect 578252 16574 578280 49671
rect 578252 16546 578648 16574
rect 577412 7608 577464 7614
rect 577412 7550 577464 7556
rect 576952 3528 577004 3534
rect 576952 3470 577004 3476
rect 576308 3460 576360 3466
rect 576308 3402 576360 3408
rect 575756 3392 575808 3398
rect 575756 3334 575808 3340
rect 575572 3052 575624 3058
rect 575572 2994 575624 3000
rect 576320 480 576348 3402
rect 577424 480 577452 7550
rect 578620 480 578648 16546
rect 580276 3330 580304 50351
rect 582286 50280 582342 50289
rect 582342 50238 582420 50266
rect 582286 50215 582342 50224
rect 582392 11762 582420 50238
rect 582470 49736 582526 49745
rect 582470 49671 582526 49680
rect 582380 11756 582432 11762
rect 582380 11698 582432 11704
rect 582484 6914 582512 49671
rect 583392 11756 583444 11762
rect 583392 11698 583444 11704
rect 582392 6886 582512 6914
rect 582392 3482 582420 6886
rect 582208 3454 582420 3482
rect 580264 3324 580316 3330
rect 580264 3266 580316 3272
rect 581000 3324 581052 3330
rect 581000 3266 581052 3272
rect 581012 480 581040 3266
rect 582208 480 582236 3454
rect 583404 480 583432 11698
rect 569102 354 569214 480
rect 568684 326 569214 354
rect 569102 -960 569214 326
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 181626 50768 181682 50824
rect 449162 50768 449218 50824
rect 162122 50632 162178 50688
rect 99378 50224 99434 50280
rect 97998 49816 98054 49872
rect 98642 49680 98698 49736
rect 6458 3304 6514 3360
rect 178682 50632 178738 50688
rect 180706 50632 180762 50688
rect 181442 50632 181498 50688
rect 102782 50496 102838 50552
rect 109038 50496 109094 50552
rect 113822 50496 113878 50552
rect 133142 50496 133198 50552
rect 142802 50496 142858 50552
rect 152462 50496 152518 50552
rect 160742 50496 160798 50552
rect 101586 50360 101642 50416
rect 101402 49544 101458 49600
rect 104162 49816 104218 49872
rect 105910 50360 105966 50416
rect 108118 50360 108174 50416
rect 108302 50360 108358 50416
rect 106922 50224 106978 50280
rect 105726 49680 105782 49736
rect 108118 50088 108174 50144
rect 108486 49680 108542 49736
rect 112442 50360 112498 50416
rect 111062 49816 111118 49872
rect 112626 49680 112682 49736
rect 119342 50360 119398 50416
rect 123482 50360 123538 50416
rect 131762 50360 131818 50416
rect 115202 49816 115258 49872
rect 115386 49680 115442 49736
rect 116674 50224 116730 50280
rect 116674 49952 116730 50008
rect 118606 49816 118662 49872
rect 116674 49680 116730 49736
rect 117962 49680 118018 49736
rect 122470 50224 122526 50280
rect 120722 49816 120778 49872
rect 122102 49680 122158 49736
rect 126426 50224 126482 50280
rect 125046 49816 125102 49872
rect 124862 49680 124918 49736
rect 126518 49952 126574 50008
rect 127622 49816 127678 49872
rect 126518 49680 126574 49736
rect 129002 49680 129058 49736
rect 129278 50224 129334 50280
rect 130382 49544 130438 49600
rect 131946 49680 132002 49736
rect 138662 50360 138718 50416
rect 141606 50360 141662 50416
rect 136086 50224 136142 50280
rect 134706 49816 134762 49872
rect 134522 49680 134578 49736
rect 136178 49952 136234 50008
rect 137282 49816 137338 49872
rect 136178 49680 136234 49736
rect 140042 50224 140098 50280
rect 138846 49680 138902 49736
rect 141422 49680 141478 49736
rect 148506 50360 148562 50416
rect 151082 50360 151138 50416
rect 145838 50224 145894 50280
rect 148322 50224 148378 50280
rect 144182 49816 144238 49872
rect 144366 49680 144422 49736
rect 145930 49952 145986 50008
rect 145930 49680 145986 49736
rect 146942 49680 146998 49736
rect 150530 49816 150586 49872
rect 149794 49680 149850 49736
rect 151726 50224 151782 50280
rect 151726 49680 151782 49736
rect 153842 49816 153898 49872
rect 155590 50360 155646 50416
rect 157798 50360 157854 50416
rect 156602 50224 156658 50280
rect 155406 49680 155462 49736
rect 159454 50224 159510 50280
rect 157798 50088 157854 50144
rect 158166 49816 158222 49872
rect 157982 49680 158038 49736
rect 159546 49952 159602 50008
rect 159546 49680 159602 49736
rect 160926 49680 160982 49736
rect 170402 50496 170458 50552
rect 163502 49816 163558 49872
rect 165342 50360 165398 50416
rect 167642 50360 167698 50416
rect 166262 50224 166318 50280
rect 167642 50224 167698 50280
rect 165066 49680 165122 49736
rect 167826 50360 167882 50416
rect 167734 50088 167790 50144
rect 169022 49816 169078 49872
rect 174726 50360 174782 50416
rect 177118 50360 177174 50416
rect 177486 50360 177542 50416
rect 173162 50224 173218 50280
rect 172150 49816 172206 49872
rect 171782 49680 171838 49736
rect 173254 49952 173310 50008
rect 173254 49680 173310 49736
rect 174542 49680 174598 49736
rect 176014 50224 176070 50280
rect 177118 50088 177174 50144
rect 177302 49680 177358 49736
rect 180062 50496 180118 50552
rect 180706 50360 180762 50416
rect 200762 50632 200818 50688
rect 278686 50632 278742 50688
rect 288346 50632 288402 50688
rect 363050 50632 363106 50688
rect 410522 50632 410578 50688
rect 421746 50632 421802 50688
rect 424506 50632 424562 50688
rect 431314 50632 431370 50688
rect 434626 50632 434682 50688
rect 185582 50496 185638 50552
rect 195242 50496 195298 50552
rect 199382 50496 199438 50552
rect 184846 50360 184902 50416
rect 182822 49816 182878 49872
rect 184202 49680 184258 49736
rect 188526 50360 188582 50416
rect 190918 50360 190974 50416
rect 193862 50360 193918 50416
rect 186962 49680 187018 49736
rect 188342 49544 188398 49600
rect 189722 50224 189778 50280
rect 190918 50088 190974 50144
rect 191102 49816 191158 49872
rect 191286 49680 191342 49736
rect 192574 50224 192630 50280
rect 192574 49952 192630 50008
rect 192574 49680 192630 49736
rect 194046 49680 194102 49736
rect 196622 49680 196678 49736
rect 198462 50360 198518 50416
rect 198186 49544 198242 49600
rect 199382 3304 199438 3360
rect 214562 50496 214618 50552
rect 221462 50496 221518 50552
rect 225602 50496 225658 50552
rect 227718 50496 227774 50552
rect 250994 50496 251050 50552
rect 259366 50496 259422 50552
rect 269026 50496 269082 50552
rect 277306 50496 277362 50552
rect 211802 50360 211858 50416
rect 203522 50224 203578 50280
rect 206282 50224 206338 50280
rect 209134 50224 209190 50280
rect 202142 49816 202198 49872
rect 200946 49680 201002 49736
rect 204258 49952 204314 50008
rect 203890 49816 203946 49872
rect 204902 49816 204958 49872
rect 205086 49680 205142 49736
rect 208122 49816 208178 49872
rect 207662 49544 207718 49600
rect 211066 49816 211122 49872
rect 210606 49680 210662 49736
rect 213182 49680 213238 49736
rect 218702 50360 218758 50416
rect 214930 50224 214986 50280
rect 217322 49816 217378 49872
rect 215942 49680 215998 49736
rect 217506 49544 217562 49600
rect 220082 49680 220138 49736
rect 221830 50224 221886 50280
rect 222842 49816 222898 49872
rect 224682 50224 224738 50280
rect 224406 49680 224462 49736
rect 226982 49816 227038 49872
rect 227166 49680 227222 49736
rect 233146 50360 233202 50416
rect 234434 50360 234490 50416
rect 249706 50360 249762 50416
rect 231490 50224 231546 50280
rect 230386 49816 230442 49872
rect 231674 49680 231730 49736
rect 235906 50224 235962 50280
rect 238482 50224 238538 50280
rect 241426 50224 241482 50280
rect 248050 50224 248106 50280
rect 234526 49816 234582 49872
rect 237286 49680 237342 49736
rect 241242 49816 241298 49872
rect 238666 49680 238722 49736
rect 242714 49952 242770 50008
rect 246762 49952 246818 50008
rect 242806 49680 242862 49736
rect 245566 49680 245622 49736
rect 246946 49816 247002 49872
rect 246854 49544 246910 49600
rect 248234 49680 248290 49736
rect 250810 49816 250866 49872
rect 253754 50360 253810 50416
rect 253570 50224 253626 50280
rect 252466 49680 252522 49736
rect 257894 50224 257950 50280
rect 257802 49836 257858 49872
rect 257802 49816 257804 49836
rect 257804 49816 257856 49836
rect 257856 49816 257858 49836
rect 255226 49680 255282 49736
rect 257802 49680 257858 49736
rect 266266 50360 266322 50416
rect 262126 50224 262182 50280
rect 264794 50224 264850 50280
rect 260654 49816 260710 49872
rect 260470 49680 260526 49736
rect 262678 49952 262734 50008
rect 262310 49816 262366 49872
rect 263506 49816 263562 49872
rect 264610 49680 264666 49736
rect 267554 49816 267610 49872
rect 267370 49680 267426 49736
rect 271786 50224 271842 50280
rect 274362 50224 274418 50280
rect 270406 49816 270462 49872
rect 270222 49680 270278 49736
rect 272430 49952 272486 50008
rect 272062 49816 272118 49872
rect 273166 49816 273222 49872
rect 274546 49680 274602 49736
rect 277214 49680 277270 49736
rect 275926 49544 275982 49600
rect 286690 50496 286746 50552
rect 281170 50360 281226 50416
rect 285586 50360 285642 50416
rect 282734 49816 282790 49872
rect 281354 49680 281410 49736
rect 283102 49816 283158 49872
rect 284022 49680 284078 49736
rect 286322 49816 286378 49872
rect 286966 49816 287022 49872
rect 292486 50496 292542 50552
rect 315946 50496 316002 50552
rect 330482 50496 330538 50552
rect 336002 50496 336058 50552
rect 343638 50496 343694 50552
rect 354678 50496 354734 50552
rect 289726 49680 289782 49736
rect 290922 50360 290978 50416
rect 291014 49680 291070 49736
rect 297730 50360 297786 50416
rect 304814 50360 304870 50416
rect 307482 50360 307538 50416
rect 314290 50360 314346 50416
rect 295246 50224 295302 50280
rect 293590 49816 293646 49872
rect 293774 49680 293830 49736
rect 296626 49544 296682 49600
rect 297914 50224 297970 50280
rect 300674 50224 300730 50280
rect 299386 49816 299442 49872
rect 300490 49680 300546 49736
rect 303526 50224 303582 50280
rect 303526 49680 303582 49736
rect 304906 49816 304962 49872
rect 306286 49680 306342 49736
rect 307666 50224 307722 50280
rect 310426 50224 310482 50280
rect 311806 50224 311862 50280
rect 310242 49816 310298 49872
rect 311714 49952 311770 50008
rect 313186 49680 313242 49736
rect 314474 49544 314530 49600
rect 324134 50360 324190 50416
rect 326158 50360 326214 50416
rect 327722 50360 327778 50416
rect 318706 50224 318762 50280
rect 321466 50224 321522 50280
rect 318154 49952 318210 50008
rect 317142 49816 317198 49872
rect 317326 49680 317382 49736
rect 318154 49680 318210 49736
rect 321098 49952 321154 50008
rect 320086 49816 320142 49872
rect 319994 49680 320050 49736
rect 321098 49680 321154 49736
rect 322846 49680 322902 49736
rect 323950 49544 324006 49600
rect 324962 50224 325018 50280
rect 326158 50088 326214 50144
rect 326342 49816 326398 49872
rect 326526 49680 326582 49736
rect 329194 49816 329250 49872
rect 331862 50224 331918 50280
rect 330666 49680 330722 49736
rect 333702 50360 333758 50416
rect 334714 50224 334770 50280
rect 333426 49680 333482 49736
rect 336186 49680 336242 49736
rect 342258 49680 342314 49736
rect 345202 50360 345258 50416
rect 345018 49952 345074 50008
rect 345110 49680 345166 49736
rect 346490 50224 346546 50280
rect 351918 50224 351974 50280
rect 346398 49816 346454 49872
rect 351826 49836 351882 49872
rect 351826 49816 351828 49836
rect 351828 49816 351880 49836
rect 351880 49816 351882 49836
rect 347962 49680 348018 49736
rect 348146 49680 348202 49736
rect 352194 49680 352250 49736
rect 356058 50360 356114 50416
rect 354862 49816 354918 49872
rect 357714 50224 357770 50280
rect 360198 50224 360254 50280
rect 357530 49680 357586 49736
rect 358910 49816 358966 49872
rect 360658 49952 360714 50008
rect 361578 49816 361634 49872
rect 360658 49680 360714 49736
rect 361578 49680 361634 49736
rect 364614 50496 364670 50552
rect 382278 50496 382334 50552
rect 398930 50496 398986 50552
rect 364430 49816 364486 49872
rect 365718 50360 365774 50416
rect 374366 50360 374422 50416
rect 367282 50224 367338 50280
rect 369950 50224 370006 50280
rect 367098 49680 367154 49736
rect 368754 50020 368810 50076
rect 368478 49816 368534 49872
rect 369858 49816 369914 49872
rect 371422 49680 371478 49736
rect 374182 49680 374238 49736
rect 376850 50224 376906 50280
rect 379518 50224 379574 50280
rect 375194 49816 375250 49872
rect 375378 49680 375434 49736
rect 378322 49680 378378 49736
rect 380070 49952 380126 50008
rect 380898 49816 380954 49872
rect 380070 49680 380126 49736
rect 381082 49680 381138 49736
rect 383750 50360 383806 50416
rect 385038 50360 385094 50416
rect 387982 50360 388038 50416
rect 393410 50360 393466 50416
rect 395066 50360 395122 50416
rect 383934 49816 383990 49872
rect 386510 50224 386566 50280
rect 387798 49952 387854 50008
rect 389178 50224 389234 50280
rect 388166 49816 388222 49872
rect 391938 49816 391994 49872
rect 390742 49680 390798 49736
rect 394698 49816 394754 49872
rect 394698 49680 394754 49736
rect 396170 50224 396226 50280
rect 397458 49680 397514 49736
rect 400494 50360 400550 50416
rect 400310 49680 400366 49736
rect 403070 50224 403126 50280
rect 404542 50224 404598 50280
rect 407762 50224 407818 50280
rect 402978 49816 403034 49872
rect 401690 49680 401746 49736
rect 407118 49816 407174 49872
rect 405830 49680 405886 49736
rect 409142 49816 409198 49872
rect 412086 50496 412142 50552
rect 411902 49680 411958 49736
rect 416686 50360 416742 50416
rect 420182 50360 420238 50416
rect 413282 50224 413338 50280
rect 412546 49952 412602 50008
rect 412546 49680 412602 49736
rect 414846 49816 414902 49872
rect 414662 49680 414718 49736
rect 417422 50224 417478 50280
rect 418802 49816 418858 49872
rect 417606 49680 417662 49736
rect 422942 50224 422998 50280
rect 421746 50088 421802 50144
rect 421562 49816 421618 49872
rect 421746 49680 421802 49736
rect 424322 49544 424378 49600
rect 427082 50496 427138 50552
rect 425702 49680 425758 49736
rect 428462 50360 428518 50416
rect 429750 50224 429806 50280
rect 429658 49952 429714 50008
rect 428646 49680 428702 49736
rect 429658 49680 429714 49736
rect 432602 50360 432658 50416
rect 431314 50088 431370 50144
rect 431406 49816 431462 49872
rect 431222 49680 431278 49736
rect 429658 3304 429714 3360
rect 433982 50224 434038 50280
rect 441066 50360 441122 50416
rect 445666 50360 445722 50416
rect 438122 50224 438178 50280
rect 436466 49952 436522 50008
rect 435362 49680 435418 49736
rect 436558 49816 436614 49872
rect 440422 49816 440478 49872
rect 439502 49680 439558 49736
rect 442262 49816 442318 49872
rect 445022 49680 445078 49736
rect 443734 49544 443790 49600
rect 446310 50224 446366 50280
rect 446218 49952 446274 50008
rect 446218 49680 446274 49736
rect 447966 49816 448022 49872
rect 447782 49680 447838 49736
rect 450542 50632 450598 50688
rect 461030 50632 461086 50688
rect 498290 50632 498346 50688
rect 545210 50632 545266 50688
rect 453302 50496 453358 50552
rect 451922 49816 451978 49872
rect 450726 49680 450782 49736
rect 454682 50360 454738 50416
rect 454406 49952 454462 50008
rect 454038 49680 454094 49736
rect 456982 50224 457038 50280
rect 455510 49816 455566 49872
rect 458270 49680 458326 49736
rect 459558 49680 459614 49736
rect 462410 50496 462466 50552
rect 491298 50496 491354 50552
rect 461214 49816 461270 49872
rect 463790 50360 463846 50416
rect 466550 50360 466606 50416
rect 470690 50360 470746 50416
rect 470966 50360 471022 50416
rect 473358 50360 473414 50416
rect 476486 50360 476542 50416
rect 478878 50360 478934 50416
rect 483294 50360 483350 50416
rect 488538 50360 488594 50416
rect 465170 50224 465226 50280
rect 463974 49680 464030 49736
rect 467654 50224 467710 50280
rect 466734 49816 466790 49872
rect 469218 49680 469274 49736
rect 470598 49680 470654 49736
rect 471978 50224 472034 50280
rect 470966 50088 471022 50144
rect 470874 49816 470930 49872
rect 474462 49680 474518 49736
rect 476302 49680 476358 49736
rect 477498 49680 477554 49736
rect 480350 50224 480406 50280
rect 480258 49952 480314 50008
rect 480350 49816 480406 49872
rect 480258 49680 480314 49736
rect 481362 49680 481418 49736
rect 483110 49680 483166 49736
rect 484306 50224 484362 50280
rect 484582 49952 484638 50008
rect 487434 49816 487490 49872
rect 485778 49680 485834 49736
rect 490194 49816 490250 49872
rect 490010 49680 490066 49736
rect 492862 50224 492918 50280
rect 495438 50224 495494 50280
rect 492678 49680 492734 49736
rect 494150 49680 494206 49736
rect 495898 49952 495954 50008
rect 496910 49816 496966 49872
rect 495898 49680 495954 49736
rect 497094 49680 497150 49736
rect 499670 50496 499726 50552
rect 501050 50496 501106 50552
rect 507950 50496 508006 50552
rect 514850 50496 514906 50552
rect 530030 50496 530086 50552
rect 499854 49816 499910 49872
rect 503718 50360 503774 50416
rect 502338 49680 502394 49736
rect 505098 50224 505154 50280
rect 503902 49680 503958 49736
rect 505650 49952 505706 50008
rect 506570 49816 506626 49872
rect 505650 49680 505706 49736
rect 506754 49680 506810 49736
rect 509514 50360 509570 50416
rect 509330 49680 509386 49736
rect 512090 50224 512146 50280
rect 510710 49680 510766 49736
rect 512458 49952 512514 50008
rect 513654 49816 513710 49872
rect 512458 49680 512514 49736
rect 513470 49680 513526 49736
rect 516138 50360 516194 50416
rect 518990 50360 519046 50416
rect 517702 49952 517758 50008
rect 517518 49816 517574 49872
rect 516322 49680 516378 49736
rect 520278 50224 520334 50280
rect 519174 49680 519230 49736
rect 523038 50224 523094 50280
rect 525890 50224 525946 50280
rect 527086 50224 527142 50280
rect 524142 49816 524198 49872
rect 523222 49680 523278 49736
rect 526074 49680 526130 49736
rect 528558 49680 528614 49736
rect 532698 50360 532754 50416
rect 536838 50360 536894 50416
rect 531318 50224 531374 50280
rect 530214 49680 530270 49736
rect 534170 50224 534226 50280
rect 532882 49816 532938 49872
rect 535458 49680 535514 49736
rect 537482 50360 537538 50416
rect 539690 50360 539746 50416
rect 538310 50224 538366 50280
rect 537482 50088 537538 50144
rect 537114 49816 537170 49872
rect 537114 3304 537170 3360
rect 539690 49680 539746 49736
rect 542358 50360 542414 50416
rect 540702 49816 540758 49872
rect 543830 49816 543886 49872
rect 542542 49680 542598 49736
rect 546774 50496 546830 50552
rect 546590 49680 546646 49736
rect 549534 50360 549590 50416
rect 553490 50360 553546 50416
rect 556158 50360 556214 50416
rect 565910 50360 565966 50416
rect 570234 50360 570290 50416
rect 573086 50360 573142 50416
rect 575570 50360 575626 50416
rect 580262 50360 580318 50416
rect 549350 50224 549406 50280
rect 548062 49816 548118 49872
rect 552018 50224 552074 50280
rect 550730 49680 550786 49736
rect 554870 50224 554926 50280
rect 553674 49816 553730 49872
rect 557538 50224 557594 50280
rect 559102 50224 559158 50280
rect 561770 50224 561826 50280
rect 564530 50224 564586 50280
rect 556250 49816 556306 49872
rect 557630 50088 557686 50144
rect 560390 49816 560446 49872
rect 560298 49680 560354 49736
rect 563242 49680 563298 49736
rect 567106 50224 567162 50280
rect 566002 49816 566058 49872
rect 570050 49816 570106 49872
rect 568670 49680 568726 49736
rect 571338 50224 571394 50280
rect 572810 49816 572866 49872
rect 574098 50224 574154 50280
rect 576950 50224 577006 50280
rect 575754 49816 575810 49872
rect 578238 49680 578294 49736
rect 582286 50224 582342 50280
rect 582470 49680 582526 49736
<< metal3 >>
rect 583520 697084 584960 697324
rect -960 692052 480 692292
rect 583520 683756 584960 683996
rect 583520 670564 584960 670804
rect -960 668524 480 668764
rect 583520 657236 584960 657476
rect -960 645132 480 645372
rect 583520 643908 584960 644148
rect 583520 630716 584960 630956
rect -960 621604 480 621844
rect 583520 617388 584960 617628
rect 583520 604060 584960 604300
rect -960 598212 480 598452
rect 583520 590868 584960 591108
rect 583520 577540 584960 577780
rect -960 574684 480 574924
rect 583520 564212 584960 564452
rect -960 551292 480 551532
rect 583520 551020 584960 551260
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect 583520 511172 584960 511412
rect -960 504372 480 504612
rect 583520 497844 584960 498084
rect 583520 484516 584960 484756
rect -960 480844 480 481084
rect 583520 471324 584960 471564
rect 583520 457996 584960 458236
rect -960 457452 480 457692
rect 583520 444668 584960 444908
rect -960 433924 480 434164
rect 583520 431476 584960 431716
rect 583520 418148 584960 418388
rect -960 410532 480 410772
rect 583520 404820 584960 405060
rect 583520 391628 584960 391868
rect -960 387004 480 387244
rect 583520 378300 584960 378540
rect 583520 364972 584960 365212
rect -960 363612 480 363852
rect 583520 351780 584960 352020
rect -960 340084 480 340324
rect 583520 338452 584960 338692
rect 583520 325124 584960 325364
rect -960 316556 480 316796
rect 583520 311932 584960 312172
rect 583520 298604 584960 298844
rect -960 293164 480 293404
rect 583520 285276 584960 285516
rect 583520 272084 584960 272324
rect -960 269636 480 269876
rect 583520 258756 584960 258996
rect -960 246244 480 246484
rect 583520 245428 584960 245668
rect 583520 232236 584960 232476
rect -960 222716 480 222956
rect 583520 218908 584960 219148
rect 583520 205580 584960 205820
rect -960 199324 480 199564
rect 583520 192388 584960 192628
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 152404 480 152644
rect 583520 152540 584960 152780
rect 583520 139212 584960 139452
rect -960 128876 480 129116
rect 583520 125884 584960 126124
rect 583520 112692 584960 112932
rect -960 105484 480 105724
rect 583520 99364 584960 99604
rect 583520 86036 584960 86276
rect -960 81956 480 82196
rect 583520 72844 584960 73084
rect 583520 59516 584960 59756
rect -960 58564 480 58804
rect 181621 50826 181687 50829
rect 449157 50826 449223 50829
rect 181621 50824 184716 50826
rect 181621 50768 181626 50824
rect 181682 50768 184716 50824
rect 181621 50766 184716 50768
rect 181621 50763 181687 50766
rect 162117 50690 162183 50693
rect 178677 50690 178743 50693
rect 180701 50690 180767 50693
rect 162117 50688 165212 50690
rect 162117 50632 162122 50688
rect 162178 50632 165212 50688
rect 162117 50630 165212 50632
rect 162117 50627 162183 50630
rect 102777 50554 102843 50557
rect 109033 50554 109099 50557
rect 113817 50554 113883 50557
rect 133137 50554 133203 50557
rect 142797 50554 142863 50557
rect 152457 50554 152523 50557
rect 160737 50554 160803 50557
rect 102777 50552 105780 50554
rect 102777 50496 102782 50552
rect 102838 50496 105780 50552
rect 102777 50494 105780 50496
rect 102777 50491 102843 50494
rect 101581 50418 101647 50421
rect 101581 50416 104860 50418
rect 101581 50360 101586 50416
rect 101642 50360 104860 50416
rect 101581 50358 104860 50360
rect 101581 50355 101647 50358
rect 99373 50282 99439 50285
rect 99373 50280 102928 50282
rect 99373 50224 99378 50280
rect 99434 50224 102928 50280
rect 99373 50222 102928 50224
rect 99373 50219 99439 50222
rect 102868 50116 102928 50222
rect 104800 50116 104860 50358
rect 105720 50116 105780 50494
rect 109033 50552 112362 50554
rect 109033 50496 109038 50552
rect 109094 50496 112362 50552
rect 109033 50494 112362 50496
rect 109033 50491 109099 50494
rect 105905 50418 105971 50421
rect 108113 50418 108179 50421
rect 105905 50416 108179 50418
rect 105905 50360 105910 50416
rect 105966 50360 108118 50416
rect 108174 50360 108179 50416
rect 105905 50358 108179 50360
rect 105905 50355 105971 50358
rect 108113 50355 108179 50358
rect 108297 50418 108363 50421
rect 108297 50416 111668 50418
rect 108297 50360 108302 50416
rect 108358 50360 111668 50416
rect 108297 50358 111668 50360
rect 108297 50355 108363 50358
rect 106917 50282 106983 50285
rect 106917 50280 109736 50282
rect 106917 50224 106922 50280
rect 106978 50224 109736 50280
rect 106917 50222 109736 50224
rect 106917 50219 106983 50222
rect 108113 50146 108179 50149
rect 108113 50144 108694 50146
rect 108113 50088 108118 50144
rect 108174 50088 108694 50144
rect 109676 50116 109736 50222
rect 111608 50116 111668 50358
rect 112302 50282 112362 50494
rect 113817 50552 116544 50554
rect 113817 50496 113822 50552
rect 113878 50496 116544 50552
rect 113817 50494 116544 50496
rect 113817 50491 113883 50494
rect 112437 50418 112503 50421
rect 112437 50416 115532 50418
rect 112437 50360 112442 50416
rect 112498 50360 115532 50416
rect 112437 50358 115532 50360
rect 112437 50355 112503 50358
rect 112302 50222 112680 50282
rect 112620 50116 112680 50222
rect 115472 50116 115532 50358
rect 116484 50116 116544 50494
rect 133137 50552 135956 50554
rect 133137 50496 133142 50552
rect 133198 50496 135956 50552
rect 133137 50494 135956 50496
rect 133137 50491 133203 50494
rect 119337 50418 119403 50421
rect 123477 50418 123543 50421
rect 131757 50418 131823 50421
rect 119337 50416 122340 50418
rect 119337 50360 119342 50416
rect 119398 50360 122340 50416
rect 119337 50358 122340 50360
rect 119337 50355 119403 50358
rect 116669 50282 116735 50285
rect 116669 50280 119488 50282
rect 116669 50224 116674 50280
rect 116730 50224 119488 50280
rect 116669 50222 119488 50224
rect 116669 50219 116735 50222
rect 119428 50116 119488 50222
rect 120214 50222 121420 50282
rect 108113 50086 108694 50088
rect 108113 50083 108179 50086
rect 97993 49874 98059 49877
rect 100936 49874 100996 50048
rect 97993 49872 100996 49874
rect 97993 49816 97998 49872
rect 98054 49816 100996 49872
rect 97993 49814 100996 49816
rect 97993 49811 98059 49814
rect 98637 49738 98703 49741
rect 101856 49738 101916 50048
rect 103788 49738 103848 50048
rect 104157 49874 104223 49877
rect 106732 49874 106792 50048
rect 104157 49872 106792 49874
rect 104157 49816 104162 49872
rect 104218 49816 106792 49872
rect 104157 49814 106792 49816
rect 104157 49811 104223 49814
rect 98637 49736 101916 49738
rect 98637 49680 98642 49736
rect 98698 49680 101916 49736
rect 98637 49678 101916 49680
rect 101998 49678 103848 49738
rect 105721 49738 105787 49741
rect 107744 49738 107804 50048
rect 105721 49736 107804 49738
rect 105721 49680 105726 49736
rect 105782 49680 107804 49736
rect 105721 49678 107804 49680
rect 108481 49738 108547 49741
rect 110596 49738 110656 50048
rect 111057 49874 111123 49877
rect 113540 49874 113600 50048
rect 111057 49872 113600 49874
rect 111057 49816 111062 49872
rect 111118 49816 113600 49872
rect 111057 49814 113600 49816
rect 111057 49811 111123 49814
rect 108481 49736 110656 49738
rect 108481 49680 108486 49736
rect 108542 49680 110656 49736
rect 108481 49678 110656 49680
rect 112621 49738 112687 49741
rect 114552 49738 114612 50048
rect 116669 50010 116735 50013
rect 117404 50010 117464 50048
rect 116669 50008 117464 50010
rect 116669 49952 116674 50008
rect 116730 49952 117464 50008
rect 116669 49950 117464 49952
rect 116669 49947 116735 49950
rect 115197 49874 115263 49877
rect 118416 49874 118476 50048
rect 115197 49872 118476 49874
rect 115197 49816 115202 49872
rect 115258 49816 118476 49872
rect 115197 49814 118476 49816
rect 118601 49874 118667 49877
rect 120214 49874 120274 50222
rect 121360 50116 121420 50222
rect 122280 50116 122340 50358
rect 123477 50416 126296 50418
rect 123477 50360 123482 50416
rect 123538 50360 126296 50416
rect 123477 50358 126296 50360
rect 123477 50355 123543 50358
rect 122465 50282 122531 50285
rect 122465 50280 125284 50282
rect 122465 50224 122470 50280
rect 122526 50224 125284 50280
rect 122465 50222 125284 50224
rect 122465 50219 122531 50222
rect 125224 50116 125284 50222
rect 126236 50116 126296 50358
rect 131757 50416 135036 50418
rect 131757 50360 131762 50416
rect 131818 50360 135036 50416
rect 131757 50358 135036 50360
rect 131757 50355 131823 50358
rect 126421 50282 126487 50285
rect 129273 50282 129339 50285
rect 126421 50280 129148 50282
rect 126421 50224 126426 50280
rect 126482 50224 129148 50280
rect 126421 50222 129148 50224
rect 126421 50219 126487 50222
rect 129088 50116 129148 50222
rect 129273 50280 132092 50282
rect 129273 50224 129278 50280
rect 129334 50224 132092 50280
rect 129273 50222 132092 50224
rect 129273 50219 129339 50222
rect 132032 50116 132092 50222
rect 132450 50222 133104 50282
rect 118601 49872 120274 49874
rect 118601 49816 118606 49872
rect 118662 49816 120274 49872
rect 118601 49814 120274 49816
rect 115197 49811 115263 49814
rect 118601 49811 118667 49814
rect 112621 49736 114612 49738
rect 112621 49680 112626 49736
rect 112682 49680 114612 49736
rect 112621 49678 114612 49680
rect 115381 49738 115447 49741
rect 116669 49738 116735 49741
rect 115381 49736 116735 49738
rect 115381 49680 115386 49736
rect 115442 49680 116674 49736
rect 116730 49680 116735 49736
rect 115381 49678 116735 49680
rect 98637 49675 98703 49678
rect 101397 49602 101463 49605
rect 101998 49602 102058 49678
rect 105721 49675 105787 49678
rect 108481 49675 108547 49678
rect 112621 49675 112687 49678
rect 115381 49675 115447 49678
rect 116669 49675 116735 49678
rect 117957 49738 118023 49741
rect 120348 49738 120408 50048
rect 120717 49874 120783 49877
rect 123292 49874 123352 50048
rect 120717 49872 123352 49874
rect 120717 49816 120722 49872
rect 120778 49816 123352 49872
rect 120717 49814 123352 49816
rect 120717 49811 120783 49814
rect 117957 49736 120408 49738
rect 117957 49680 117962 49736
rect 118018 49680 120408 49736
rect 117957 49678 120408 49680
rect 122097 49738 122163 49741
rect 124304 49738 124364 50048
rect 126513 50010 126579 50013
rect 127156 50010 127216 50048
rect 128168 50010 128228 50048
rect 126513 50008 127216 50010
rect 126513 49952 126518 50008
rect 126574 49952 127216 50008
rect 126513 49950 127216 49952
rect 127390 49950 128228 50010
rect 126513 49947 126579 49950
rect 125041 49874 125107 49877
rect 127390 49874 127450 49950
rect 125041 49872 127450 49874
rect 125041 49816 125046 49872
rect 125102 49816 127450 49872
rect 125041 49814 127450 49816
rect 127617 49874 127683 49877
rect 130100 49874 130160 50048
rect 127617 49872 130160 49874
rect 127617 49816 127622 49872
rect 127678 49816 130160 49872
rect 127617 49814 130160 49816
rect 125041 49811 125107 49814
rect 127617 49811 127683 49814
rect 122097 49736 124364 49738
rect 122097 49680 122102 49736
rect 122158 49680 124364 49736
rect 122097 49678 124364 49680
rect 124857 49738 124923 49741
rect 126513 49738 126579 49741
rect 124857 49736 126579 49738
rect 124857 49680 124862 49736
rect 124918 49680 126518 49736
rect 126574 49680 126579 49736
rect 124857 49678 126579 49680
rect 117957 49675 118023 49678
rect 122097 49675 122163 49678
rect 124857 49675 124923 49678
rect 126513 49675 126579 49678
rect 128997 49738 129063 49741
rect 131112 49738 131172 50048
rect 132450 49874 132510 50222
rect 133044 50116 133104 50222
rect 134976 50116 135036 50358
rect 135896 50116 135956 50494
rect 142797 50552 145708 50554
rect 142797 50496 142802 50552
rect 142858 50496 145708 50552
rect 142797 50494 145708 50496
rect 142797 50491 142863 50494
rect 138657 50418 138723 50421
rect 141601 50418 141667 50421
rect 138657 50416 141434 50418
rect 138657 50360 138662 50416
rect 138718 50360 141434 50416
rect 138657 50358 141434 50360
rect 138657 50355 138723 50358
rect 136081 50282 136147 50285
rect 140037 50282 140103 50285
rect 141374 50282 141434 50358
rect 141601 50416 144788 50418
rect 141601 50360 141606 50416
rect 141662 50360 144788 50416
rect 141601 50358 144788 50360
rect 141601 50355 141667 50358
rect 136081 50280 138900 50282
rect 136081 50224 136086 50280
rect 136142 50224 138900 50280
rect 136081 50222 138900 50224
rect 136081 50219 136147 50222
rect 138840 50116 138900 50222
rect 140037 50280 141066 50282
rect 140037 50224 140042 50280
rect 140098 50224 141066 50280
rect 140037 50222 141066 50224
rect 141374 50222 141844 50282
rect 140037 50219 140103 50222
rect 128997 49736 131172 49738
rect 128997 49680 129002 49736
rect 129058 49680 131172 49736
rect 128997 49678 131172 49680
rect 131254 49814 132510 49874
rect 128997 49675 129063 49678
rect 101397 49600 102058 49602
rect 101397 49544 101402 49600
rect 101458 49544 102058 49600
rect 101397 49542 102058 49544
rect 130377 49602 130443 49605
rect 131254 49602 131314 49814
rect 131941 49738 132007 49741
rect 133964 49738 134024 50048
rect 136173 50010 136239 50013
rect 136908 50010 136968 50048
rect 137920 50010 137980 50048
rect 136173 50008 136968 50010
rect 136173 49952 136178 50008
rect 136234 49952 136968 50008
rect 136173 49950 136968 49952
rect 137142 49950 137980 50010
rect 136173 49947 136239 49950
rect 134701 49874 134767 49877
rect 137142 49874 137202 49950
rect 134701 49872 137202 49874
rect 134701 49816 134706 49872
rect 134762 49816 137202 49872
rect 134701 49814 137202 49816
rect 137277 49874 137343 49877
rect 139852 49874 139912 50048
rect 137277 49872 139912 49874
rect 137277 49816 137282 49872
rect 137338 49816 139912 49872
rect 137277 49814 139912 49816
rect 134701 49811 134767 49814
rect 137277 49811 137343 49814
rect 131941 49736 134024 49738
rect 131941 49680 131946 49736
rect 132002 49680 134024 49736
rect 131941 49678 134024 49680
rect 134517 49738 134583 49741
rect 136173 49738 136239 49741
rect 134517 49736 136239 49738
rect 134517 49680 134522 49736
rect 134578 49680 136178 49736
rect 136234 49680 136239 49736
rect 134517 49678 136239 49680
rect 131941 49675 132007 49678
rect 134517 49675 134583 49678
rect 136173 49675 136239 49678
rect 138841 49738 138907 49741
rect 140772 49738 140832 50048
rect 141006 49874 141066 50222
rect 141784 50116 141844 50222
rect 144728 50116 144788 50358
rect 145648 50116 145708 50494
rect 152457 50552 155460 50554
rect 152457 50496 152462 50552
rect 152518 50496 155460 50552
rect 152457 50494 155460 50496
rect 152457 50491 152523 50494
rect 148501 50418 148567 50421
rect 151077 50418 151143 50421
rect 148501 50416 151002 50418
rect 148501 50360 148506 50416
rect 148562 50360 151002 50416
rect 148501 50358 151002 50360
rect 148501 50355 148567 50358
rect 145833 50282 145899 50285
rect 148317 50282 148383 50285
rect 150942 50282 151002 50358
rect 151077 50416 154540 50418
rect 151077 50360 151082 50416
rect 151138 50360 154540 50416
rect 151077 50358 154540 50360
rect 151077 50355 151143 50358
rect 151721 50282 151787 50285
rect 145833 50280 147874 50282
rect 145833 50224 145838 50280
rect 145894 50224 147874 50280
rect 145833 50222 147874 50224
rect 145833 50219 145899 50222
rect 147814 50146 147874 50222
rect 148317 50280 150584 50282
rect 148317 50224 148322 50280
rect 148378 50224 150584 50280
rect 148317 50222 150584 50224
rect 150942 50222 151596 50282
rect 148317 50219 148383 50222
rect 147814 50086 148622 50146
rect 150524 50116 150584 50222
rect 151536 50116 151596 50222
rect 151721 50280 152516 50282
rect 151721 50224 151726 50280
rect 151782 50224 152516 50280
rect 151721 50222 152516 50224
rect 151721 50219 151787 50222
rect 152456 50116 152516 50222
rect 154480 50116 154540 50358
rect 155400 50116 155460 50494
rect 160737 50552 164200 50554
rect 160737 50496 160742 50552
rect 160798 50496 164200 50552
rect 160737 50494 164200 50496
rect 160737 50491 160803 50494
rect 155585 50418 155651 50421
rect 157793 50418 157859 50421
rect 155585 50416 157859 50418
rect 155585 50360 155590 50416
rect 155646 50360 157798 50416
rect 157854 50360 157859 50416
rect 155585 50358 157859 50360
rect 155585 50355 155651 50358
rect 157793 50355 157859 50358
rect 156597 50282 156663 50285
rect 159449 50282 159515 50285
rect 156597 50280 159324 50282
rect 156597 50224 156602 50280
rect 156658 50224 159324 50280
rect 156597 50222 159324 50224
rect 156597 50219 156663 50222
rect 157793 50146 157859 50149
rect 157793 50144 158374 50146
rect 157793 50088 157798 50144
rect 157854 50088 158374 50144
rect 159264 50116 159324 50222
rect 159449 50280 162268 50282
rect 159449 50224 159454 50280
rect 159510 50224 162268 50280
rect 159449 50222 162268 50224
rect 159449 50219 159515 50222
rect 162208 50116 162268 50222
rect 164140 50116 164200 50494
rect 165152 50116 165212 50630
rect 178677 50688 180767 50690
rect 178677 50632 178682 50688
rect 178738 50632 180706 50688
rect 180762 50632 180767 50688
rect 178677 50630 180767 50632
rect 178677 50627 178743 50630
rect 180701 50627 180767 50630
rect 181437 50690 181503 50693
rect 181437 50688 183704 50690
rect 181437 50632 181442 50688
rect 181498 50632 183704 50688
rect 181437 50630 183704 50632
rect 181437 50627 181503 50630
rect 170397 50554 170463 50557
rect 180057 50554 180123 50557
rect 170397 50552 173032 50554
rect 170397 50496 170402 50552
rect 170458 50496 173032 50552
rect 170397 50494 173032 50496
rect 170397 50491 170463 50494
rect 165337 50418 165403 50421
rect 167637 50418 167703 50421
rect 165337 50416 167703 50418
rect 165337 50360 165342 50416
rect 165398 50360 167642 50416
rect 167698 50360 167703 50416
rect 165337 50358 167703 50360
rect 165337 50355 165403 50358
rect 167637 50355 167703 50358
rect 167821 50418 167887 50421
rect 167821 50416 171008 50418
rect 167821 50360 167826 50416
rect 167882 50360 171008 50416
rect 167821 50358 171008 50360
rect 167821 50355 167887 50358
rect 166257 50282 166323 50285
rect 167637 50282 167703 50285
rect 166257 50280 167562 50282
rect 166257 50224 166262 50280
rect 166318 50224 167562 50280
rect 166257 50222 167562 50224
rect 166257 50219 166323 50222
rect 157793 50086 158374 50088
rect 157793 50083 157859 50086
rect 142796 49874 142856 50048
rect 141006 49814 142856 49874
rect 138841 49736 140832 49738
rect 138841 49680 138846 49736
rect 138902 49680 140832 49736
rect 138841 49678 140832 49680
rect 141417 49738 141483 49741
rect 143716 49738 143776 50048
rect 145925 50010 145991 50013
rect 146660 50010 146720 50048
rect 145925 50008 146720 50010
rect 145925 49952 145930 50008
rect 145986 49952 146720 50008
rect 145925 49950 146720 49952
rect 145925 49947 145991 49950
rect 144177 49874 144243 49877
rect 147580 49874 147640 50048
rect 144177 49872 147640 49874
rect 144177 49816 144182 49872
rect 144238 49816 147640 49872
rect 144177 49814 147640 49816
rect 144177 49811 144243 49814
rect 141417 49736 143776 49738
rect 141417 49680 141422 49736
rect 141478 49680 143776 49736
rect 141417 49678 143776 49680
rect 144361 49738 144427 49741
rect 145925 49738 145991 49741
rect 144361 49736 145991 49738
rect 144361 49680 144366 49736
rect 144422 49680 145930 49736
rect 145986 49680 145991 49736
rect 144361 49678 145991 49680
rect 138841 49675 138907 49678
rect 141417 49675 141483 49678
rect 144361 49675 144427 49678
rect 145925 49675 145991 49678
rect 146937 49738 147003 49741
rect 149604 49738 149664 50048
rect 150525 49874 150591 49877
rect 153468 49874 153528 50048
rect 150525 49872 153528 49874
rect 150525 49816 150530 49872
rect 150586 49816 153528 49872
rect 150525 49814 153528 49816
rect 153837 49874 153903 49877
rect 156412 49874 156472 50048
rect 153837 49872 156472 49874
rect 153837 49816 153842 49872
rect 153898 49816 156472 49872
rect 153837 49814 156472 49816
rect 150525 49811 150591 49814
rect 153837 49811 153903 49814
rect 146937 49736 149664 49738
rect 146937 49680 146942 49736
rect 146998 49680 149664 49736
rect 146937 49678 149664 49680
rect 149789 49738 149855 49741
rect 151721 49738 151787 49741
rect 149789 49736 151787 49738
rect 149789 49680 149794 49736
rect 149850 49680 151726 49736
rect 151782 49680 151787 49736
rect 149789 49678 151787 49680
rect 146937 49675 147003 49678
rect 149789 49675 149855 49678
rect 151721 49675 151787 49678
rect 155401 49738 155467 49741
rect 157332 49738 157392 50048
rect 159541 50010 159607 50013
rect 160276 50010 160336 50048
rect 159541 50008 160336 50010
rect 159541 49952 159546 50008
rect 159602 49952 160336 50008
rect 159541 49950 160336 49952
rect 159541 49947 159607 49950
rect 158161 49874 158227 49877
rect 161288 49874 161348 50048
rect 158161 49872 161348 49874
rect 158161 49816 158166 49872
rect 158222 49816 161348 49872
rect 158161 49814 161348 49816
rect 158161 49811 158227 49814
rect 155401 49736 157392 49738
rect 155401 49680 155406 49736
rect 155462 49680 157392 49736
rect 155401 49678 157392 49680
rect 157977 49738 158043 49741
rect 159541 49738 159607 49741
rect 157977 49736 159607 49738
rect 157977 49680 157982 49736
rect 158038 49680 159546 49736
rect 159602 49680 159607 49736
rect 157977 49678 159607 49680
rect 155401 49675 155467 49678
rect 157977 49675 158043 49678
rect 159541 49675 159607 49678
rect 160921 49738 160987 49741
rect 163220 49738 163280 50048
rect 163497 49874 163563 49877
rect 166072 49874 166132 50048
rect 163497 49872 166132 49874
rect 163497 49816 163502 49872
rect 163558 49816 166132 49872
rect 163497 49814 166132 49816
rect 163497 49811 163563 49814
rect 160921 49736 163280 49738
rect 160921 49680 160926 49736
rect 160982 49680 163280 49736
rect 160921 49678 163280 49680
rect 165061 49738 165127 49741
rect 167084 49738 167144 50048
rect 167502 49874 167562 50222
rect 167637 50280 170088 50282
rect 167637 50224 167642 50280
rect 167698 50224 170088 50280
rect 167637 50222 170088 50224
rect 167637 50219 167703 50222
rect 167729 50146 167795 50149
rect 167729 50144 168126 50146
rect 167729 50088 167734 50144
rect 167790 50088 168126 50144
rect 170028 50116 170088 50222
rect 170948 50116 171008 50358
rect 172972 50116 173032 50494
rect 180057 50552 182692 50554
rect 180057 50496 180062 50552
rect 180118 50496 182692 50552
rect 180057 50494 182692 50496
rect 180057 50491 180123 50494
rect 174721 50418 174787 50421
rect 177113 50418 177179 50421
rect 174721 50416 177179 50418
rect 174721 50360 174726 50416
rect 174782 50360 177118 50416
rect 177174 50360 177179 50416
rect 174721 50358 177179 50360
rect 174721 50355 174787 50358
rect 177113 50355 177179 50358
rect 177481 50418 177547 50421
rect 180701 50418 180767 50421
rect 177481 50416 180626 50418
rect 177481 50360 177486 50416
rect 177542 50360 180626 50416
rect 177481 50358 180626 50360
rect 177481 50355 177547 50358
rect 173157 50282 173223 50285
rect 176009 50282 176075 50285
rect 180566 50282 180626 50358
rect 180701 50416 181772 50418
rect 180701 50360 180706 50416
rect 180762 50360 181772 50416
rect 180701 50358 181772 50360
rect 180701 50355 180767 50358
rect 173157 50280 175884 50282
rect 173157 50224 173162 50280
rect 173218 50224 175884 50280
rect 173157 50222 175884 50224
rect 173157 50219 173223 50222
rect 175824 50116 175884 50222
rect 176009 50280 178828 50282
rect 176009 50224 176014 50280
rect 176070 50224 178828 50280
rect 176009 50222 178828 50224
rect 180566 50222 180760 50282
rect 176009 50219 176075 50222
rect 177113 50146 177179 50149
rect 177113 50144 177786 50146
rect 167729 50086 168126 50088
rect 177113 50088 177118 50144
rect 177174 50088 177786 50144
rect 178768 50116 178828 50222
rect 180700 50116 180760 50222
rect 181712 50116 181772 50358
rect 182632 50116 182692 50494
rect 183644 50116 183704 50630
rect 184656 50116 184716 50766
rect 446488 50824 449223 50826
rect 446488 50768 449162 50824
rect 449218 50768 449223 50824
rect 446488 50766 449223 50768
rect 200757 50690 200823 50693
rect 278681 50690 278747 50693
rect 288341 50690 288407 50693
rect 363045 50690 363111 50693
rect 410517 50690 410583 50693
rect 200757 50688 203208 50690
rect 200757 50632 200762 50688
rect 200818 50632 203208 50688
rect 200757 50630 203208 50632
rect 200757 50627 200823 50630
rect 185577 50554 185643 50557
rect 195237 50554 195303 50557
rect 199377 50554 199443 50557
rect 185577 50552 188354 50554
rect 185577 50496 185582 50552
rect 185638 50496 188354 50552
rect 185577 50494 188354 50496
rect 185577 50491 185643 50494
rect 184841 50418 184907 50421
rect 184841 50416 187568 50418
rect 184841 50360 184846 50416
rect 184902 50360 187568 50416
rect 184841 50358 187568 50360
rect 184841 50355 184907 50358
rect 187508 50116 187568 50358
rect 188294 50282 188354 50494
rect 195237 50552 198332 50554
rect 195237 50496 195242 50552
rect 195298 50496 198332 50552
rect 195237 50494 198332 50496
rect 195237 50491 195303 50494
rect 188521 50418 188587 50421
rect 190913 50418 190979 50421
rect 193857 50418 193923 50421
rect 188521 50416 190979 50418
rect 188521 50360 188526 50416
rect 188582 50360 190918 50416
rect 190974 50360 190979 50416
rect 188521 50358 190979 50360
rect 188521 50355 188587 50358
rect 190913 50355 190979 50358
rect 191238 50358 192444 50418
rect 189717 50282 189783 50285
rect 191238 50282 191298 50358
rect 188294 50222 188580 50282
rect 188520 50116 188580 50222
rect 189717 50280 191298 50282
rect 189717 50224 189722 50280
rect 189778 50224 191298 50280
rect 189717 50222 191298 50224
rect 189717 50219 189783 50222
rect 190913 50146 190979 50149
rect 190913 50144 191494 50146
rect 177113 50086 177786 50088
rect 190913 50088 190918 50144
rect 190974 50088 191494 50144
rect 192384 50116 192444 50358
rect 193857 50416 197320 50418
rect 193857 50360 193862 50416
rect 193918 50360 197320 50416
rect 193857 50358 197320 50360
rect 193857 50355 193923 50358
rect 192569 50282 192635 50285
rect 192569 50280 195388 50282
rect 192569 50224 192574 50280
rect 192630 50224 195388 50280
rect 192569 50222 195388 50224
rect 192569 50219 192635 50222
rect 195328 50116 195388 50222
rect 197260 50116 197320 50358
rect 198272 50116 198332 50494
rect 199377 50552 202196 50554
rect 199377 50496 199382 50552
rect 199438 50496 202196 50552
rect 199377 50494 202196 50496
rect 199377 50491 199443 50494
rect 198457 50418 198523 50421
rect 198457 50416 201184 50418
rect 198457 50360 198462 50416
rect 198518 50360 201184 50416
rect 198457 50358 201184 50360
rect 198457 50355 198523 50358
rect 201124 50116 201184 50358
rect 202136 50116 202196 50494
rect 203148 50116 203208 50630
rect 278681 50688 281040 50690
rect 278681 50632 278686 50688
rect 278742 50632 281040 50688
rect 278681 50630 281040 50632
rect 278681 50627 278747 50630
rect 214557 50554 214623 50557
rect 221457 50554 221523 50557
rect 225597 50554 225663 50557
rect 227713 50554 227779 50557
rect 250989 50554 251055 50557
rect 259361 50554 259427 50557
rect 269021 50554 269087 50557
rect 277301 50554 277367 50557
rect 214557 50552 217744 50554
rect 214557 50496 214562 50552
rect 214618 50496 217744 50552
rect 214557 50494 217744 50496
rect 214557 50491 214623 50494
rect 211797 50418 211863 50421
rect 211797 50416 214800 50418
rect 211797 50360 211802 50416
rect 211858 50360 214800 50416
rect 211797 50358 214800 50360
rect 211797 50355 211863 50358
rect 203517 50282 203583 50285
rect 206277 50282 206343 50285
rect 209129 50282 209195 50285
rect 203517 50280 206060 50282
rect 203517 50224 203522 50280
rect 203578 50224 206060 50280
rect 203517 50222 206060 50224
rect 203517 50219 203583 50222
rect 206000 50116 206060 50222
rect 206277 50280 209004 50282
rect 206277 50224 206282 50280
rect 206338 50224 209004 50280
rect 206277 50222 209004 50224
rect 206277 50219 206343 50222
rect 208944 50116 209004 50222
rect 209129 50280 211948 50282
rect 209129 50224 209134 50280
rect 209190 50224 211948 50280
rect 209129 50222 211948 50224
rect 209129 50219 209195 50222
rect 211888 50116 211948 50222
rect 212582 50222 213880 50282
rect 190913 50086 191494 50088
rect 167729 50083 167795 50086
rect 177113 50083 177179 50086
rect 190913 50083 190979 50086
rect 169016 50010 169076 50048
rect 168790 49950 169076 50010
rect 168790 49874 168850 49950
rect 167502 49814 168850 49874
rect 169017 49874 169083 49877
rect 171960 49874 172020 50048
rect 173249 50010 173315 50013
rect 173892 50010 173952 50048
rect 173249 50008 173952 50010
rect 173249 49952 173254 50008
rect 173310 49952 173952 50008
rect 173249 49950 173952 49952
rect 173249 49947 173315 49950
rect 169017 49872 172020 49874
rect 169017 49816 169022 49872
rect 169078 49816 172020 49872
rect 169017 49814 172020 49816
rect 172145 49874 172211 49877
rect 174904 49874 174964 50048
rect 172145 49872 174964 49874
rect 172145 49816 172150 49872
rect 172206 49816 174964 49872
rect 172145 49814 174964 49816
rect 169017 49811 169083 49814
rect 172145 49811 172211 49814
rect 165061 49736 167144 49738
rect 165061 49680 165066 49736
rect 165122 49680 167144 49736
rect 165061 49678 167144 49680
rect 171777 49738 171843 49741
rect 173249 49738 173315 49741
rect 171777 49736 173315 49738
rect 171777 49680 171782 49736
rect 171838 49680 173254 49736
rect 173310 49680 173315 49736
rect 171777 49678 173315 49680
rect 160921 49675 160987 49678
rect 165061 49675 165127 49678
rect 171777 49675 171843 49678
rect 173249 49675 173315 49678
rect 174537 49738 174603 49741
rect 176836 49738 176896 50048
rect 174537 49736 176896 49738
rect 174537 49680 174542 49736
rect 174598 49680 176896 49736
rect 174537 49678 176896 49680
rect 177297 49738 177363 49741
rect 179780 49738 179840 50048
rect 182817 49874 182883 49877
rect 185576 49874 185636 50048
rect 182817 49872 185636 49874
rect 182817 49816 182822 49872
rect 182878 49816 185636 49872
rect 182817 49814 185636 49816
rect 182817 49811 182883 49814
rect 177297 49736 179840 49738
rect 177297 49680 177302 49736
rect 177358 49680 179840 49736
rect 177297 49678 179840 49680
rect 184197 49738 184263 49741
rect 186588 49738 186648 50048
rect 184197 49736 186648 49738
rect 184197 49680 184202 49736
rect 184258 49680 186648 49736
rect 184197 49678 186648 49680
rect 186957 49738 187023 49741
rect 189440 49738 189500 50048
rect 190452 49738 190512 50048
rect 192569 50010 192635 50013
rect 193396 50010 193456 50048
rect 192569 50008 193456 50010
rect 192569 49952 192574 50008
rect 192630 49952 193456 50008
rect 192569 49950 193456 49952
rect 192569 49947 192635 49950
rect 191097 49874 191163 49877
rect 194316 49874 194376 50048
rect 191097 49872 194376 49874
rect 191097 49816 191102 49872
rect 191158 49816 194376 49872
rect 191097 49814 194376 49816
rect 191097 49811 191163 49814
rect 186957 49736 189500 49738
rect 186957 49680 186962 49736
rect 187018 49680 189500 49736
rect 186957 49678 189500 49680
rect 189582 49678 190512 49738
rect 191281 49738 191347 49741
rect 192569 49738 192635 49741
rect 191281 49736 192635 49738
rect 191281 49680 191286 49736
rect 191342 49680 192574 49736
rect 192630 49680 192635 49736
rect 191281 49678 192635 49680
rect 174537 49675 174603 49678
rect 177297 49675 177363 49678
rect 184197 49675 184263 49678
rect 186957 49675 187023 49678
rect 130377 49600 131314 49602
rect 130377 49544 130382 49600
rect 130438 49544 131314 49600
rect 130377 49542 131314 49544
rect 188337 49602 188403 49605
rect 189582 49602 189642 49678
rect 191281 49675 191347 49678
rect 192569 49675 192635 49678
rect 194041 49738 194107 49741
rect 196248 49738 196308 50048
rect 194041 49736 196308 49738
rect 194041 49680 194046 49736
rect 194102 49680 196308 49736
rect 194041 49678 196308 49680
rect 196617 49738 196683 49741
rect 199192 49738 199252 50048
rect 200204 49738 200264 50048
rect 202137 49874 202203 49877
rect 203885 49874 203951 49877
rect 202137 49872 203951 49874
rect 202137 49816 202142 49872
rect 202198 49816 203890 49872
rect 203946 49816 203951 49872
rect 202137 49814 203951 49816
rect 202137 49811 202203 49814
rect 203885 49811 203951 49814
rect 196617 49736 199252 49738
rect 196617 49680 196622 49736
rect 196678 49680 199252 49736
rect 196617 49678 199252 49680
rect 199334 49678 200264 49738
rect 200941 49738 201007 49741
rect 204068 49738 204128 50048
rect 204253 50010 204319 50013
rect 205080 50010 205140 50048
rect 207012 50010 207072 50048
rect 204253 50008 205140 50010
rect 204253 49952 204258 50008
rect 204314 49952 205140 50008
rect 204253 49950 205140 49952
rect 206878 49950 207072 50010
rect 204253 49947 204319 49950
rect 204897 49874 204963 49877
rect 206878 49874 206938 49950
rect 204897 49872 206938 49874
rect 204897 49816 204902 49872
rect 204958 49816 206938 49872
rect 204897 49814 206938 49816
rect 204897 49811 204963 49814
rect 200941 49736 204128 49738
rect 200941 49680 200946 49736
rect 201002 49680 204128 49736
rect 200941 49678 204128 49680
rect 205081 49738 205147 49741
rect 207932 49738 207992 50048
rect 209956 50010 210016 50048
rect 209086 49950 210016 50010
rect 208117 49874 208183 49877
rect 209086 49874 209146 49950
rect 210876 49874 210936 50048
rect 208117 49872 209146 49874
rect 208117 49816 208122 49872
rect 208178 49816 209146 49872
rect 208117 49814 209146 49816
rect 209730 49814 210936 49874
rect 211061 49874 211127 49877
rect 212582 49874 212642 50222
rect 213820 50116 213880 50222
rect 214740 50116 214800 50358
rect 214925 50282 214991 50285
rect 214925 50280 216824 50282
rect 214925 50224 214930 50280
rect 214986 50224 216824 50280
rect 214925 50222 216824 50224
rect 214925 50219 214991 50222
rect 216764 50116 216824 50222
rect 217684 50116 217744 50494
rect 221457 50552 224552 50554
rect 221457 50496 221462 50552
rect 221518 50496 224552 50552
rect 221457 50494 224552 50496
rect 221457 50491 221523 50494
rect 218697 50418 218763 50421
rect 218697 50416 221700 50418
rect 218697 50360 218702 50416
rect 218758 50360 221700 50416
rect 218697 50358 221700 50360
rect 218697 50355 218763 50358
rect 217918 50222 220688 50282
rect 211061 49872 212642 49874
rect 211061 49816 211066 49872
rect 211122 49816 212642 49872
rect 211061 49814 212642 49816
rect 208117 49811 208183 49814
rect 209730 49738 209790 49814
rect 211061 49811 211127 49814
rect 205081 49736 207992 49738
rect 205081 49680 205086 49736
rect 205142 49680 207992 49736
rect 205081 49678 207992 49680
rect 208166 49678 209790 49738
rect 210601 49738 210667 49741
rect 212808 49738 212868 50048
rect 210601 49736 212868 49738
rect 210601 49680 210606 49736
rect 210662 49680 212868 49736
rect 210601 49678 212868 49680
rect 213177 49738 213243 49741
rect 215752 49738 215812 50048
rect 217317 49874 217383 49877
rect 217918 49874 217978 50222
rect 220628 50116 220688 50222
rect 221640 50116 221700 50358
rect 221825 50282 221891 50285
rect 221825 50280 223632 50282
rect 221825 50224 221830 50280
rect 221886 50224 223632 50280
rect 221825 50222 223632 50224
rect 221825 50219 221891 50222
rect 223572 50116 223632 50222
rect 224492 50116 224552 50494
rect 225597 50552 227546 50554
rect 225597 50496 225602 50552
rect 225658 50496 227546 50552
rect 225597 50494 227546 50496
rect 225597 50491 225663 50494
rect 227486 50418 227546 50494
rect 227713 50552 231360 50554
rect 227713 50496 227718 50552
rect 227774 50496 231360 50552
rect 227713 50494 231360 50496
rect 227713 50491 227779 50494
rect 227486 50358 228508 50418
rect 224677 50282 224743 50285
rect 224677 50280 226810 50282
rect 224677 50224 224682 50280
rect 224738 50224 226810 50280
rect 224677 50222 226810 50224
rect 224677 50219 224743 50222
rect 226750 50146 226810 50222
rect 226750 50086 227466 50146
rect 228448 50116 228508 50358
rect 229050 50222 230440 50282
rect 217317 49872 217978 49874
rect 217317 49816 217322 49872
rect 217378 49816 217978 49872
rect 217317 49814 217978 49816
rect 217317 49811 217383 49814
rect 213177 49736 215812 49738
rect 213177 49680 213182 49736
rect 213238 49680 215812 49736
rect 213177 49678 215812 49680
rect 215937 49738 216003 49741
rect 218696 49738 218756 50048
rect 219616 49738 219676 50048
rect 215937 49736 218756 49738
rect 215937 49680 215942 49736
rect 215998 49680 218756 49736
rect 215937 49678 218756 49680
rect 218838 49678 219676 49738
rect 220077 49738 220143 49741
rect 222560 49738 222620 50048
rect 222837 49874 222903 49877
rect 225504 49874 225564 50048
rect 222837 49872 225564 49874
rect 222837 49816 222842 49872
rect 222898 49816 225564 49872
rect 222837 49814 225564 49816
rect 222837 49811 222903 49814
rect 220077 49736 222620 49738
rect 220077 49680 220082 49736
rect 220138 49680 222620 49736
rect 220077 49678 222620 49680
rect 224401 49738 224467 49741
rect 226424 49738 226484 50048
rect 226977 49874 227043 49877
rect 229050 49874 229110 50222
rect 230380 50116 230440 50222
rect 231300 50116 231360 50494
rect 250989 50552 252202 50554
rect 250989 50496 250994 50552
rect 251050 50496 252202 50552
rect 250989 50494 252202 50496
rect 250989 50491 251055 50494
rect 233141 50418 233207 50421
rect 234429 50418 234495 50421
rect 249701 50418 249767 50421
rect 233141 50416 234354 50418
rect 233141 50360 233146 50416
rect 233202 50360 234354 50416
rect 233141 50358 234354 50360
rect 233141 50355 233207 50358
rect 231485 50282 231551 50285
rect 234294 50282 234354 50358
rect 234429 50416 235642 50418
rect 234429 50360 234434 50416
rect 234490 50360 235642 50416
rect 234429 50358 235642 50360
rect 234429 50355 234495 50358
rect 231485 50280 233618 50282
rect 231485 50224 231490 50280
rect 231546 50224 233618 50280
rect 231485 50222 233618 50224
rect 234294 50222 235316 50282
rect 231485 50219 231551 50222
rect 233558 50146 233618 50222
rect 233558 50086 234274 50146
rect 235256 50116 235316 50222
rect 235582 50146 235642 50358
rect 249701 50416 251876 50418
rect 249701 50360 249706 50416
rect 249762 50360 251876 50416
rect 249701 50358 251876 50360
rect 249701 50355 249767 50358
rect 235901 50282 235967 50285
rect 238477 50282 238543 50285
rect 241421 50282 241487 50285
rect 248045 50282 248111 50285
rect 235901 50280 238168 50282
rect 235901 50224 235906 50280
rect 235962 50224 238168 50280
rect 235901 50222 238168 50224
rect 235901 50219 235967 50222
rect 235582 50086 236206 50146
rect 238108 50116 238168 50222
rect 238477 50280 241112 50282
rect 238477 50224 238482 50280
rect 238538 50224 241112 50280
rect 238477 50222 241112 50224
rect 238477 50219 238543 50222
rect 241052 50116 241112 50222
rect 241421 50280 244056 50282
rect 241421 50224 241426 50280
rect 241482 50224 244056 50280
rect 241421 50222 244056 50224
rect 241421 50219 241487 50222
rect 243996 50116 244056 50222
rect 248045 50280 250864 50282
rect 248045 50224 248050 50280
rect 248106 50224 250864 50280
rect 248045 50222 250864 50224
rect 248045 50219 248111 50222
rect 250804 50116 250864 50222
rect 251816 50116 251876 50358
rect 252142 50146 252202 50494
rect 259361 50552 261536 50554
rect 259361 50496 259366 50552
rect 259422 50496 261536 50552
rect 259361 50494 261536 50496
rect 259361 50491 259427 50494
rect 253749 50418 253815 50421
rect 253749 50416 256660 50418
rect 253749 50360 253754 50416
rect 253810 50360 256660 50416
rect 253749 50358 256660 50360
rect 253749 50355 253815 50358
rect 253565 50282 253631 50285
rect 253565 50280 255740 50282
rect 253565 50224 253570 50280
rect 253626 50224 255740 50280
rect 253565 50222 255740 50224
rect 253565 50219 253631 50222
rect 252142 50086 252766 50146
rect 255680 50116 255740 50222
rect 256600 50116 256660 50358
rect 257889 50282 257955 50285
rect 257889 50280 260616 50282
rect 257889 50224 257894 50280
rect 257950 50224 260616 50280
rect 257889 50222 260616 50224
rect 257889 50219 257955 50222
rect 260556 50116 260616 50222
rect 261476 50116 261536 50494
rect 269021 50552 271288 50554
rect 269021 50496 269026 50552
rect 269082 50496 271288 50552
rect 269021 50494 271288 50496
rect 269021 50491 269087 50494
rect 266261 50418 266327 50421
rect 266261 50416 268344 50418
rect 266261 50360 266266 50416
rect 266322 50360 268344 50416
rect 266261 50358 268344 50360
rect 266261 50355 266327 50358
rect 262121 50282 262187 50285
rect 264789 50282 264855 50285
rect 262121 50280 264480 50282
rect 262121 50224 262126 50280
rect 262182 50224 264480 50280
rect 262121 50222 264480 50224
rect 262121 50219 262187 50222
rect 264420 50116 264480 50222
rect 264789 50280 267424 50282
rect 264789 50224 264794 50280
rect 264850 50224 267424 50280
rect 264789 50222 267424 50224
rect 264789 50219 264855 50222
rect 267364 50116 267424 50222
rect 268284 50116 268344 50358
rect 269070 50222 270368 50282
rect 226977 49872 229110 49874
rect 226977 49816 226982 49872
rect 227038 49816 229110 49872
rect 226977 49814 229110 49816
rect 226977 49811 227043 49814
rect 224401 49736 226484 49738
rect 224401 49680 224406 49736
rect 224462 49680 226484 49736
rect 224401 49678 226484 49680
rect 227161 49738 227227 49741
rect 229368 49738 229428 50048
rect 230381 49874 230447 49877
rect 232312 49874 232372 50048
rect 230381 49872 232372 49874
rect 230381 49816 230386 49872
rect 230442 49816 232372 49872
rect 230381 49814 232372 49816
rect 230381 49811 230447 49814
rect 227161 49736 229428 49738
rect 227161 49680 227166 49736
rect 227222 49680 229428 49736
rect 227161 49678 229428 49680
rect 231669 49738 231735 49741
rect 233324 49738 233384 50048
rect 234521 49874 234587 49877
rect 237188 49874 237248 50048
rect 239120 49874 239180 50048
rect 234521 49872 237248 49874
rect 234521 49816 234526 49872
rect 234582 49816 237248 49872
rect 234521 49814 237248 49816
rect 237422 49814 239180 49874
rect 234521 49811 234587 49814
rect 231669 49736 233384 49738
rect 231669 49680 231674 49736
rect 231730 49680 233384 49736
rect 231669 49678 233384 49680
rect 237281 49738 237347 49741
rect 237422 49738 237482 49814
rect 237281 49736 237482 49738
rect 237281 49680 237286 49736
rect 237342 49680 237482 49736
rect 237281 49678 237482 49680
rect 238661 49738 238727 49741
rect 240132 49738 240192 50048
rect 242064 50010 242124 50048
rect 242709 50010 242775 50013
rect 242064 50008 242775 50010
rect 242064 49952 242714 50008
rect 242770 49952 242775 50008
rect 242064 49950 242775 49952
rect 242709 49947 242775 49950
rect 241237 49874 241303 49877
rect 242984 49874 243044 50048
rect 241237 49872 243044 49874
rect 241237 49816 241242 49872
rect 241298 49816 243044 49872
rect 241237 49814 243044 49816
rect 241237 49811 241303 49814
rect 238661 49736 240192 49738
rect 238661 49680 238666 49736
rect 238722 49680 240192 49736
rect 238661 49678 240192 49680
rect 242801 49738 242867 49741
rect 244916 49738 244976 50048
rect 245928 49874 245988 50048
rect 246757 50010 246823 50013
rect 246940 50010 247000 50048
rect 246757 50008 247000 50010
rect 246757 49952 246762 50008
rect 246818 49952 247000 50008
rect 246757 49950 247000 49952
rect 246757 49947 246823 49950
rect 246941 49874 247007 49877
rect 245928 49872 247007 49874
rect 245928 49816 246946 49872
rect 247002 49816 247007 49872
rect 245928 49814 247007 49816
rect 246941 49811 247007 49814
rect 242801 49736 244976 49738
rect 242801 49680 242806 49736
rect 242862 49680 244976 49736
rect 242801 49678 244976 49680
rect 245561 49738 245627 49741
rect 247860 49738 247920 50048
rect 248872 49874 248932 50048
rect 245561 49736 247920 49738
rect 245561 49680 245566 49736
rect 245622 49680 247920 49736
rect 245561 49678 247920 49680
rect 248094 49814 248932 49874
rect 194041 49675 194107 49678
rect 196617 49675 196683 49678
rect 188337 49600 189642 49602
rect 188337 49544 188342 49600
rect 188398 49544 189642 49600
rect 188337 49542 189642 49544
rect 198181 49602 198247 49605
rect 199334 49602 199394 49678
rect 200941 49675 201007 49678
rect 205081 49675 205147 49678
rect 198181 49600 199394 49602
rect 198181 49544 198186 49600
rect 198242 49544 199394 49600
rect 198181 49542 199394 49544
rect 207657 49602 207723 49605
rect 208166 49602 208226 49678
rect 210601 49675 210667 49678
rect 213177 49675 213243 49678
rect 215937 49675 216003 49678
rect 207657 49600 208226 49602
rect 207657 49544 207662 49600
rect 207718 49544 208226 49600
rect 207657 49542 208226 49544
rect 217501 49602 217567 49605
rect 218838 49602 218898 49678
rect 220077 49675 220143 49678
rect 224401 49675 224467 49678
rect 227161 49675 227227 49678
rect 231669 49675 231735 49678
rect 237281 49675 237347 49678
rect 238661 49675 238727 49678
rect 242801 49675 242867 49678
rect 245561 49675 245627 49678
rect 217501 49600 218898 49602
rect 217501 49544 217506 49600
rect 217562 49544 218898 49600
rect 217501 49542 218898 49544
rect 246849 49602 246915 49605
rect 248094 49602 248154 49814
rect 248229 49738 248295 49741
rect 249792 49738 249852 50048
rect 253748 50010 253808 50048
rect 253614 49950 253808 50010
rect 250805 49874 250871 49877
rect 253614 49874 253674 49950
rect 250805 49872 253674 49874
rect 250805 49816 250810 49872
rect 250866 49816 253674 49872
rect 250805 49814 253674 49816
rect 250805 49811 250871 49814
rect 248229 49736 249852 49738
rect 248229 49680 248234 49736
rect 248290 49680 249852 49736
rect 248229 49678 249852 49680
rect 252461 49738 252527 49741
rect 254668 49738 254728 50048
rect 252461 49736 254728 49738
rect 252461 49680 252466 49736
rect 252522 49680 254728 49736
rect 252461 49678 254728 49680
rect 255221 49738 255287 49741
rect 257612 49738 257672 50048
rect 257797 49874 257863 49877
rect 258624 49874 258684 50048
rect 257797 49872 258684 49874
rect 257797 49816 257802 49872
rect 257858 49816 258684 49872
rect 257797 49814 258684 49816
rect 257797 49811 257863 49814
rect 255221 49736 257672 49738
rect 255221 49680 255226 49736
rect 255282 49680 257672 49736
rect 255221 49678 257672 49680
rect 257797 49738 257863 49741
rect 259544 49738 259604 50048
rect 260649 49874 260715 49877
rect 262305 49874 262371 49877
rect 260649 49872 262371 49874
rect 260649 49816 260654 49872
rect 260710 49816 262310 49872
rect 262366 49816 262371 49872
rect 260649 49814 262371 49816
rect 260649 49811 260715 49814
rect 262305 49811 262371 49814
rect 257797 49736 259604 49738
rect 257797 49680 257802 49736
rect 257858 49680 259604 49736
rect 257797 49678 259604 49680
rect 260465 49738 260531 49741
rect 262488 49738 262548 50048
rect 262673 50010 262739 50013
rect 263500 50010 263560 50048
rect 262673 50008 263560 50010
rect 262673 49952 262678 50008
rect 262734 49952 263560 50008
rect 262673 49950 263560 49952
rect 262673 49947 262739 49950
rect 263501 49874 263567 49877
rect 265432 49874 265492 50048
rect 263501 49872 265492 49874
rect 263501 49816 263506 49872
rect 263562 49816 265492 49872
rect 263501 49814 265492 49816
rect 263501 49811 263567 49814
rect 260465 49736 262548 49738
rect 260465 49680 260470 49736
rect 260526 49680 262548 49736
rect 260465 49678 262548 49680
rect 264605 49738 264671 49741
rect 266352 49738 266412 50048
rect 267549 49874 267615 49877
rect 269070 49874 269130 50222
rect 270308 50116 270368 50222
rect 271228 50116 271288 50494
rect 277301 50552 280028 50554
rect 277301 50496 277306 50552
rect 277362 50496 280028 50552
rect 277301 50494 280028 50496
rect 277301 50491 277367 50494
rect 271781 50282 271847 50285
rect 274357 50282 274423 50285
rect 271781 50280 274232 50282
rect 271781 50224 271786 50280
rect 271842 50224 274232 50280
rect 271781 50222 274232 50224
rect 271781 50219 271847 50222
rect 274172 50116 274232 50222
rect 274357 50280 277176 50282
rect 274357 50224 274362 50280
rect 274418 50224 277176 50280
rect 274357 50222 277176 50224
rect 274357 50219 274423 50222
rect 277116 50116 277176 50222
rect 279968 50116 280028 50494
rect 280980 50116 281040 50630
rect 288341 50688 290792 50690
rect 288341 50632 288346 50688
rect 288402 50632 290792 50688
rect 288341 50630 290792 50632
rect 288341 50627 288407 50630
rect 286685 50554 286751 50557
rect 286685 50552 288860 50554
rect 286685 50496 286690 50552
rect 286746 50496 288860 50552
rect 286685 50494 288860 50496
rect 286685 50491 286751 50494
rect 281165 50418 281231 50421
rect 285581 50418 285647 50421
rect 281165 50416 283984 50418
rect 281165 50360 281170 50416
rect 281226 50360 283984 50416
rect 281165 50358 283984 50360
rect 281165 50355 281231 50358
rect 283924 50116 283984 50358
rect 285581 50416 287848 50418
rect 285581 50360 285586 50416
rect 285642 50360 287848 50416
rect 285581 50358 287848 50360
rect 285581 50355 285647 50358
rect 287788 50116 287848 50358
rect 288800 50116 288860 50494
rect 290732 50116 290792 50630
rect 360836 50688 363111 50690
rect 360836 50632 363050 50688
rect 363106 50632 363111 50688
rect 360836 50630 363111 50632
rect 292481 50554 292547 50557
rect 315941 50554 316007 50557
rect 330477 50554 330543 50557
rect 335997 50554 336063 50557
rect 343633 50554 343699 50557
rect 354673 50554 354739 50557
rect 292481 50552 294656 50554
rect 292481 50496 292486 50552
rect 292542 50496 294656 50552
rect 292481 50494 294656 50496
rect 292481 50491 292547 50494
rect 290917 50418 290983 50421
rect 290917 50416 293736 50418
rect 290917 50360 290922 50416
rect 290978 50360 293736 50416
rect 290917 50358 293736 50360
rect 290917 50355 290983 50358
rect 293676 50116 293736 50358
rect 294596 50116 294656 50494
rect 315941 50552 318024 50554
rect 315941 50496 315946 50552
rect 316002 50496 318024 50552
rect 315941 50494 318024 50496
rect 315941 50491 316007 50494
rect 297725 50418 297791 50421
rect 304809 50418 304875 50421
rect 307477 50418 307543 50421
rect 314285 50418 314351 50421
rect 297725 50416 300544 50418
rect 297725 50360 297730 50416
rect 297786 50360 300544 50416
rect 297725 50358 300544 50360
rect 297725 50355 297791 50358
rect 295241 50282 295307 50285
rect 297909 50282 297975 50285
rect 295241 50280 297600 50282
rect 295241 50224 295246 50280
rect 295302 50224 297600 50280
rect 295241 50222 297600 50224
rect 295241 50219 295307 50222
rect 297540 50116 297600 50222
rect 297909 50280 299532 50282
rect 297909 50224 297914 50280
rect 297970 50224 299532 50280
rect 297909 50222 299532 50224
rect 297909 50219 297975 50222
rect 299472 50116 299532 50222
rect 300484 50116 300544 50358
rect 304809 50416 306390 50418
rect 304809 50360 304814 50416
rect 304870 50360 306390 50416
rect 304809 50358 306390 50360
rect 304809 50355 304875 50358
rect 300669 50282 300735 50285
rect 303521 50282 303587 50285
rect 306330 50282 306390 50358
rect 307477 50416 310204 50418
rect 307477 50360 307482 50416
rect 307538 50360 310204 50416
rect 307477 50358 310204 50360
rect 307477 50355 307543 50358
rect 307661 50282 307727 50285
rect 300669 50280 303396 50282
rect 300669 50224 300674 50280
rect 300730 50224 303396 50280
rect 300669 50222 303396 50224
rect 300669 50219 300735 50222
rect 303336 50116 303396 50222
rect 303521 50280 305746 50282
rect 303521 50224 303526 50280
rect 303582 50224 305746 50280
rect 303521 50222 305746 50224
rect 306330 50222 307352 50282
rect 303521 50219 303587 50222
rect 305686 50146 305746 50222
rect 305686 50086 306310 50146
rect 307292 50116 307352 50222
rect 307661 50280 309284 50282
rect 307661 50224 307666 50280
rect 307722 50224 309284 50280
rect 307661 50222 309284 50224
rect 307661 50219 307727 50222
rect 309224 50116 309284 50222
rect 310144 50116 310204 50358
rect 314285 50416 317012 50418
rect 314285 50360 314290 50416
rect 314346 50360 317012 50416
rect 314285 50358 317012 50360
rect 314285 50355 314351 50358
rect 310421 50282 310487 50285
rect 311801 50282 311867 50285
rect 310421 50280 311634 50282
rect 310421 50224 310426 50280
rect 310482 50224 311634 50280
rect 310421 50222 311634 50224
rect 310421 50219 310487 50222
rect 311574 50146 311634 50222
rect 311801 50280 314160 50282
rect 311801 50224 311806 50280
rect 311862 50224 314160 50280
rect 311801 50222 314160 50224
rect 311801 50219 311867 50222
rect 311574 50086 312198 50146
rect 314100 50116 314160 50222
rect 316952 50116 317012 50358
rect 317964 50116 318024 50494
rect 330477 50552 333572 50554
rect 330477 50496 330482 50552
rect 330538 50496 333572 50552
rect 330477 50494 333572 50496
rect 330477 50491 330543 50494
rect 324129 50418 324195 50421
rect 326153 50418 326219 50421
rect 327717 50418 327783 50421
rect 324129 50416 326219 50418
rect 324129 50360 324134 50416
rect 324190 50360 326158 50416
rect 326214 50360 326219 50416
rect 324129 50358 326219 50360
rect 324129 50355 324195 50358
rect 326153 50355 326219 50358
rect 326478 50358 326906 50418
rect 318701 50282 318767 50285
rect 321461 50282 321527 50285
rect 324957 50282 325023 50285
rect 326478 50282 326538 50358
rect 318701 50280 320968 50282
rect 318701 50224 318706 50280
rect 318762 50224 320968 50280
rect 318701 50222 320968 50224
rect 318701 50219 318767 50222
rect 320908 50116 320968 50222
rect 321461 50280 323912 50282
rect 321461 50224 321466 50280
rect 321522 50224 323912 50280
rect 321461 50222 323912 50224
rect 321461 50219 321527 50222
rect 323852 50116 323912 50222
rect 324957 50280 326538 50282
rect 324957 50224 324962 50280
rect 325018 50224 326538 50280
rect 324957 50222 326538 50224
rect 326846 50282 326906 50358
rect 327717 50416 330720 50418
rect 327717 50360 327722 50416
rect 327778 50360 330720 50416
rect 327717 50358 330720 50360
rect 327717 50355 327783 50358
rect 326846 50222 327776 50282
rect 324957 50219 325023 50222
rect 326153 50146 326219 50149
rect 326153 50144 326734 50146
rect 326153 50088 326158 50144
rect 326214 50088 326734 50144
rect 327716 50116 327776 50222
rect 328502 50222 329708 50282
rect 326153 50086 326734 50088
rect 326153 50083 326219 50086
rect 267549 49872 269130 49874
rect 267549 49816 267554 49872
rect 267610 49816 269130 49872
rect 267549 49814 269130 49816
rect 267549 49811 267615 49814
rect 264605 49736 266412 49738
rect 264605 49680 264610 49736
rect 264666 49680 266412 49736
rect 264605 49678 266412 49680
rect 267365 49738 267431 49741
rect 269296 49738 269356 50048
rect 270401 49874 270467 49877
rect 272057 49874 272123 49877
rect 270401 49872 272123 49874
rect 270401 49816 270406 49872
rect 270462 49816 272062 49872
rect 272118 49816 272123 49872
rect 270401 49814 272123 49816
rect 270401 49811 270467 49814
rect 272057 49811 272123 49814
rect 267365 49736 269356 49738
rect 267365 49680 267370 49736
rect 267426 49680 269356 49736
rect 267365 49678 269356 49680
rect 270217 49738 270283 49741
rect 272240 49738 272300 50048
rect 272425 50010 272491 50013
rect 273160 50010 273220 50048
rect 272425 50008 273220 50010
rect 272425 49952 272430 50008
rect 272486 49952 273220 50008
rect 272425 49950 273220 49952
rect 272425 49947 272491 49950
rect 273161 49874 273227 49877
rect 275092 49874 275152 50048
rect 273161 49872 275152 49874
rect 273161 49816 273166 49872
rect 273222 49816 275152 49872
rect 273161 49814 275152 49816
rect 273161 49811 273227 49814
rect 270217 49736 272300 49738
rect 270217 49680 270222 49736
rect 270278 49680 272300 49736
rect 270217 49678 272300 49680
rect 274541 49738 274607 49741
rect 276104 49738 276164 50048
rect 278036 49874 278096 50048
rect 274541 49736 276164 49738
rect 274541 49680 274546 49736
rect 274602 49680 276164 49736
rect 274541 49678 276164 49680
rect 276246 49814 278096 49874
rect 248229 49675 248295 49678
rect 252461 49675 252527 49678
rect 255221 49675 255287 49678
rect 257797 49675 257863 49678
rect 260465 49675 260531 49678
rect 264605 49675 264671 49678
rect 267365 49675 267431 49678
rect 270217 49675 270283 49678
rect 274541 49675 274607 49678
rect 246849 49600 248154 49602
rect 246849 49544 246854 49600
rect 246910 49544 248154 49600
rect 246849 49542 248154 49544
rect 275921 49602 275987 49605
rect 276246 49602 276306 49814
rect 277209 49738 277275 49741
rect 279048 49738 279108 50048
rect 281992 49874 282052 50048
rect 282729 49874 282795 49877
rect 281992 49872 282795 49874
rect 281992 49816 282734 49872
rect 282790 49816 282795 49872
rect 281992 49814 282795 49816
rect 282729 49811 282795 49814
rect 277209 49736 279108 49738
rect 277209 49680 277214 49736
rect 277270 49680 279108 49736
rect 277209 49678 279108 49680
rect 281349 49738 281415 49741
rect 282912 49738 282972 50048
rect 283097 49874 283163 49877
rect 284844 49874 284904 50048
rect 283097 49872 284904 49874
rect 283097 49816 283102 49872
rect 283158 49816 284904 49872
rect 283097 49814 284904 49816
rect 285856 49874 285916 50048
rect 286317 49874 286383 49877
rect 285856 49872 286383 49874
rect 285856 49816 286322 49872
rect 286378 49816 286383 49872
rect 285856 49814 286383 49816
rect 283097 49811 283163 49814
rect 286317 49811 286383 49814
rect 281349 49736 282972 49738
rect 281349 49680 281354 49736
rect 281410 49680 282972 49736
rect 281349 49678 282972 49680
rect 284017 49738 284083 49741
rect 286776 49738 286836 50048
rect 286961 49874 287027 49877
rect 289720 49874 289780 50048
rect 291652 49874 291712 50048
rect 286961 49872 289780 49874
rect 286961 49816 286966 49872
rect 287022 49816 289780 49872
rect 286961 49814 289780 49816
rect 290782 49814 291712 49874
rect 286961 49811 287027 49814
rect 284017 49736 286836 49738
rect 284017 49680 284022 49736
rect 284078 49680 286836 49736
rect 284017 49678 286836 49680
rect 289721 49738 289787 49741
rect 290782 49738 290842 49814
rect 289721 49736 290842 49738
rect 289721 49680 289726 49736
rect 289782 49680 290842 49736
rect 289721 49678 290842 49680
rect 291009 49738 291075 49741
rect 292664 49738 292724 50048
rect 293585 49874 293651 49877
rect 295608 49874 295668 50048
rect 293585 49872 295668 49874
rect 293585 49816 293590 49872
rect 293646 49816 295668 49872
rect 293585 49814 295668 49816
rect 293585 49811 293651 49814
rect 291009 49736 292724 49738
rect 291009 49680 291014 49736
rect 291070 49680 292724 49736
rect 291009 49678 292724 49680
rect 293769 49738 293835 49741
rect 296528 49738 296588 50048
rect 298460 49738 298520 50048
rect 299381 49874 299447 49877
rect 301404 49874 301464 50048
rect 299381 49872 301464 49874
rect 299381 49816 299386 49872
rect 299442 49816 301464 49872
rect 299381 49814 301464 49816
rect 299381 49811 299447 49814
rect 293769 49736 296588 49738
rect 293769 49680 293774 49736
rect 293830 49680 296588 49736
rect 293769 49678 296588 49680
rect 296670 49678 298520 49738
rect 300485 49738 300551 49741
rect 302416 49738 302476 50048
rect 304348 49874 304408 50048
rect 304901 49874 304967 49877
rect 304348 49872 304967 49874
rect 304348 49816 304906 49872
rect 304962 49816 304967 49872
rect 304348 49814 304967 49816
rect 304901 49811 304967 49814
rect 300485 49736 302476 49738
rect 300485 49680 300490 49736
rect 300546 49680 302476 49736
rect 300485 49678 302476 49680
rect 303521 49738 303587 49741
rect 305268 49738 305328 50048
rect 303521 49736 305328 49738
rect 303521 49680 303526 49736
rect 303582 49680 305328 49736
rect 303521 49678 305328 49680
rect 306281 49738 306347 49741
rect 308212 49738 308272 50048
rect 311156 50010 311216 50048
rect 311709 50010 311775 50013
rect 311156 50008 311775 50010
rect 311156 49952 311714 50008
rect 311770 49952 311775 50008
rect 311156 49950 311775 49952
rect 311709 49947 311775 49950
rect 310237 49874 310303 49877
rect 313088 49874 313148 50048
rect 310237 49872 313148 49874
rect 310237 49816 310242 49872
rect 310298 49816 313148 49872
rect 310237 49814 313148 49816
rect 310237 49811 310303 49814
rect 306281 49736 308272 49738
rect 306281 49680 306286 49736
rect 306342 49680 308272 49736
rect 306281 49678 308272 49680
rect 313181 49738 313247 49741
rect 315020 49738 315080 50048
rect 316032 49738 316092 50048
rect 318149 50010 318215 50013
rect 318976 50010 319036 50048
rect 318149 50008 319036 50010
rect 318149 49952 318154 50008
rect 318210 49952 319036 50008
rect 318149 49950 319036 49952
rect 318149 49947 318215 49950
rect 317137 49874 317203 49877
rect 319896 49874 319956 50048
rect 321093 50010 321159 50013
rect 321828 50010 321888 50048
rect 321093 50008 321888 50010
rect 321093 49952 321098 50008
rect 321154 49952 321888 50008
rect 321093 49950 321888 49952
rect 321093 49947 321159 49950
rect 317137 49872 319956 49874
rect 317137 49816 317142 49872
rect 317198 49816 319956 49872
rect 317137 49814 319956 49816
rect 320081 49874 320147 49877
rect 322840 49874 322900 50048
rect 320081 49872 322900 49874
rect 320081 49816 320086 49872
rect 320142 49816 322900 49872
rect 320081 49814 322900 49816
rect 317137 49811 317203 49814
rect 320081 49811 320147 49814
rect 313181 49736 315080 49738
rect 313181 49680 313186 49736
rect 313242 49680 315080 49736
rect 313181 49678 315080 49680
rect 315254 49678 316092 49738
rect 317321 49738 317387 49741
rect 318149 49738 318215 49741
rect 317321 49736 318215 49738
rect 317321 49680 317326 49736
rect 317382 49680 318154 49736
rect 318210 49680 318215 49736
rect 317321 49678 318215 49680
rect 277209 49675 277275 49678
rect 281349 49675 281415 49678
rect 284017 49675 284083 49678
rect 289721 49675 289787 49678
rect 291009 49675 291075 49678
rect 293769 49675 293835 49678
rect 296670 49605 296730 49678
rect 300485 49675 300551 49678
rect 303521 49675 303587 49678
rect 306281 49675 306347 49678
rect 313181 49675 313247 49678
rect 275921 49600 276306 49602
rect 275921 49544 275926 49600
rect 275982 49544 276306 49600
rect 275921 49542 276306 49544
rect 296621 49600 296730 49605
rect 296621 49544 296626 49600
rect 296682 49544 296730 49600
rect 296621 49542 296730 49544
rect 314469 49602 314535 49605
rect 315254 49602 315314 49678
rect 317321 49675 317387 49678
rect 318149 49675 318215 49678
rect 319989 49738 320055 49741
rect 321093 49738 321159 49741
rect 319989 49736 321159 49738
rect 319989 49680 319994 49736
rect 320050 49680 321098 49736
rect 321154 49680 321159 49736
rect 319989 49678 321159 49680
rect 319989 49675 320055 49678
rect 321093 49675 321159 49678
rect 322841 49738 322907 49741
rect 324772 49738 324832 50048
rect 325784 49738 325844 50048
rect 326337 49874 326403 49877
rect 328502 49874 328562 50222
rect 329648 50116 329708 50222
rect 330660 50116 330720 50358
rect 331857 50282 331923 50285
rect 331857 50280 333346 50282
rect 331857 50224 331862 50280
rect 331918 50224 333346 50280
rect 331857 50222 333346 50224
rect 331857 50219 331923 50222
rect 326337 49872 328562 49874
rect 326337 49816 326342 49872
rect 326398 49816 328562 49872
rect 326337 49814 328562 49816
rect 326337 49811 326403 49814
rect 322841 49736 324832 49738
rect 322841 49680 322846 49736
rect 322902 49680 324832 49736
rect 322841 49678 324832 49680
rect 325006 49678 325844 49738
rect 326521 49738 326587 49741
rect 328636 49738 328696 50048
rect 329189 49874 329255 49877
rect 331580 49874 331640 50048
rect 329189 49872 331640 49874
rect 329189 49816 329194 49872
rect 329250 49816 331640 49872
rect 329189 49814 331640 49816
rect 329189 49811 329255 49814
rect 326521 49736 328696 49738
rect 326521 49680 326526 49736
rect 326582 49680 328696 49736
rect 326521 49678 328696 49680
rect 330661 49738 330727 49741
rect 332592 49738 332652 50048
rect 333286 49874 333346 50222
rect 333512 50116 333572 50494
rect 335997 50552 339460 50554
rect 335997 50496 336002 50552
rect 336058 50496 339460 50552
rect 335997 50494 339460 50496
rect 335997 50491 336063 50494
rect 333697 50418 333763 50421
rect 333697 50416 336516 50418
rect 333697 50360 333702 50416
rect 333758 50360 336516 50416
rect 333697 50358 336516 50360
rect 333697 50355 333763 50358
rect 334709 50282 334775 50285
rect 334709 50280 336290 50282
rect 334709 50224 334714 50280
rect 334770 50224 336290 50280
rect 334709 50222 336290 50224
rect 334709 50219 334775 50222
rect 334524 49874 334584 50048
rect 333286 49814 334584 49874
rect 330661 49736 332652 49738
rect 330661 49680 330666 49736
rect 330722 49680 332652 49736
rect 330661 49678 332652 49680
rect 333421 49738 333487 49741
rect 335444 49738 335504 50048
rect 336230 49874 336290 50222
rect 336456 50116 336516 50358
rect 339400 50116 339460 50494
rect 341332 50552 343699 50554
rect 341332 50496 343638 50552
rect 343694 50496 343699 50552
rect 341332 50494 343699 50496
rect 341332 50116 341392 50494
rect 343633 50491 343699 50494
rect 353016 50552 354739 50554
rect 353016 50496 354678 50552
rect 354734 50496 354739 50552
rect 353016 50494 354739 50496
rect 345197 50418 345263 50421
rect 342344 50416 345263 50418
rect 342344 50360 345202 50416
rect 345258 50360 345263 50416
rect 342344 50358 345263 50360
rect 342344 50116 342404 50358
rect 345197 50355 345263 50358
rect 346485 50282 346551 50285
rect 351913 50282 351979 50285
rect 345798 50280 346551 50282
rect 345798 50224 346490 50280
rect 346546 50224 346551 50280
rect 345798 50222 346551 50224
rect 337468 49874 337528 50048
rect 336230 49814 337528 49874
rect 333421 49736 335504 49738
rect 333421 49680 333426 49736
rect 333482 49680 335504 49736
rect 333421 49678 335504 49680
rect 336181 49738 336247 49741
rect 338388 49738 338448 50048
rect 336181 49736 338448 49738
rect 336181 49680 336186 49736
rect 336242 49680 338448 49736
rect 336181 49678 338448 49680
rect 340320 49738 340380 50048
rect 342253 49738 342319 49741
rect 340320 49736 342319 49738
rect 340320 49680 342258 49736
rect 342314 49680 342319 49736
rect 340320 49678 342319 49680
rect 343264 49738 343324 50048
rect 344276 49874 344336 50048
rect 345013 50010 345079 50013
rect 345196 50010 345256 50048
rect 345013 50008 345256 50010
rect 345013 49952 345018 50008
rect 345074 49952 345256 50008
rect 345013 49950 345256 49952
rect 345013 49947 345079 49950
rect 345798 49874 345858 50222
rect 346485 50219 346551 50222
rect 349152 50280 351979 50282
rect 349152 50224 351918 50280
rect 351974 50224 351979 50280
rect 349152 50222 351979 50224
rect 349152 50116 349212 50222
rect 351913 50219 351979 50222
rect 353016 50116 353076 50494
rect 354673 50491 354739 50494
rect 356053 50418 356119 50421
rect 353936 50416 356119 50418
rect 353936 50360 356058 50416
rect 356114 50360 356119 50416
rect 353936 50358 356119 50360
rect 353936 50116 353996 50358
rect 356053 50355 356119 50358
rect 357709 50282 357775 50285
rect 360193 50282 360259 50285
rect 354948 50280 357775 50282
rect 354948 50224 357714 50280
rect 357770 50224 357775 50280
rect 354948 50222 357775 50224
rect 354948 50116 355008 50222
rect 357709 50219 357775 50222
rect 357892 50280 360259 50282
rect 357892 50224 360198 50280
rect 360254 50224 360259 50280
rect 357892 50222 360259 50224
rect 357892 50116 357952 50222
rect 360193 50219 360259 50222
rect 360836 50116 360896 50630
rect 363045 50627 363111 50630
rect 407990 50688 410583 50690
rect 407990 50632 410522 50688
rect 410578 50632 410583 50688
rect 407990 50630 410583 50632
rect 364609 50554 364675 50557
rect 382273 50554 382339 50557
rect 398925 50554 398991 50557
rect 362768 50552 364675 50554
rect 362768 50496 364614 50552
rect 364670 50496 364675 50552
rect 362768 50494 364675 50496
rect 362768 50116 362828 50494
rect 364609 50491 364675 50494
rect 380248 50552 382339 50554
rect 380248 50496 382278 50552
rect 382334 50496 382339 50552
rect 380248 50494 382339 50496
rect 365713 50418 365779 50421
rect 374361 50418 374427 50421
rect 363688 50416 365779 50418
rect 363688 50360 365718 50416
rect 365774 50360 365779 50416
rect 363688 50358 365779 50360
rect 363688 50116 363748 50358
rect 365713 50355 365779 50358
rect 371508 50416 374427 50418
rect 371508 50360 374366 50416
rect 374422 50360 374427 50416
rect 371508 50358 374427 50360
rect 367277 50282 367343 50285
rect 369945 50282 370011 50285
rect 364700 50280 367343 50282
rect 364700 50224 367282 50280
rect 367338 50224 367343 50280
rect 364700 50222 367343 50224
rect 364700 50116 364760 50222
rect 367277 50219 367343 50222
rect 367644 50280 370011 50282
rect 367644 50224 369950 50280
rect 370006 50224 370011 50280
rect 367644 50222 370011 50224
rect 367644 50116 367704 50222
rect 369945 50219 370011 50222
rect 371508 50116 371568 50358
rect 374361 50355 374427 50358
rect 376845 50282 376911 50285
rect 379513 50282 379579 50285
rect 374452 50280 376911 50282
rect 374452 50224 376850 50280
rect 376906 50224 376911 50280
rect 374452 50222 376911 50224
rect 374452 50116 374512 50222
rect 376845 50219 376911 50222
rect 377304 50280 379579 50282
rect 377304 50224 379518 50280
rect 379574 50224 379579 50280
rect 377304 50222 379579 50224
rect 377304 50116 377364 50222
rect 379513 50219 379579 50222
rect 380248 50116 380308 50494
rect 382273 50491 382339 50494
rect 396808 50552 398991 50554
rect 396808 50496 398930 50552
rect 398986 50496 398991 50552
rect 396808 50494 398991 50496
rect 383745 50418 383811 50421
rect 385033 50418 385099 50421
rect 387977 50418 388043 50421
rect 393405 50418 393471 50421
rect 395061 50418 395127 50421
rect 382180 50416 383811 50418
rect 382180 50360 383750 50416
rect 383806 50360 383811 50416
rect 382180 50358 383811 50360
rect 382180 50116 382240 50358
rect 383745 50355 383811 50358
rect 383886 50416 385099 50418
rect 383886 50360 385038 50416
rect 385094 50360 385099 50416
rect 383886 50358 385099 50360
rect 383886 50282 383946 50358
rect 385033 50355 385099 50358
rect 386646 50416 388043 50418
rect 386646 50360 387982 50416
rect 388038 50360 388043 50416
rect 386646 50358 388043 50360
rect 386505 50282 386571 50285
rect 383192 50222 383946 50282
rect 384112 50280 386571 50282
rect 384112 50224 386510 50280
rect 386566 50224 386571 50280
rect 384112 50222 386571 50224
rect 383192 50116 383252 50222
rect 384112 50116 384172 50222
rect 386505 50219 386571 50222
rect 386646 50146 386706 50358
rect 387977 50355 388043 50358
rect 391012 50416 393471 50418
rect 391012 50360 393410 50416
rect 393466 50360 393471 50416
rect 391012 50358 393471 50360
rect 389173 50282 389239 50285
rect 386166 50086 386706 50146
rect 387056 50280 389239 50282
rect 387056 50224 389178 50280
rect 389234 50224 389239 50280
rect 387056 50222 389239 50224
rect 387056 50116 387116 50222
rect 389173 50219 389239 50222
rect 391012 50116 391072 50358
rect 393405 50355 393471 50358
rect 393638 50416 395127 50418
rect 393638 50360 395066 50416
rect 395122 50360 395127 50416
rect 393638 50358 395127 50360
rect 391932 50222 393146 50282
rect 391932 50116 391992 50222
rect 368749 50078 368815 50081
rect 368594 50076 368815 50078
rect 344276 49814 345858 49874
rect 345105 49738 345171 49741
rect 343264 49736 345171 49738
rect 343264 49680 345110 49736
rect 345166 49680 345171 49736
rect 343264 49678 345171 49680
rect 346208 49738 346268 50048
rect 346393 49874 346459 49877
rect 347128 49874 347188 50048
rect 346393 49872 347188 49874
rect 346393 49816 346398 49872
rect 346454 49816 347188 49872
rect 346393 49814 347188 49816
rect 346393 49811 346459 49814
rect 348140 49741 348200 50048
rect 347957 49738 348023 49741
rect 346208 49736 348023 49738
rect 346208 49680 347962 49736
rect 348018 49680 348023 49736
rect 346208 49678 348023 49680
rect 348140 49736 348207 49741
rect 348140 49680 348146 49736
rect 348202 49680 348207 49736
rect 348140 49678 348207 49680
rect 350072 49738 350132 50048
rect 351084 49874 351144 50048
rect 351821 49874 351887 49877
rect 351084 49872 351887 49874
rect 351084 49816 351826 49872
rect 351882 49816 351887 49872
rect 351084 49814 351887 49816
rect 352004 49874 352064 50048
rect 354857 49874 354923 49877
rect 352004 49872 354923 49874
rect 352004 49816 354862 49872
rect 354918 49816 354923 49872
rect 352004 49814 354923 49816
rect 351821 49811 351887 49814
rect 354857 49811 354923 49814
rect 352189 49738 352255 49741
rect 350072 49736 352255 49738
rect 350072 49680 352194 49736
rect 352250 49680 352255 49736
rect 350072 49678 352255 49680
rect 355960 49738 356020 50048
rect 356880 49874 356940 50048
rect 358812 50010 358872 50048
rect 359824 50010 359884 50048
rect 360653 50010 360719 50013
rect 358812 49950 359106 50010
rect 359824 50008 360719 50010
rect 359824 49952 360658 50008
rect 360714 49952 360719 50008
rect 359824 49950 360719 49952
rect 358905 49874 358971 49877
rect 356880 49872 358971 49874
rect 356880 49816 358910 49872
rect 358966 49816 358971 49872
rect 356880 49814 358971 49816
rect 359046 49874 359106 49950
rect 360653 49947 360719 49950
rect 361573 49874 361639 49877
rect 359046 49872 361639 49874
rect 359046 49816 361578 49872
rect 361634 49816 361639 49872
rect 359046 49814 361639 49816
rect 361756 49874 361816 50048
rect 364425 49874 364491 49877
rect 361756 49872 364491 49874
rect 361756 49816 364430 49872
rect 364486 49816 364491 49872
rect 361756 49814 364491 49816
rect 358905 49811 358971 49814
rect 361573 49811 361639 49814
rect 364425 49811 364491 49814
rect 357525 49738 357591 49741
rect 355960 49736 357591 49738
rect 355960 49680 357530 49736
rect 357586 49680 357591 49736
rect 355960 49678 357591 49680
rect 322841 49675 322907 49678
rect 314469 49600 315314 49602
rect 314469 49544 314474 49600
rect 314530 49544 315314 49600
rect 314469 49542 315314 49544
rect 323945 49602 324011 49605
rect 325006 49602 325066 49678
rect 326521 49675 326587 49678
rect 330661 49675 330727 49678
rect 333421 49675 333487 49678
rect 336181 49675 336247 49678
rect 342253 49675 342319 49678
rect 345105 49675 345171 49678
rect 347957 49675 348023 49678
rect 348141 49675 348207 49678
rect 352189 49675 352255 49678
rect 357525 49675 357591 49678
rect 360653 49738 360719 49741
rect 361573 49738 361639 49741
rect 360653 49736 361639 49738
rect 360653 49680 360658 49736
rect 360714 49680 361578 49736
rect 361634 49680 361639 49736
rect 360653 49678 361639 49680
rect 365620 49738 365680 50048
rect 366632 49874 366692 50048
rect 368594 50020 368754 50076
rect 368810 50020 368815 50076
rect 368594 50018 368815 50020
rect 368749 50015 368815 50018
rect 368473 49874 368539 49877
rect 366632 49872 368539 49874
rect 366632 49816 368478 49872
rect 368534 49816 368539 49872
rect 366632 49814 368539 49816
rect 368473 49811 368539 49814
rect 367093 49738 367159 49741
rect 365620 49736 367159 49738
rect 365620 49680 367098 49736
rect 367154 49680 367159 49736
rect 365620 49678 367159 49680
rect 369576 49738 369636 50048
rect 369853 49874 369919 49877
rect 370496 49874 370556 50048
rect 369853 49872 370556 49874
rect 369853 49816 369858 49872
rect 369914 49816 370556 49872
rect 369853 49814 370556 49816
rect 369853 49811 369919 49814
rect 371417 49738 371483 49741
rect 369576 49736 371483 49738
rect 369576 49680 371422 49736
rect 371478 49680 371483 49736
rect 369576 49678 371483 49680
rect 372520 49738 372580 50048
rect 373440 49874 373500 50048
rect 375189 49874 375255 49877
rect 373440 49872 375255 49874
rect 373440 49816 375194 49872
rect 375250 49816 375255 49872
rect 373440 49814 375255 49816
rect 375189 49811 375255 49814
rect 375372 49741 375432 50048
rect 374177 49738 374243 49741
rect 372520 49736 374243 49738
rect 372520 49680 374182 49736
rect 374238 49680 374243 49736
rect 372520 49678 374243 49680
rect 375372 49736 375439 49741
rect 375372 49680 375378 49736
rect 375434 49680 375439 49736
rect 375372 49678 375439 49680
rect 376384 49738 376444 50048
rect 378316 49874 378376 50048
rect 379328 50010 379388 50048
rect 380065 50010 380131 50013
rect 379328 50008 380131 50010
rect 379328 49952 380070 50008
rect 380126 49952 380131 50008
rect 379328 49950 380131 49952
rect 380065 49947 380131 49950
rect 380893 49874 380959 49877
rect 378316 49872 380959 49874
rect 378316 49816 380898 49872
rect 380954 49816 380959 49872
rect 378316 49814 380959 49816
rect 381260 49874 381320 50048
rect 383929 49874 383995 49877
rect 381260 49872 383995 49874
rect 381260 49816 383934 49872
rect 383990 49816 383995 49872
rect 381260 49814 383995 49816
rect 385124 49874 385184 50048
rect 387793 50010 387859 50013
rect 388068 50010 388128 50048
rect 387793 50008 388128 50010
rect 387793 49952 387798 50008
rect 387854 49952 388128 50008
rect 387793 49950 388128 49952
rect 387793 49947 387859 49950
rect 388161 49874 388227 49877
rect 385124 49872 388227 49874
rect 385124 49816 388166 49872
rect 388222 49816 388227 49872
rect 385124 49814 388227 49816
rect 380893 49811 380959 49814
rect 383929 49811 383995 49814
rect 388161 49811 388227 49814
rect 378317 49738 378383 49741
rect 376384 49736 378383 49738
rect 376384 49680 378322 49736
rect 378378 49680 378383 49736
rect 376384 49678 378383 49680
rect 360653 49675 360719 49678
rect 361573 49675 361639 49678
rect 367093 49675 367159 49678
rect 371417 49675 371483 49678
rect 374177 49675 374243 49678
rect 375373 49675 375439 49678
rect 378317 49675 378383 49678
rect 380065 49738 380131 49741
rect 381077 49738 381143 49741
rect 380065 49736 381143 49738
rect 380065 49680 380070 49736
rect 380126 49680 381082 49736
rect 381138 49680 381143 49736
rect 380065 49678 381143 49680
rect 388988 49738 389048 50048
rect 390000 49874 390060 50048
rect 391933 49874 391999 49877
rect 390000 49872 391999 49874
rect 390000 49816 391938 49872
rect 391994 49816 391999 49872
rect 390000 49814 391999 49816
rect 391933 49811 391999 49814
rect 390737 49738 390803 49741
rect 388988 49736 390803 49738
rect 388988 49680 390742 49736
rect 390798 49680 390803 49736
rect 388988 49678 390803 49680
rect 392944 49738 393004 50048
rect 393086 49874 393146 50222
rect 393638 49874 393698 50358
rect 395061 50355 395127 50358
rect 396165 50282 396231 50285
rect 393864 50280 396231 50282
rect 393864 50224 396170 50280
rect 396226 50224 396231 50280
rect 393864 50222 396231 50224
rect 393864 50116 393924 50222
rect 396165 50219 396231 50222
rect 396808 50116 396868 50494
rect 398925 50491 398991 50494
rect 400489 50418 400555 50421
rect 397820 50416 400555 50418
rect 397820 50360 400494 50416
rect 400550 50360 400555 50416
rect 397820 50358 400555 50360
rect 397820 50116 397880 50358
rect 400489 50355 400555 50358
rect 403065 50282 403131 50285
rect 404537 50282 404603 50285
rect 407757 50282 407823 50285
rect 400672 50280 403131 50282
rect 400672 50224 403070 50280
rect 403126 50224 403131 50280
rect 400672 50222 403131 50224
rect 400672 50116 400732 50222
rect 403065 50219 403131 50222
rect 403206 50280 404603 50282
rect 403206 50224 404542 50280
rect 404598 50224 404603 50280
rect 403206 50222 404603 50224
rect 403206 50146 403266 50222
rect 404537 50219 404603 50222
rect 405548 50280 407823 50282
rect 405548 50224 407762 50280
rect 407818 50224 407823 50280
rect 405548 50222 407823 50224
rect 402726 50086 403266 50146
rect 405548 50116 405608 50222
rect 407757 50219 407823 50222
rect 407990 50146 408050 50630
rect 410517 50627 410583 50630
rect 421741 50690 421807 50693
rect 424501 50690 424567 50693
rect 421741 50688 424567 50690
rect 421741 50632 421746 50688
rect 421802 50632 424506 50688
rect 424562 50632 424567 50688
rect 421741 50630 424567 50632
rect 421741 50627 421807 50630
rect 424501 50627 424567 50630
rect 431309 50690 431375 50693
rect 434621 50690 434687 50693
rect 431309 50688 434687 50690
rect 431309 50632 431314 50688
rect 431370 50632 434626 50688
rect 434682 50632 434687 50688
rect 431309 50630 434687 50632
rect 431309 50627 431375 50630
rect 434621 50627 434687 50630
rect 412081 50554 412147 50557
rect 427077 50554 427143 50557
rect 407510 50086 408050 50146
rect 408492 50552 412147 50554
rect 408492 50496 412086 50552
rect 412142 50496 412147 50552
rect 408492 50494 412147 50496
rect 408492 50116 408552 50494
rect 412081 50491 412147 50494
rect 424040 50552 427143 50554
rect 424040 50496 427082 50552
rect 427138 50496 427143 50552
rect 424040 50494 427143 50496
rect 416681 50418 416747 50421
rect 420177 50418 420243 50421
rect 413878 50416 416747 50418
rect 413878 50360 416686 50416
rect 416742 50360 416747 50416
rect 413878 50358 416747 50360
rect 413277 50282 413343 50285
rect 410424 50280 413343 50282
rect 410424 50224 413282 50280
rect 413338 50224 413343 50280
rect 410424 50222 413343 50224
rect 410424 50116 410484 50222
rect 413277 50219 413343 50222
rect 413878 50146 413938 50358
rect 416681 50355 416747 50358
rect 417742 50416 420243 50418
rect 417742 50360 420182 50416
rect 420238 50360 420243 50416
rect 417742 50358 420243 50360
rect 417417 50282 417483 50285
rect 413398 50086 413938 50146
rect 414288 50280 417483 50282
rect 414288 50224 417422 50280
rect 417478 50224 417483 50280
rect 414288 50222 417483 50224
rect 414288 50116 414348 50222
rect 417417 50219 417483 50222
rect 417742 50146 417802 50358
rect 420177 50355 420243 50358
rect 421054 50358 422310 50418
rect 421054 50282 421114 50358
rect 417262 50086 417802 50146
rect 418244 50222 419458 50282
rect 418244 50116 418304 50222
rect 394693 49874 394759 49877
rect 393086 49814 393698 49874
rect 394006 49872 394759 49874
rect 394006 49816 394698 49872
rect 394754 49816 394759 49872
rect 394006 49814 394759 49816
rect 394006 49738 394066 49814
rect 394693 49811 394759 49814
rect 392944 49678 394066 49738
rect 394693 49738 394759 49741
rect 394876 49738 394936 50048
rect 394693 49736 394936 49738
rect 394693 49680 394698 49736
rect 394754 49680 394936 49736
rect 394693 49678 394936 49680
rect 395796 49738 395856 50048
rect 397453 49738 397519 49741
rect 395796 49736 397519 49738
rect 395796 49680 397458 49736
rect 397514 49680 397519 49736
rect 395796 49678 397519 49680
rect 398740 49738 398800 50048
rect 399752 49874 399812 50048
rect 401684 49874 401744 50048
rect 402973 49874 403039 49877
rect 399752 49814 400506 49874
rect 401684 49872 403039 49874
rect 401684 49816 402978 49872
rect 403034 49816 403039 49872
rect 401684 49814 403039 49816
rect 400305 49738 400371 49741
rect 398740 49736 400371 49738
rect 398740 49680 400310 49736
rect 400366 49680 400371 49736
rect 398740 49678 400371 49680
rect 400446 49738 400506 49814
rect 402973 49811 403039 49814
rect 401685 49738 401751 49741
rect 400446 49736 401751 49738
rect 400446 49680 401690 49736
rect 401746 49680 401751 49736
rect 400446 49678 401751 49680
rect 403616 49738 403676 50048
rect 404628 49874 404688 50048
rect 406560 50010 406620 50048
rect 406560 49950 407314 50010
rect 407113 49874 407179 49877
rect 404628 49872 407179 49874
rect 404628 49816 407118 49872
rect 407174 49816 407179 49872
rect 404628 49814 407179 49816
rect 407254 49874 407314 49950
rect 409137 49874 409203 49877
rect 407254 49872 409203 49874
rect 407254 49816 409142 49872
rect 409198 49816 409203 49872
rect 407254 49814 409203 49816
rect 407113 49811 407179 49814
rect 409137 49811 409203 49814
rect 405825 49738 405891 49741
rect 403616 49736 405891 49738
rect 403616 49680 405830 49736
rect 405886 49680 405891 49736
rect 403616 49678 405891 49680
rect 409504 49738 409564 50048
rect 411436 49874 411496 50048
rect 412356 50010 412416 50048
rect 412541 50010 412607 50013
rect 412356 50008 412607 50010
rect 412356 49952 412546 50008
rect 412602 49952 412607 50008
rect 412356 49950 412607 49952
rect 412541 49947 412607 49950
rect 414841 49874 414907 49877
rect 411436 49872 414907 49874
rect 411436 49816 414846 49872
rect 414902 49816 414907 49872
rect 411436 49814 414907 49816
rect 414841 49811 414907 49814
rect 411897 49738 411963 49741
rect 409504 49736 411963 49738
rect 409504 49680 411902 49736
rect 411958 49680 411963 49736
rect 409504 49678 411963 49680
rect 380065 49675 380131 49678
rect 381077 49675 381143 49678
rect 390737 49675 390803 49678
rect 394693 49675 394759 49678
rect 397453 49675 397519 49678
rect 400305 49675 400371 49678
rect 401685 49675 401751 49678
rect 405825 49675 405891 49678
rect 411897 49675 411963 49678
rect 412541 49738 412607 49741
rect 414657 49738 414723 49741
rect 412541 49736 414723 49738
rect 412541 49680 412546 49736
rect 412602 49680 414662 49736
rect 414718 49680 414723 49736
rect 412541 49678 414723 49680
rect 415300 49738 415360 50048
rect 416312 49874 416372 50048
rect 418797 49874 418863 49877
rect 416312 49872 418863 49874
rect 416312 49816 418802 49872
rect 418858 49816 418863 49872
rect 416312 49814 418863 49816
rect 418797 49811 418863 49814
rect 417601 49738 417667 49741
rect 415300 49736 417667 49738
rect 415300 49680 417606 49736
rect 417662 49680 417667 49736
rect 415300 49678 417667 49680
rect 419164 49738 419224 50048
rect 419398 49874 419458 50222
rect 420176 50222 421114 50282
rect 422250 50282 422310 50358
rect 422937 50282 423003 50285
rect 422250 50280 423003 50282
rect 422250 50224 422942 50280
rect 422998 50224 423003 50280
rect 422250 50222 423003 50224
rect 420176 50116 420236 50222
rect 422937 50219 423003 50222
rect 421741 50146 421807 50149
rect 421218 50144 421807 50146
rect 421218 50088 421746 50144
rect 421802 50088 421807 50144
rect 424040 50116 424100 50494
rect 427077 50491 427143 50494
rect 428457 50418 428523 50421
rect 432597 50418 432663 50421
rect 441061 50418 441127 50421
rect 445661 50418 445727 50421
rect 425052 50416 428523 50418
rect 425052 50360 428462 50416
rect 428518 50360 428523 50416
rect 425052 50358 428523 50360
rect 425052 50116 425112 50358
rect 428457 50355 428523 50358
rect 429928 50416 432663 50418
rect 429928 50360 432602 50416
rect 432658 50360 432663 50416
rect 429928 50358 432663 50360
rect 429745 50282 429811 50285
rect 426984 50280 429811 50282
rect 426984 50224 429750 50280
rect 429806 50224 429811 50280
rect 426984 50222 429811 50224
rect 426984 50116 427044 50222
rect 429745 50219 429811 50222
rect 429928 50116 429988 50358
rect 432597 50355 432663 50358
rect 438668 50416 441127 50418
rect 438668 50360 441066 50416
rect 441122 50360 441127 50416
rect 438668 50358 441127 50360
rect 433977 50282 434043 50285
rect 438117 50282 438183 50285
rect 431910 50280 434043 50282
rect 431910 50224 433982 50280
rect 434038 50224 434043 50280
rect 431910 50222 434043 50224
rect 431309 50146 431375 50149
rect 430878 50144 431375 50146
rect 421218 50086 421807 50088
rect 430878 50088 431314 50144
rect 431370 50088 431375 50144
rect 430878 50086 431375 50088
rect 421741 50083 421807 50086
rect 431309 50083 431375 50086
rect 431910 50048 431970 50222
rect 433977 50219 434043 50222
rect 434804 50280 438183 50282
rect 434804 50224 438122 50280
rect 438178 50224 438183 50280
rect 434804 50222 438183 50224
rect 434804 50116 434864 50222
rect 438117 50219 438183 50222
rect 438668 50116 438728 50358
rect 441061 50355 441127 50358
rect 441612 50416 445727 50418
rect 441612 50360 445666 50416
rect 445722 50360 445727 50416
rect 441612 50358 445727 50360
rect 439680 50222 440802 50282
rect 439680 50116 439740 50222
rect 421557 49874 421623 49877
rect 419398 49872 421623 49874
rect 419398 49816 421562 49872
rect 421618 49816 421623 49872
rect 419398 49814 421623 49816
rect 421557 49811 421623 49814
rect 421741 49738 421807 49741
rect 419164 49736 421807 49738
rect 419164 49680 421746 49736
rect 421802 49680 421807 49736
rect 419164 49678 421807 49680
rect 422108 49738 422168 50048
rect 423120 49738 423180 50048
rect 425697 49738 425763 49741
rect 422108 49678 422954 49738
rect 423120 49736 425763 49738
rect 423120 49680 425702 49736
rect 425758 49680 425763 49736
rect 423120 49678 425763 49680
rect 425972 49738 426032 50048
rect 427996 49874 428056 50048
rect 428916 50010 428976 50048
rect 429653 50010 429719 50013
rect 428916 50008 429719 50010
rect 428916 49952 429658 50008
rect 429714 49952 429719 50008
rect 428916 49950 429719 49952
rect 429653 49947 429719 49950
rect 431401 49874 431467 49877
rect 427996 49872 431467 49874
rect 427996 49816 431406 49872
rect 431462 49816 431467 49872
rect 427996 49814 431467 49816
rect 431401 49811 431467 49814
rect 428641 49738 428707 49741
rect 425972 49736 428707 49738
rect 425972 49680 428646 49736
rect 428702 49680 428707 49736
rect 425972 49678 428707 49680
rect 412541 49675 412607 49678
rect 414657 49675 414723 49678
rect 417601 49675 417667 49678
rect 421741 49675 421807 49678
rect 323945 49600 325066 49602
rect 323945 49544 323950 49600
rect 324006 49544 325066 49600
rect 323945 49542 325066 49544
rect 422894 49602 422954 49678
rect 425697 49675 425763 49678
rect 428641 49675 428707 49678
rect 429653 49738 429719 49741
rect 431217 49738 431283 49741
rect 429653 49736 431283 49738
rect 429653 49680 429658 49736
rect 429714 49680 431222 49736
rect 431278 49680 431283 49736
rect 429653 49678 431283 49680
rect 431860 49678 431970 50048
rect 432872 49738 432932 50048
rect 433792 49874 433852 50048
rect 435724 50010 435784 50048
rect 436461 50010 436527 50013
rect 435724 50008 436527 50010
rect 435724 49952 436466 50008
rect 436522 49952 436527 50008
rect 435724 49950 436527 49952
rect 436461 49947 436527 49950
rect 436553 49874 436619 49877
rect 433792 49872 436619 49874
rect 433792 49816 436558 49872
rect 436614 49816 436619 49872
rect 433792 49814 436619 49816
rect 436553 49811 436619 49814
rect 435357 49738 435423 49741
rect 432872 49736 435423 49738
rect 432872 49680 435362 49736
rect 435418 49680 435423 49736
rect 432872 49678 435423 49680
rect 436736 49738 436796 50048
rect 437656 49874 437716 50048
rect 440417 49874 440483 49877
rect 437656 49872 440483 49874
rect 437656 49816 440422 49872
rect 440478 49816 440483 49872
rect 437656 49814 440483 49816
rect 440417 49811 440483 49814
rect 439497 49738 439563 49741
rect 436736 49736 439563 49738
rect 436736 49680 439502 49736
rect 439558 49680 439563 49736
rect 436736 49678 439563 49680
rect 440600 49738 440660 50048
rect 440742 49874 440802 50222
rect 441612 50116 441672 50358
rect 445661 50355 445727 50358
rect 446305 50282 446371 50285
rect 443544 50280 446371 50282
rect 443544 50224 446310 50280
rect 446366 50224 446371 50280
rect 443544 50222 446371 50224
rect 443544 50116 443604 50222
rect 446305 50219 446371 50222
rect 446488 50116 446548 50766
rect 449157 50763 449223 50766
rect 450537 50690 450603 50693
rect 461025 50690 461091 50693
rect 498285 50690 498351 50693
rect 545205 50690 545271 50693
rect 447408 50688 450603 50690
rect 447408 50632 450542 50688
rect 450598 50632 450603 50688
rect 447408 50630 450603 50632
rect 447408 50116 447468 50630
rect 450537 50627 450603 50630
rect 458172 50688 461091 50690
rect 458172 50632 461030 50688
rect 461086 50632 461091 50688
rect 458172 50630 461091 50632
rect 453297 50554 453363 50557
rect 450352 50552 453363 50554
rect 450352 50496 453302 50552
rect 453358 50496 453363 50552
rect 450352 50494 453363 50496
rect 450352 50116 450412 50494
rect 453297 50491 453363 50494
rect 454677 50418 454743 50421
rect 451364 50416 454743 50418
rect 451364 50360 454682 50416
rect 454738 50360 454743 50416
rect 451364 50358 454743 50360
rect 451364 50116 451424 50358
rect 454677 50355 454743 50358
rect 456977 50282 457043 50285
rect 454216 50280 457043 50282
rect 454216 50224 456982 50280
rect 457038 50224 457043 50280
rect 454216 50222 457043 50224
rect 454216 50116 454276 50222
rect 456977 50219 457043 50222
rect 458172 50116 458232 50630
rect 461025 50627 461091 50630
rect 496076 50688 498351 50690
rect 496076 50632 498290 50688
rect 498346 50632 498351 50688
rect 496076 50630 498351 50632
rect 462405 50554 462471 50557
rect 491293 50554 491359 50557
rect 460104 50552 462471 50554
rect 460104 50496 462410 50552
rect 462466 50496 462471 50552
rect 460104 50494 462471 50496
rect 460104 50116 460164 50494
rect 462405 50491 462471 50494
rect 489268 50552 491359 50554
rect 489268 50496 491298 50552
rect 491354 50496 491359 50552
rect 489268 50494 491359 50496
rect 463785 50418 463851 50421
rect 466545 50418 466611 50421
rect 470685 50418 470751 50421
rect 461024 50416 463851 50418
rect 461024 50360 463790 50416
rect 463846 50360 463851 50416
rect 461024 50358 463851 50360
rect 461024 50116 461084 50358
rect 463785 50355 463851 50358
rect 465582 50416 466611 50418
rect 465582 50360 466550 50416
rect 466606 50360 466611 50416
rect 465582 50358 466611 50360
rect 465165 50282 465231 50285
rect 463048 50280 465231 50282
rect 463048 50224 465170 50280
rect 465226 50224 465231 50280
rect 463048 50222 465231 50224
rect 463048 50116 463108 50222
rect 465165 50219 465231 50222
rect 465582 50146 465642 50358
rect 466545 50355 466611 50358
rect 467832 50416 470751 50418
rect 467832 50360 470690 50416
rect 470746 50360 470751 50416
rect 467832 50358 470751 50360
rect 467649 50282 467715 50285
rect 465010 50086 465642 50146
rect 465900 50280 467715 50282
rect 465900 50224 467654 50280
rect 467710 50224 467715 50280
rect 465900 50222 467715 50224
rect 465900 50116 465960 50222
rect 467649 50219 467715 50222
rect 467832 50116 467892 50358
rect 470685 50355 470751 50358
rect 470961 50418 471027 50421
rect 473353 50418 473419 50421
rect 476481 50418 476547 50421
rect 478873 50418 478939 50421
rect 483289 50418 483355 50421
rect 488533 50418 488599 50421
rect 470961 50416 473419 50418
rect 470961 50360 470966 50416
rect 471022 50360 473358 50416
rect 473414 50360 473419 50416
rect 470961 50358 473419 50360
rect 470961 50355 471027 50358
rect 473353 50355 473419 50358
rect 473720 50416 476547 50418
rect 473720 50360 476486 50416
rect 476542 50360 476547 50416
rect 473720 50358 476547 50360
rect 471973 50282 472039 50285
rect 469856 50280 472039 50282
rect 469856 50224 471978 50280
rect 472034 50224 472039 50280
rect 469856 50222 472039 50224
rect 469856 50116 469916 50222
rect 471973 50219 472039 50222
rect 470961 50146 471027 50149
rect 470806 50144 471027 50146
rect 470806 50088 470966 50144
rect 471022 50088 471027 50144
rect 473720 50116 473780 50358
rect 476481 50355 476547 50358
rect 476664 50416 478939 50418
rect 476664 50360 478878 50416
rect 478934 50360 478939 50416
rect 476664 50358 478939 50360
rect 476664 50116 476724 50358
rect 478873 50355 478939 50358
rect 480528 50416 483355 50418
rect 480528 50360 483294 50416
rect 483350 50360 483355 50416
rect 480528 50358 483355 50360
rect 480345 50282 480411 50285
rect 478596 50280 480411 50282
rect 478596 50224 480350 50280
rect 480406 50224 480411 50280
rect 478596 50222 480411 50224
rect 478596 50116 478656 50222
rect 480345 50219 480411 50222
rect 480528 50116 480588 50358
rect 483289 50355 483355 50358
rect 486324 50416 488599 50418
rect 486324 50360 488538 50416
rect 488594 50360 488599 50416
rect 486324 50358 488599 50360
rect 484301 50282 484367 50285
rect 482460 50280 484367 50282
rect 482460 50224 484306 50280
rect 484362 50224 484367 50280
rect 482460 50222 484367 50224
rect 482460 50116 482520 50222
rect 484301 50219 484367 50222
rect 486324 50116 486384 50358
rect 488533 50355 488599 50358
rect 487336 50222 488642 50282
rect 487336 50116 487396 50222
rect 470806 50086 471027 50088
rect 470961 50083 471027 50086
rect 442257 49874 442323 49877
rect 440742 49872 442323 49874
rect 440742 49816 442262 49872
rect 442318 49816 442323 49872
rect 440742 49814 442323 49816
rect 442257 49811 442323 49814
rect 442532 49738 442592 50048
rect 444464 49874 444524 50048
rect 445476 50010 445536 50048
rect 446213 50010 446279 50013
rect 445476 50008 446279 50010
rect 445476 49952 446218 50008
rect 446274 49952 446279 50008
rect 445476 49950 446279 49952
rect 446213 49947 446279 49950
rect 447961 49874 448027 49877
rect 444464 49872 448027 49874
rect 444464 49816 447966 49872
rect 448022 49816 448027 49872
rect 444464 49814 448027 49816
rect 447961 49811 448027 49814
rect 445017 49738 445083 49741
rect 440600 49678 442458 49738
rect 442532 49736 445083 49738
rect 442532 49680 445022 49736
rect 445078 49680 445083 49736
rect 442532 49678 445083 49680
rect 429653 49675 429719 49678
rect 431217 49675 431283 49678
rect 435357 49675 435423 49678
rect 439497 49675 439563 49678
rect 424317 49602 424383 49605
rect 422894 49600 424383 49602
rect 422894 49544 424322 49600
rect 424378 49544 424383 49600
rect 422894 49542 424383 49544
rect 442398 49602 442458 49678
rect 445017 49675 445083 49678
rect 446213 49738 446279 49741
rect 447777 49738 447843 49741
rect 446213 49736 447843 49738
rect 446213 49680 446218 49736
rect 446274 49680 447782 49736
rect 447838 49680 447843 49736
rect 446213 49678 447843 49680
rect 448420 49738 448480 50048
rect 449340 49874 449400 50048
rect 451917 49874 451983 49877
rect 449340 49872 451983 49874
rect 449340 49816 451922 49872
rect 451978 49816 451983 49872
rect 449340 49814 451983 49816
rect 451917 49811 451983 49814
rect 450721 49738 450787 49741
rect 448420 49736 450787 49738
rect 448420 49680 450726 49736
rect 450782 49680 450787 49736
rect 448420 49678 450787 49680
rect 452284 49738 452344 50048
rect 453296 49874 453356 50048
rect 454401 50010 454467 50013
rect 455228 50010 455288 50048
rect 454401 50008 455288 50010
rect 454401 49952 454406 50008
rect 454462 49952 455288 50008
rect 454401 49950 455288 49952
rect 454401 49947 454467 49950
rect 455505 49874 455571 49877
rect 453296 49872 455571 49874
rect 453296 49816 455510 49872
rect 455566 49816 455571 49872
rect 453296 49814 455571 49816
rect 455505 49811 455571 49814
rect 454033 49738 454099 49741
rect 452284 49736 454099 49738
rect 452284 49680 454038 49736
rect 454094 49680 454099 49736
rect 452284 49678 454099 49680
rect 456148 49738 456208 50048
rect 457160 49874 457220 50048
rect 459092 49874 459152 50048
rect 461209 49874 461275 49877
rect 457160 49814 458466 49874
rect 459092 49872 461275 49874
rect 459092 49816 461214 49872
rect 461270 49816 461275 49872
rect 459092 49814 461275 49816
rect 458265 49738 458331 49741
rect 456148 49736 458331 49738
rect 456148 49680 458270 49736
rect 458326 49680 458331 49736
rect 456148 49678 458331 49680
rect 458406 49738 458466 49814
rect 461209 49811 461275 49814
rect 459553 49738 459619 49741
rect 458406 49736 459619 49738
rect 458406 49680 459558 49736
rect 459614 49680 459619 49736
rect 458406 49678 459619 49680
rect 462036 49738 462096 50048
rect 463968 49874 464028 50048
rect 466729 49874 466795 49877
rect 463968 49872 466795 49874
rect 463968 49816 466734 49872
rect 466790 49816 466795 49872
rect 463968 49814 466795 49816
rect 466729 49811 466795 49814
rect 463969 49738 464035 49741
rect 462036 49736 464035 49738
rect 462036 49680 463974 49736
rect 464030 49680 464035 49736
rect 462036 49678 464035 49680
rect 466912 49738 466972 50048
rect 468844 49874 468904 50048
rect 470869 49874 470935 49877
rect 468844 49872 470935 49874
rect 468844 49816 470874 49872
rect 470930 49816 470935 49872
rect 468844 49814 470935 49816
rect 470869 49811 470935 49814
rect 469213 49738 469279 49741
rect 466912 49736 469279 49738
rect 466912 49680 469218 49736
rect 469274 49680 469279 49736
rect 466912 49678 469279 49680
rect 446213 49675 446279 49678
rect 447777 49675 447843 49678
rect 450721 49675 450787 49678
rect 454033 49675 454099 49678
rect 458265 49675 458331 49678
rect 459553 49675 459619 49678
rect 463969 49675 464035 49678
rect 469213 49675 469279 49678
rect 470593 49738 470659 49741
rect 471788 49738 471848 50048
rect 470593 49736 471848 49738
rect 470593 49680 470598 49736
rect 470654 49680 471848 49736
rect 470593 49678 471848 49680
rect 472708 49738 472768 50048
rect 474457 49738 474523 49741
rect 472708 49736 474523 49738
rect 472708 49680 474462 49736
rect 474518 49680 474523 49736
rect 472708 49678 474523 49680
rect 474640 49738 474700 50048
rect 475652 49874 475712 50048
rect 477584 49874 477644 50048
rect 479516 50010 479576 50048
rect 480253 50010 480319 50013
rect 479516 50008 480319 50010
rect 479516 49952 480258 50008
rect 480314 49952 480319 50008
rect 479516 49950 480319 49952
rect 480253 49947 480319 49950
rect 480345 49874 480411 49877
rect 475652 49814 476498 49874
rect 477584 49872 480411 49874
rect 477584 49816 480350 49872
rect 480406 49816 480411 49872
rect 477584 49814 480411 49816
rect 476297 49738 476363 49741
rect 474640 49736 476363 49738
rect 474640 49680 476302 49736
rect 476358 49680 476363 49736
rect 474640 49678 476363 49680
rect 476438 49738 476498 49814
rect 480345 49811 480411 49814
rect 477493 49738 477559 49741
rect 476438 49736 477559 49738
rect 476438 49680 477498 49736
rect 477554 49680 477559 49736
rect 476438 49678 477559 49680
rect 470593 49675 470659 49678
rect 474457 49675 474523 49678
rect 476297 49675 476363 49678
rect 477493 49675 477559 49678
rect 480253 49738 480319 49741
rect 481357 49738 481423 49741
rect 480253 49736 481423 49738
rect 480253 49680 480258 49736
rect 480314 49680 481362 49736
rect 481418 49680 481423 49736
rect 480253 49678 481423 49680
rect 481540 49738 481600 50048
rect 483105 49738 483171 49741
rect 481540 49736 483171 49738
rect 481540 49680 483110 49736
rect 483166 49680 483171 49736
rect 481540 49678 483171 49680
rect 483472 49738 483532 50048
rect 484392 49874 484452 50048
rect 484577 50010 484643 50013
rect 485404 50010 485464 50048
rect 484577 50008 485464 50010
rect 484577 49952 484582 50008
rect 484638 49952 485464 50008
rect 484577 49950 485464 49952
rect 484577 49947 484643 49950
rect 487429 49874 487495 49877
rect 484392 49872 487495 49874
rect 484392 49816 487434 49872
rect 487490 49816 487495 49872
rect 484392 49814 487495 49816
rect 487429 49811 487495 49814
rect 485773 49738 485839 49741
rect 483472 49736 485839 49738
rect 483472 49680 485778 49736
rect 485834 49680 485839 49736
rect 483472 49678 485839 49680
rect 488348 49738 488408 50048
rect 488582 49874 488642 50222
rect 489268 50116 489328 50494
rect 491293 50491 491359 50494
rect 492857 50282 492923 50285
rect 495433 50282 495499 50285
rect 490280 50280 492923 50282
rect 490280 50224 492862 50280
rect 492918 50224 492923 50280
rect 490280 50222 492923 50224
rect 490280 50116 490340 50222
rect 492857 50219 492923 50222
rect 493224 50280 495499 50282
rect 493224 50224 495438 50280
rect 495494 50224 495499 50280
rect 493224 50222 495499 50224
rect 493224 50116 493284 50222
rect 495433 50219 495499 50222
rect 496076 50116 496136 50630
rect 498285 50627 498351 50630
rect 542812 50688 545271 50690
rect 542812 50632 545210 50688
rect 545266 50632 545271 50688
rect 542812 50630 545271 50632
rect 499665 50554 499731 50557
rect 501045 50554 501111 50557
rect 507945 50554 508011 50557
rect 514845 50554 514911 50557
rect 530025 50554 530091 50557
rect 498008 50552 499731 50554
rect 498008 50496 499670 50552
rect 499726 50496 499731 50552
rect 498008 50494 499731 50496
rect 498008 50116 498068 50494
rect 499665 50491 499731 50494
rect 500358 50552 501111 50554
rect 500358 50496 501050 50552
rect 501106 50496 501111 50552
rect 500358 50494 501111 50496
rect 500358 50418 500418 50494
rect 501045 50491 501111 50494
rect 505828 50552 508011 50554
rect 505828 50496 507950 50552
rect 508006 50496 508011 50552
rect 505828 50494 508011 50496
rect 503713 50418 503779 50421
rect 499020 50358 500418 50418
rect 500952 50416 503779 50418
rect 500952 50360 503718 50416
rect 503774 50360 503779 50416
rect 500952 50358 503779 50360
rect 499020 50116 499080 50358
rect 500952 50116 501012 50358
rect 503713 50355 503779 50358
rect 505093 50282 505159 50285
rect 502884 50280 505159 50282
rect 502884 50224 505098 50280
rect 505154 50224 505159 50280
rect 502884 50222 505159 50224
rect 502884 50116 502944 50222
rect 505093 50219 505159 50222
rect 505828 50116 505888 50494
rect 507945 50491 508011 50494
rect 512636 50552 514911 50554
rect 512636 50496 514850 50552
rect 514906 50496 514911 50552
rect 512636 50494 514911 50496
rect 509509 50418 509575 50421
rect 506840 50416 509575 50418
rect 506840 50360 509514 50416
rect 509570 50360 509575 50416
rect 506840 50358 509575 50360
rect 506840 50116 506900 50358
rect 509509 50355 509575 50358
rect 512085 50282 512151 50285
rect 509692 50280 512151 50282
rect 509692 50224 512090 50280
rect 512146 50224 512151 50280
rect 509692 50222 512151 50224
rect 509692 50116 509752 50222
rect 512085 50219 512151 50222
rect 512636 50116 512696 50494
rect 514845 50491 514911 50494
rect 527264 50552 530091 50554
rect 527264 50496 530030 50552
rect 530086 50496 530091 50552
rect 527264 50494 530091 50496
rect 516133 50418 516199 50421
rect 518985 50418 519051 50421
rect 513648 50416 516199 50418
rect 513648 50360 516138 50416
rect 516194 50360 516199 50416
rect 513648 50358 516199 50360
rect 513648 50116 513708 50358
rect 516133 50355 516199 50358
rect 516500 50416 519051 50418
rect 516500 50360 518990 50416
rect 519046 50360 519051 50416
rect 516500 50358 519051 50360
rect 516500 50116 516560 50358
rect 518985 50355 519051 50358
rect 520273 50282 520339 50285
rect 523033 50282 523099 50285
rect 525885 50282 525951 50285
rect 527081 50282 527147 50285
rect 518524 50280 520339 50282
rect 518524 50224 520278 50280
rect 520334 50224 520339 50280
rect 518524 50222 520339 50224
rect 518524 50116 518584 50222
rect 520273 50219 520339 50222
rect 520456 50280 523099 50282
rect 520456 50224 523038 50280
rect 523094 50224 523099 50280
rect 520456 50222 523099 50224
rect 520456 50116 520516 50222
rect 523033 50219 523099 50222
rect 523308 50280 525951 50282
rect 523308 50224 525890 50280
rect 525946 50224 525951 50280
rect 523308 50222 525951 50224
rect 523308 50116 523368 50222
rect 525885 50219 525951 50222
rect 526118 50280 527147 50282
rect 526118 50224 527086 50280
rect 527142 50224 527147 50280
rect 526118 50222 527147 50224
rect 526118 50146 526178 50222
rect 527081 50219 527147 50222
rect 525362 50086 526178 50146
rect 527264 50116 527324 50494
rect 530025 50491 530091 50494
rect 532693 50418 532759 50421
rect 536833 50418 536899 50421
rect 531638 50416 532759 50418
rect 531638 50360 532698 50416
rect 532754 50360 532759 50416
rect 531638 50358 532759 50360
rect 531313 50282 531379 50285
rect 529196 50280 531379 50282
rect 529196 50224 531318 50280
rect 531374 50224 531379 50280
rect 529196 50222 531379 50224
rect 529196 50116 529256 50222
rect 531313 50219 531379 50222
rect 531638 50146 531698 50358
rect 532693 50355 532759 50358
rect 534582 50416 536899 50418
rect 534582 50360 536838 50416
rect 536894 50360 536899 50416
rect 534582 50358 536899 50360
rect 534165 50282 534231 50285
rect 531158 50086 531698 50146
rect 532140 50280 534231 50282
rect 532140 50224 534170 50280
rect 534226 50224 534231 50280
rect 532140 50222 534231 50224
rect 532140 50116 532200 50222
rect 534165 50219 534231 50222
rect 534582 50146 534642 50358
rect 536833 50355 536899 50358
rect 537477 50418 537543 50421
rect 539685 50418 539751 50421
rect 542353 50418 542419 50421
rect 537477 50416 539751 50418
rect 537477 50360 537482 50416
rect 537538 50360 539690 50416
rect 539746 50360 539751 50416
rect 537477 50358 539751 50360
rect 537477 50355 537543 50358
rect 539685 50355 539751 50358
rect 539868 50416 542419 50418
rect 539868 50360 542358 50416
rect 542414 50360 542419 50416
rect 539868 50358 542419 50360
rect 538305 50282 538371 50285
rect 534102 50086 534642 50146
rect 536004 50280 538371 50282
rect 536004 50224 538310 50280
rect 538366 50224 538371 50280
rect 536004 50222 538371 50224
rect 536004 50116 536064 50222
rect 538305 50219 538371 50222
rect 537477 50146 537543 50149
rect 537046 50144 537543 50146
rect 537046 50088 537482 50144
rect 537538 50088 537543 50144
rect 539868 50116 539928 50358
rect 542353 50355 542419 50358
rect 542812 50116 542872 50630
rect 545205 50627 545271 50630
rect 546769 50554 546835 50557
rect 543824 50552 546835 50554
rect 543824 50496 546774 50552
rect 546830 50496 546835 50552
rect 543824 50494 546835 50496
rect 543824 50116 543884 50494
rect 546769 50491 546835 50494
rect 549529 50418 549595 50421
rect 553485 50418 553551 50421
rect 556153 50418 556219 50421
rect 565905 50418 565971 50421
rect 570229 50418 570295 50421
rect 573081 50418 573147 50421
rect 575565 50418 575631 50421
rect 580257 50418 580323 50421
rect 546676 50416 549595 50418
rect 546676 50360 549534 50416
rect 549590 50360 549595 50416
rect 546676 50358 549595 50360
rect 546676 50116 546736 50358
rect 549529 50355 549595 50358
rect 552246 50416 553551 50418
rect 552246 50360 553490 50416
rect 553546 50360 553551 50416
rect 552246 50358 553551 50360
rect 549345 50282 549411 50285
rect 552013 50282 552079 50285
rect 547688 50280 549411 50282
rect 547688 50224 549350 50280
rect 549406 50224 549411 50280
rect 547688 50222 549411 50224
rect 547688 50116 547748 50222
rect 549345 50219 549411 50222
rect 549620 50280 552079 50282
rect 549620 50224 552018 50280
rect 552074 50224 552079 50280
rect 549620 50222 552079 50224
rect 549620 50116 549680 50222
rect 552013 50219 552079 50222
rect 552246 50146 552306 50358
rect 553485 50355 553551 50358
rect 555006 50416 556219 50418
rect 555006 50360 556158 50416
rect 556214 50360 556219 50416
rect 555006 50358 556219 50360
rect 554865 50282 554931 50285
rect 537046 50086 537543 50088
rect 551582 50086 552306 50146
rect 552564 50280 554931 50282
rect 552564 50224 554870 50280
rect 554926 50224 554931 50280
rect 552564 50222 554931 50224
rect 552564 50116 552624 50222
rect 554865 50219 554931 50222
rect 555006 50146 555066 50358
rect 556153 50355 556219 50358
rect 564758 50416 565971 50418
rect 564758 50360 565910 50416
rect 565966 50360 565971 50416
rect 564758 50358 565971 50360
rect 557533 50282 557599 50285
rect 559097 50282 559163 50285
rect 561765 50282 561831 50285
rect 564525 50282 564591 50285
rect 554526 50086 555066 50146
rect 555508 50280 557599 50282
rect 555508 50224 557538 50280
rect 557594 50224 557599 50280
rect 555508 50222 557599 50224
rect 555508 50116 555568 50222
rect 557533 50219 557599 50222
rect 558134 50280 559163 50282
rect 558134 50224 559102 50280
rect 559158 50224 559163 50280
rect 558134 50222 559163 50224
rect 557625 50146 557691 50149
rect 557470 50144 557691 50146
rect 557470 50088 557630 50144
rect 557686 50088 557691 50144
rect 557470 50086 557691 50088
rect 537477 50083 537543 50086
rect 557625 50083 557691 50086
rect 490189 49874 490255 49877
rect 488582 49872 490255 49874
rect 488582 49816 490194 49872
rect 490250 49816 490255 49872
rect 488582 49814 490255 49816
rect 490189 49811 490255 49814
rect 490005 49738 490071 49741
rect 488348 49736 490071 49738
rect 488348 49680 490010 49736
rect 490066 49680 490071 49736
rect 488348 49678 490071 49680
rect 491200 49738 491260 50048
rect 492212 49874 492272 50048
rect 494144 49874 494204 50048
rect 495156 50010 495216 50048
rect 495893 50010 495959 50013
rect 495156 50008 495959 50010
rect 495156 49952 495898 50008
rect 495954 49952 495959 50008
rect 495156 49950 495959 49952
rect 495893 49947 495959 49950
rect 496905 49874 496971 49877
rect 492212 49814 492874 49874
rect 494144 49872 496971 49874
rect 494144 49816 496910 49872
rect 496966 49816 496971 49872
rect 494144 49814 496971 49816
rect 497088 49874 497148 50048
rect 499849 49874 499915 49877
rect 497088 49872 499915 49874
rect 497088 49816 499854 49872
rect 499910 49816 499915 49872
rect 497088 49814 499915 49816
rect 492673 49738 492739 49741
rect 491200 49736 492739 49738
rect 491200 49680 492678 49736
rect 492734 49680 492739 49736
rect 491200 49678 492739 49680
rect 492814 49738 492874 49814
rect 496905 49811 496971 49814
rect 499849 49811 499915 49814
rect 494145 49738 494211 49741
rect 492814 49736 494211 49738
rect 492814 49680 494150 49736
rect 494206 49680 494211 49736
rect 492814 49678 494211 49680
rect 480253 49675 480319 49678
rect 481357 49675 481423 49678
rect 483105 49675 483171 49678
rect 485773 49675 485839 49678
rect 490005 49675 490071 49678
rect 492673 49675 492739 49678
rect 494145 49675 494211 49678
rect 495893 49738 495959 49741
rect 497089 49738 497155 49741
rect 495893 49736 497155 49738
rect 495893 49680 495898 49736
rect 495954 49680 497094 49736
rect 497150 49680 497155 49736
rect 495893 49678 497155 49680
rect 500032 49738 500092 50048
rect 501964 49874 502024 50048
rect 503896 49874 503956 50048
rect 504816 50010 504876 50048
rect 505645 50010 505711 50013
rect 504816 50008 505711 50010
rect 504816 49952 505650 50008
rect 505706 49952 505711 50008
rect 504816 49950 505711 49952
rect 505645 49947 505711 49950
rect 506565 49874 506631 49877
rect 501964 49814 502626 49874
rect 503896 49872 506631 49874
rect 503896 49816 506570 49872
rect 506626 49816 506631 49872
rect 503896 49814 506631 49816
rect 502333 49738 502399 49741
rect 500032 49736 502399 49738
rect 500032 49680 502338 49736
rect 502394 49680 502399 49736
rect 500032 49678 502399 49680
rect 502566 49738 502626 49814
rect 506565 49811 506631 49814
rect 503897 49738 503963 49741
rect 502566 49736 503963 49738
rect 502566 49680 503902 49736
rect 503958 49680 503963 49736
rect 502566 49678 503963 49680
rect 495893 49675 495959 49678
rect 497089 49675 497155 49678
rect 502333 49675 502399 49678
rect 503897 49675 503963 49678
rect 505645 49738 505711 49741
rect 506749 49738 506815 49741
rect 505645 49736 506815 49738
rect 505645 49680 505650 49736
rect 505706 49680 506754 49736
rect 506810 49680 506815 49736
rect 505645 49678 506815 49680
rect 507760 49738 507820 50048
rect 508772 49874 508832 50048
rect 510704 49874 510764 50048
rect 511716 50010 511776 50048
rect 512453 50010 512519 50013
rect 511716 50008 512519 50010
rect 511716 49952 512458 50008
rect 512514 49952 512519 50008
rect 511716 49950 512519 49952
rect 512453 49947 512519 49950
rect 513649 49874 513715 49877
rect 508772 49814 509986 49874
rect 510704 49872 513715 49874
rect 510704 49816 513654 49872
rect 513710 49816 513715 49872
rect 510704 49814 513715 49816
rect 509325 49738 509391 49741
rect 507760 49736 509391 49738
rect 507760 49680 509330 49736
rect 509386 49680 509391 49736
rect 507760 49678 509391 49680
rect 509926 49738 509986 49814
rect 513649 49811 513715 49814
rect 510705 49738 510771 49741
rect 509926 49736 510771 49738
rect 509926 49680 510710 49736
rect 510766 49680 510771 49736
rect 509926 49678 510771 49680
rect 505645 49675 505711 49678
rect 506749 49675 506815 49678
rect 509325 49675 509391 49678
rect 510705 49675 510771 49678
rect 512453 49738 512519 49741
rect 513465 49738 513531 49741
rect 512453 49736 513531 49738
rect 512453 49680 512458 49736
rect 512514 49680 513470 49736
rect 513526 49680 513531 49736
rect 512453 49678 513531 49680
rect 514568 49738 514628 50048
rect 515580 49874 515640 50048
rect 517512 50010 517572 50048
rect 517697 50010 517763 50013
rect 517512 50008 517763 50010
rect 517512 49952 517702 50008
rect 517758 49952 517763 50008
rect 517512 49950 517763 49952
rect 517697 49947 517763 49950
rect 517513 49874 517579 49877
rect 515580 49872 517579 49874
rect 515580 49816 517518 49872
rect 517574 49816 517579 49872
rect 515580 49814 517579 49816
rect 517513 49811 517579 49814
rect 516317 49738 516383 49741
rect 514568 49736 516383 49738
rect 514568 49680 516322 49736
rect 516378 49680 516383 49736
rect 514568 49678 516383 49680
rect 512453 49675 512519 49678
rect 513465 49675 513531 49678
rect 516317 49675 516383 49678
rect 519169 49738 519235 49741
rect 519444 49738 519504 50048
rect 519169 49736 519504 49738
rect 519169 49680 519174 49736
rect 519230 49680 519504 49736
rect 519169 49678 519504 49680
rect 521376 49738 521436 50048
rect 522388 49874 522448 50048
rect 524137 49874 524203 49877
rect 522388 49872 524203 49874
rect 522388 49816 524142 49872
rect 524198 49816 524203 49872
rect 522388 49814 524203 49816
rect 524137 49811 524203 49814
rect 523217 49738 523283 49741
rect 521376 49736 523283 49738
rect 521376 49680 523222 49736
rect 523278 49680 523283 49736
rect 521376 49678 523283 49680
rect 524320 49738 524380 50048
rect 526069 49738 526135 49741
rect 524320 49736 526135 49738
rect 524320 49680 526074 49736
rect 526130 49680 526135 49736
rect 524320 49678 526135 49680
rect 526252 49738 526312 50048
rect 528184 49874 528244 50048
rect 530208 49874 530268 50048
rect 532877 49874 532943 49877
rect 528184 49814 529490 49874
rect 530208 49872 532943 49874
rect 530208 49816 532882 49872
rect 532938 49816 532943 49872
rect 530208 49814 532943 49816
rect 528553 49738 528619 49741
rect 526252 49736 528619 49738
rect 526252 49680 528558 49736
rect 528614 49680 528619 49736
rect 526252 49678 528619 49680
rect 529430 49738 529490 49814
rect 532877 49811 532943 49814
rect 530209 49738 530275 49741
rect 529430 49736 530275 49738
rect 529430 49680 530214 49736
rect 530270 49680 530275 49736
rect 529430 49678 530275 49680
rect 533060 49738 533120 50048
rect 534992 49874 535052 50048
rect 537109 49874 537175 49877
rect 534992 49872 537175 49874
rect 534992 49816 537114 49872
rect 537170 49816 537175 49872
rect 534992 49814 537175 49816
rect 537109 49811 537175 49814
rect 535453 49738 535519 49741
rect 533060 49736 535519 49738
rect 533060 49680 535458 49736
rect 535514 49680 535519 49736
rect 533060 49678 535519 49680
rect 537936 49738 537996 50048
rect 538948 49874 539008 50048
rect 540697 49874 540763 49877
rect 538948 49872 540763 49874
rect 538948 49816 540702 49872
rect 540758 49816 540763 49872
rect 538948 49814 540763 49816
rect 540697 49811 540763 49814
rect 539685 49738 539751 49741
rect 537936 49736 539751 49738
rect 537936 49680 539690 49736
rect 539746 49680 539751 49736
rect 537936 49678 539751 49680
rect 540880 49738 540940 50048
rect 541892 49874 541952 50048
rect 543825 49874 543891 49877
rect 541892 49872 543891 49874
rect 541892 49816 543830 49872
rect 543886 49816 543891 49872
rect 541892 49814 543891 49816
rect 543825 49811 543891 49814
rect 542537 49738 542603 49741
rect 540880 49736 542603 49738
rect 540880 49680 542542 49736
rect 542598 49680 542603 49736
rect 540880 49678 542603 49680
rect 544744 49738 544804 50048
rect 545756 49874 545816 50048
rect 548057 49874 548123 49877
rect 545756 49872 548123 49874
rect 545756 49816 548062 49872
rect 548118 49816 548123 49872
rect 545756 49814 548123 49816
rect 548057 49811 548123 49814
rect 546585 49738 546651 49741
rect 544744 49736 546651 49738
rect 544744 49680 546590 49736
rect 546646 49680 546651 49736
rect 544744 49678 546651 49680
rect 548700 49738 548760 50048
rect 550632 49874 550692 50048
rect 553484 50010 553544 50048
rect 553484 49950 553962 50010
rect 553669 49874 553735 49877
rect 550632 49872 553735 49874
rect 550632 49816 553674 49872
rect 553730 49816 553735 49872
rect 550632 49814 553735 49816
rect 553902 49874 553962 49950
rect 556245 49874 556311 49877
rect 553902 49872 556311 49874
rect 553902 49816 556250 49872
rect 556306 49816 556311 49872
rect 553902 49814 556311 49816
rect 556428 49874 556488 50048
rect 558134 49874 558194 50222
rect 559097 50219 559163 50222
rect 559372 50280 561831 50282
rect 559372 50224 561770 50280
rect 561826 50224 561831 50280
rect 559372 50222 561831 50224
rect 559372 50116 559432 50222
rect 561765 50219 561831 50222
rect 562316 50280 564591 50282
rect 562316 50224 564530 50280
rect 564586 50224 564591 50280
rect 562316 50222 564591 50224
rect 562316 50116 562376 50222
rect 564525 50219 564591 50222
rect 564758 50146 564818 50358
rect 565905 50355 565971 50358
rect 567702 50416 570295 50418
rect 567702 50360 570234 50416
rect 570290 50360 570295 50416
rect 567702 50358 570295 50360
rect 567101 50282 567167 50285
rect 564278 50086 564818 50146
rect 565168 50280 567167 50282
rect 565168 50224 567106 50280
rect 567162 50224 567167 50280
rect 565168 50222 567167 50224
rect 565168 50116 565228 50222
rect 567101 50219 567167 50222
rect 567702 50146 567762 50358
rect 570229 50355 570295 50358
rect 571566 50416 573147 50418
rect 571566 50360 573086 50416
rect 573142 50360 573147 50416
rect 571566 50358 573147 50360
rect 571333 50282 571399 50285
rect 567222 50086 567762 50146
rect 569124 50280 571399 50282
rect 569124 50224 571338 50280
rect 571394 50224 571399 50280
rect 569124 50222 571399 50224
rect 569124 50116 569184 50222
rect 571333 50219 571399 50222
rect 571566 50146 571626 50358
rect 573081 50355 573147 50358
rect 574510 50416 575631 50418
rect 574510 50360 575570 50416
rect 575626 50360 575631 50416
rect 574510 50358 575631 50360
rect 574093 50282 574159 50285
rect 571086 50086 571626 50146
rect 572068 50280 574159 50282
rect 572068 50224 574098 50280
rect 574154 50224 574159 50280
rect 572068 50222 574159 50224
rect 572068 50116 572128 50222
rect 574093 50219 574159 50222
rect 574510 50146 574570 50358
rect 575565 50355 575631 50358
rect 577864 50416 580323 50418
rect 577864 50360 580262 50416
rect 580318 50360 580323 50416
rect 577864 50358 580323 50360
rect 576945 50282 577011 50285
rect 574030 50086 574570 50146
rect 574920 50280 577011 50282
rect 574920 50224 576950 50280
rect 577006 50224 577011 50280
rect 574920 50222 577011 50224
rect 574920 50116 574980 50222
rect 576945 50219 577011 50222
rect 577864 50116 577924 50358
rect 580257 50355 580323 50358
rect 582281 50282 582347 50285
rect 578876 50280 582347 50282
rect 578876 50224 582286 50280
rect 582342 50224 582347 50280
rect 578876 50222 582347 50224
rect 578876 50116 578936 50222
rect 582281 50219 582347 50222
rect 556428 49814 558194 49874
rect 553669 49811 553735 49814
rect 556245 49811 556311 49814
rect 550725 49738 550791 49741
rect 548700 49736 550791 49738
rect 548700 49680 550730 49736
rect 550786 49680 550791 49736
rect 548700 49678 550791 49680
rect 558360 49738 558420 50048
rect 560384 49877 560444 50048
rect 560384 49872 560451 49877
rect 560384 49816 560390 49872
rect 560446 49816 560451 49872
rect 560384 49814 560451 49816
rect 560385 49811 560451 49814
rect 560293 49738 560359 49741
rect 558360 49736 560359 49738
rect 558360 49680 560298 49736
rect 560354 49680 560359 49736
rect 558360 49678 560359 49680
rect 561304 49738 561364 50048
rect 563236 49874 563296 50048
rect 565997 49874 566063 49877
rect 563236 49872 566063 49874
rect 563236 49816 566002 49872
rect 566058 49816 566063 49872
rect 563236 49814 566063 49816
rect 565997 49811 566063 49814
rect 563237 49738 563303 49741
rect 561304 49736 563303 49738
rect 561304 49680 563242 49736
rect 563298 49680 563303 49736
rect 561304 49678 563303 49680
rect 566180 49738 566240 50048
rect 568112 49874 568172 50048
rect 570044 50010 570104 50048
rect 570044 49950 570338 50010
rect 570045 49874 570111 49877
rect 568112 49872 570111 49874
rect 568112 49816 570050 49872
rect 570106 49816 570111 49872
rect 568112 49814 570111 49816
rect 570278 49874 570338 49950
rect 572805 49874 572871 49877
rect 570278 49872 572871 49874
rect 570278 49816 572810 49872
rect 572866 49816 572871 49872
rect 570278 49814 572871 49816
rect 572988 49874 573048 50048
rect 575749 49874 575815 49877
rect 572988 49872 575815 49874
rect 572988 49816 575754 49872
rect 575810 49816 575815 49872
rect 572988 49814 575815 49816
rect 570045 49811 570111 49814
rect 572805 49811 572871 49814
rect 575749 49811 575815 49814
rect 568665 49738 568731 49741
rect 566180 49736 568731 49738
rect 566180 49680 568670 49736
rect 568726 49680 568731 49736
rect 566180 49678 568731 49680
rect 575932 49738 575992 50048
rect 578233 49738 578299 49741
rect 575932 49736 578299 49738
rect 575932 49680 578238 49736
rect 578294 49680 578299 49736
rect 575932 49678 578299 49680
rect 579612 49738 579672 50048
rect 582465 49738 582531 49741
rect 579612 49736 582531 49738
rect 579612 49680 582470 49736
rect 582526 49680 582531 49736
rect 579612 49678 582531 49680
rect 519169 49675 519235 49678
rect 523217 49675 523283 49678
rect 526069 49675 526135 49678
rect 528553 49675 528619 49678
rect 530209 49675 530275 49678
rect 535453 49675 535519 49678
rect 539685 49675 539751 49678
rect 542537 49675 542603 49678
rect 546585 49675 546651 49678
rect 550725 49675 550791 49678
rect 560293 49675 560359 49678
rect 563237 49675 563303 49678
rect 568665 49675 568731 49678
rect 578233 49675 578299 49678
rect 582465 49675 582531 49678
rect 443729 49602 443795 49605
rect 442398 49600 443795 49602
rect 442398 49544 443734 49600
rect 443790 49544 443795 49600
rect 442398 49542 443795 49544
rect 101397 49539 101463 49542
rect 130377 49539 130443 49542
rect 188337 49539 188403 49542
rect 198181 49539 198247 49542
rect 207657 49539 207723 49542
rect 217501 49539 217567 49542
rect 246849 49539 246915 49542
rect 275921 49539 275987 49542
rect 296621 49539 296687 49542
rect 314469 49539 314535 49542
rect 323945 49539 324011 49542
rect 424317 49539 424383 49542
rect 443729 49539 443795 49542
rect 583520 46188 584960 46428
rect -960 35036 480 35276
rect 583520 32996 584960 33236
rect 583520 19668 584960 19908
rect -960 11644 480 11884
rect 583520 6476 584960 6716
rect 6453 3362 6519 3365
rect 199377 3362 199443 3365
rect 6453 3360 199443 3362
rect 6453 3304 6458 3360
rect 6514 3304 199382 3360
rect 199438 3304 199443 3360
rect 6453 3302 199443 3304
rect 6453 3299 6519 3302
rect 199377 3299 199443 3302
rect 429653 3362 429719 3365
rect 537109 3362 537175 3365
rect 429653 3360 537175 3362
rect 429653 3304 429658 3360
rect 429714 3304 537114 3360
rect 537170 3304 537175 3360
rect 429653 3302 537175 3304
rect 429653 3299 429719 3302
rect 537109 3299 537175 3302
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 356614 67574 392058
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176614 67574 212058
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66954 140614 67574 176058
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 104614 67574 140058
rect 66954 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 67574 104614
rect 66954 104294 67574 104378
rect 66954 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 67574 104294
rect 66954 68614 67574 104058
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 115174 78134 150618
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 77514 79174 78134 114618
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 370894 81854 406338
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 262894 81854 298338
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 226894 81854 262338
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 118894 81854 154338
rect 81234 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 81854 118894
rect 81234 118574 81854 118658
rect 81234 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 81854 118574
rect 81234 82894 81854 118338
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 374614 85574 410058
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 266614 85574 302058
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 122614 85574 158058
rect 84954 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 85574 122614
rect 84954 122294 85574 122378
rect 84954 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 85574 122294
rect 84954 86614 85574 122058
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 552004 99854 568338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 552004 103574 572058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 552004 110414 578898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 552004 114134 582618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 552004 117854 586338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 552004 121574 554058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 552004 128414 560898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 552004 132134 564618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 552004 135854 568338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 552004 139574 572058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 552004 146414 578898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 552004 150134 582618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 552004 153854 586338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 552004 157574 554058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 552004 164414 560898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 552004 168134 564618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 552004 171854 568338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 552004 175574 572058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 552004 182414 578898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 552004 186134 582618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 552004 189854 586338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 552004 193574 554058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 552004 200414 560898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 552004 204134 564618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 552004 207854 568338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 552004 211574 572058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 552004 218414 578898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 552004 222134 582618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 552004 225854 586338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 552004 229574 554058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 552004 236414 560898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 552004 240134 564618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 552004 243854 568338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 552004 247574 572058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 552004 254414 578898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 552004 258134 582618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 552004 261854 586338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 552004 265574 554058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 552004 272414 560898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 552004 276134 564618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 552004 279854 568338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 552004 283574 572058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 552004 290414 578898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 552004 294134 582618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 552004 297854 586338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 552004 301574 554058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 552004 308414 560898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 552004 312134 564618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 552004 315854 568338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 552004 319574 572058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 552004 326414 578898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 552004 330134 582618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 552004 333854 586338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 552004 337574 554058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 552004 344414 560898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 552004 348134 564618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 552004 351854 568338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 552004 355574 572058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 552004 362414 578898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 552004 366134 582618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 552004 369854 586338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 552004 373574 554058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 552004 380414 560898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 552004 384134 564618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 552004 387854 568338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 552004 391574 572058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 552004 398414 578898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 552004 402134 582618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 552004 405854 586338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 552004 409574 554058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 552004 416414 560898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 552004 420134 564618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 552004 423854 568338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 552004 427574 572058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 552004 434414 578898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 552004 438134 582618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 552004 441854 586338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 552004 445574 554058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 552004 452414 560898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 552004 456134 564618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 552004 459854 568338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 552004 463574 572058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 552004 470414 578898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 552004 474134 582618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 552004 477854 586338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 552004 481574 554058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 552004 488414 560898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 552004 492134 564618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 552004 495854 568338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 552004 499574 572058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 552004 506414 578898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 552004 510134 582618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 552004 513854 586338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 552004 517574 554058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 552004 524414 560898
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 552004 528134 564618
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 552004 531854 568338
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 552004 535574 572058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 552004 542414 578898
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 552004 546134 582618
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 552004 549854 586338
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 552004 553574 554058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 552004 560414 560898
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 552004 564134 564618
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 552004 567854 568338
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 552004 571574 572058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 552004 578414 578898
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 552004 582134 582618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 578300 543454 578660 543486
rect 578300 543218 578362 543454
rect 578598 543218 578660 543454
rect 578300 543134 578660 543218
rect 578300 542898 578362 543134
rect 578598 542898 578660 543134
rect 578300 542866 578660 542898
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 100584 525454 100944 525486
rect 100584 525218 100646 525454
rect 100882 525218 100944 525454
rect 100584 525134 100944 525218
rect 100584 524898 100646 525134
rect 100882 524898 100944 525134
rect 100584 524866 100944 524898
rect 579020 525454 579380 525486
rect 579020 525218 579082 525454
rect 579318 525218 579380 525454
rect 579020 525134 579380 525218
rect 579020 524898 579082 525134
rect 579318 524898 579380 525134
rect 579020 524866 579380 524898
rect 101304 507454 101664 507486
rect 101304 507218 101366 507454
rect 101602 507218 101664 507454
rect 101304 507134 101664 507218
rect 101304 506898 101366 507134
rect 101602 506898 101664 507134
rect 101304 506866 101664 506898
rect 578300 507454 578660 507486
rect 578300 507218 578362 507454
rect 578598 507218 578660 507454
rect 578300 507134 578660 507218
rect 578300 506898 578362 507134
rect 578598 506898 578660 507134
rect 578300 506866 578660 506898
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 100584 489454 100944 489486
rect 100584 489218 100646 489454
rect 100882 489218 100944 489454
rect 100584 489134 100944 489218
rect 100584 488898 100646 489134
rect 100882 488898 100944 489134
rect 100584 488866 100944 488898
rect 141798 489454 142158 489486
rect 141798 489218 141860 489454
rect 142096 489218 142158 489454
rect 141798 489134 142158 489218
rect 141798 488898 141860 489134
rect 142096 488898 142158 489134
rect 141798 488866 142158 488898
rect 540286 489454 540646 489486
rect 540286 489218 540348 489454
rect 540584 489218 540646 489454
rect 540286 489134 540646 489218
rect 540286 488898 540348 489134
rect 540584 488898 540646 489134
rect 540286 488866 540646 488898
rect 579020 489454 579380 489486
rect 579020 489218 579082 489454
rect 579318 489218 579380 489454
rect 579020 489134 579380 489218
rect 579020 488898 579082 489134
rect 579318 488898 579380 489134
rect 579020 488866 579380 488898
rect 101304 471454 101664 471486
rect 101304 471218 101366 471454
rect 101602 471218 101664 471454
rect 101304 471134 101664 471218
rect 101304 470898 101366 471134
rect 101602 470898 101664 471134
rect 101304 470866 101664 470898
rect 142518 471454 142878 471486
rect 142518 471218 142580 471454
rect 142816 471218 142878 471454
rect 142518 471134 142878 471218
rect 142518 470898 142580 471134
rect 142816 470898 142878 471134
rect 142518 470866 142878 470898
rect 151290 471454 151638 471486
rect 151290 471218 151346 471454
rect 151582 471218 151638 471454
rect 151290 471134 151638 471218
rect 151290 470898 151346 471134
rect 151582 470898 151638 471134
rect 151290 470866 151638 470898
rect 244994 471454 245342 471486
rect 244994 471218 245050 471454
rect 245286 471218 245342 471454
rect 244994 471134 245342 471218
rect 244994 470898 245050 471134
rect 245286 470898 245342 471134
rect 244994 470866 245342 470898
rect 436666 471454 437014 471486
rect 436666 471218 436722 471454
rect 436958 471218 437014 471454
rect 436666 471134 437014 471218
rect 436666 470898 436722 471134
rect 436958 470898 437014 471134
rect 436666 470866 437014 470898
rect 530370 471454 530718 471486
rect 530370 471218 530426 471454
rect 530662 471218 530718 471454
rect 530370 471134 530718 471218
rect 530370 470898 530426 471134
rect 530662 470898 530718 471134
rect 530370 470866 530718 470898
rect 539566 471454 539926 471486
rect 539566 471218 539628 471454
rect 539864 471218 539926 471454
rect 539566 471134 539926 471218
rect 539566 470898 539628 471134
rect 539864 470898 539926 471134
rect 539566 470866 539926 470898
rect 578300 471454 578660 471486
rect 578300 471218 578362 471454
rect 578598 471218 578660 471454
rect 578300 471134 578660 471218
rect 578300 470898 578362 471134
rect 578598 470898 578660 471134
rect 578300 470866 578660 470898
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 421174 96134 456618
rect 100584 453454 100944 453486
rect 100584 453218 100646 453454
rect 100882 453218 100944 453454
rect 100584 453134 100944 453218
rect 100584 452898 100646 453134
rect 100882 452898 100944 453134
rect 100584 452866 100944 452898
rect 141798 453454 142158 453486
rect 141798 453218 141860 453454
rect 142096 453218 142158 453454
rect 141798 453134 142158 453218
rect 141798 452898 141860 453134
rect 142096 452898 142158 453134
rect 141798 452866 142158 452898
rect 150610 453454 150958 453486
rect 150610 453218 150666 453454
rect 150902 453218 150958 453454
rect 150610 453134 150958 453218
rect 150610 452898 150666 453134
rect 150902 452898 150958 453134
rect 150610 452866 150958 452898
rect 245674 453454 246022 453486
rect 245674 453218 245730 453454
rect 245966 453218 246022 453454
rect 245674 453134 246022 453218
rect 245674 452898 245730 453134
rect 245966 452898 246022 453134
rect 245674 452866 246022 452898
rect 435986 453454 436334 453486
rect 435986 453218 436042 453454
rect 436278 453218 436334 453454
rect 435986 453134 436334 453218
rect 435986 452898 436042 453134
rect 436278 452898 436334 453134
rect 435986 452866 436334 452898
rect 531050 453454 531398 453486
rect 531050 453218 531106 453454
rect 531342 453218 531398 453454
rect 531050 453134 531398 453218
rect 531050 452898 531106 453134
rect 531342 452898 531398 453134
rect 531050 452866 531398 452898
rect 540286 453454 540646 453486
rect 540286 453218 540348 453454
rect 540584 453218 540646 453454
rect 540286 453134 540646 453218
rect 540286 452898 540348 453134
rect 540584 452898 540646 453134
rect 540286 452866 540646 452898
rect 579020 453454 579380 453486
rect 579020 453218 579082 453454
rect 579318 453218 579380 453454
rect 579020 453134 579380 453218
rect 579020 452898 579082 453134
rect 579318 452898 579380 453134
rect 579020 452866 579380 452898
rect 101304 435454 101664 435486
rect 101304 435218 101366 435454
rect 101602 435218 101664 435454
rect 101304 435134 101664 435218
rect 101304 434898 101366 435134
rect 101602 434898 101664 435134
rect 101304 434866 101664 434898
rect 142518 435454 142878 435486
rect 142518 435218 142580 435454
rect 142816 435218 142878 435454
rect 142518 435134 142878 435218
rect 142518 434898 142580 435134
rect 142816 434898 142878 435134
rect 142518 434866 142878 434898
rect 151290 435454 151638 435486
rect 151290 435218 151346 435454
rect 151582 435218 151638 435454
rect 151290 435134 151638 435218
rect 151290 434898 151346 435134
rect 151582 434898 151638 435134
rect 151290 434866 151638 434898
rect 244994 435454 245342 435486
rect 244994 435218 245050 435454
rect 245286 435218 245342 435454
rect 244994 435134 245342 435218
rect 244994 434898 245050 435134
rect 245286 434898 245342 435134
rect 244994 434866 245342 434898
rect 436666 435454 437014 435486
rect 436666 435218 436722 435454
rect 436958 435218 437014 435454
rect 436666 435134 437014 435218
rect 436666 434898 436722 435134
rect 436958 434898 437014 435134
rect 436666 434866 437014 434898
rect 530370 435454 530718 435486
rect 530370 435218 530426 435454
rect 530662 435218 530718 435454
rect 530370 435134 530718 435218
rect 530370 434898 530426 435134
rect 530662 434898 530718 435134
rect 530370 434866 530718 434898
rect 539566 435454 539926 435486
rect 539566 435218 539628 435454
rect 539864 435218 539926 435454
rect 539566 435134 539926 435218
rect 539566 434898 539628 435134
rect 539864 434898 539926 435134
rect 539566 434866 539926 434898
rect 578300 435454 578660 435486
rect 578300 435218 578362 435454
rect 578598 435218 578660 435454
rect 578300 435134 578660 435218
rect 578300 434898 578362 435134
rect 578598 434898 578660 435134
rect 578300 434866 578660 434898
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 385174 96134 420618
rect 100584 417454 100944 417486
rect 100584 417218 100646 417454
rect 100882 417218 100944 417454
rect 100584 417134 100944 417218
rect 100584 416898 100646 417134
rect 100882 416898 100944 417134
rect 100584 416866 100944 416898
rect 141798 417454 142158 417486
rect 141798 417218 141860 417454
rect 142096 417218 142158 417454
rect 141798 417134 142158 417218
rect 141798 416898 141860 417134
rect 142096 416898 142158 417134
rect 141798 416866 142158 416898
rect 150610 417454 150958 417486
rect 150610 417218 150666 417454
rect 150902 417218 150958 417454
rect 150610 417134 150958 417218
rect 150610 416898 150666 417134
rect 150902 416898 150958 417134
rect 150610 416866 150958 416898
rect 245674 417454 246022 417486
rect 245674 417218 245730 417454
rect 245966 417218 246022 417454
rect 245674 417134 246022 417218
rect 245674 416898 245730 417134
rect 245966 416898 246022 417134
rect 245674 416866 246022 416898
rect 435986 417454 436334 417486
rect 435986 417218 436042 417454
rect 436278 417218 436334 417454
rect 435986 417134 436334 417218
rect 435986 416898 436042 417134
rect 436278 416898 436334 417134
rect 435986 416866 436334 416898
rect 531050 417454 531398 417486
rect 531050 417218 531106 417454
rect 531342 417218 531398 417454
rect 531050 417134 531398 417218
rect 531050 416898 531106 417134
rect 531342 416898 531398 417134
rect 531050 416866 531398 416898
rect 540286 417454 540646 417486
rect 540286 417218 540348 417454
rect 540584 417218 540646 417454
rect 540286 417134 540646 417218
rect 540286 416898 540348 417134
rect 540584 416898 540646 417134
rect 540286 416866 540646 416898
rect 579020 417454 579380 417486
rect 579020 417218 579082 417454
rect 579318 417218 579380 417454
rect 579020 417134 579380 417218
rect 579020 416898 579082 417134
rect 579318 416898 579380 417134
rect 579020 416866 579380 416898
rect 101304 399454 101664 399486
rect 101304 399218 101366 399454
rect 101602 399218 101664 399454
rect 101304 399134 101664 399218
rect 101304 398898 101366 399134
rect 101602 398898 101664 399134
rect 101304 398866 101664 398898
rect 142518 399454 142878 399486
rect 142518 399218 142580 399454
rect 142816 399218 142878 399454
rect 142518 399134 142878 399218
rect 142518 398898 142580 399134
rect 142816 398898 142878 399134
rect 142518 398866 142878 398898
rect 539566 399454 539926 399486
rect 539566 399218 539628 399454
rect 539864 399218 539926 399454
rect 539566 399134 539926 399218
rect 539566 398898 539628 399134
rect 539864 398898 539926 399134
rect 539566 398866 539926 398898
rect 578300 399454 578660 399486
rect 578300 399218 578362 399454
rect 578598 399218 578660 399454
rect 578300 399134 578660 399218
rect 578300 398898 578362 399134
rect 578598 398898 578660 399134
rect 578300 398866 578660 398898
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 100584 381454 100944 381486
rect 100584 381218 100646 381454
rect 100882 381218 100944 381454
rect 100584 381134 100944 381218
rect 100584 380898 100646 381134
rect 100882 380898 100944 381134
rect 100584 380866 100944 380898
rect 141798 381454 142158 381486
rect 141798 381218 141860 381454
rect 142096 381218 142158 381454
rect 141798 381134 142158 381218
rect 141798 380898 141860 381134
rect 142096 380898 142158 381134
rect 141798 380866 142158 380898
rect 150610 381454 150958 381486
rect 150610 381218 150666 381454
rect 150902 381218 150958 381454
rect 150610 381134 150958 381218
rect 150610 380898 150666 381134
rect 150902 380898 150958 381134
rect 150610 380866 150958 380898
rect 245674 381454 246022 381486
rect 245674 381218 245730 381454
rect 245966 381218 246022 381454
rect 245674 381134 246022 381218
rect 245674 380898 245730 381134
rect 245966 380898 246022 381134
rect 245674 380866 246022 380898
rect 435986 381454 436334 381486
rect 435986 381218 436042 381454
rect 436278 381218 436334 381454
rect 435986 381134 436334 381218
rect 435986 380898 436042 381134
rect 436278 380898 436334 381134
rect 435986 380866 436334 380898
rect 531050 381454 531398 381486
rect 531050 381218 531106 381454
rect 531342 381218 531398 381454
rect 531050 381134 531398 381218
rect 531050 380898 531106 381134
rect 531342 380898 531398 381134
rect 531050 380866 531398 380898
rect 540286 381454 540646 381486
rect 540286 381218 540348 381454
rect 540584 381218 540646 381454
rect 540286 381134 540646 381218
rect 540286 380898 540348 381134
rect 540584 380898 540646 381134
rect 540286 380866 540646 380898
rect 579020 381454 579380 381486
rect 579020 381218 579082 381454
rect 579318 381218 579380 381454
rect 579020 381134 579380 381218
rect 579020 380898 579082 381134
rect 579318 380898 579380 381134
rect 579020 380866 579380 380898
rect 101304 363454 101664 363486
rect 101304 363218 101366 363454
rect 101602 363218 101664 363454
rect 101304 363134 101664 363218
rect 101304 362898 101366 363134
rect 101602 362898 101664 363134
rect 101304 362866 101664 362898
rect 142518 363454 142878 363486
rect 142518 363218 142580 363454
rect 142816 363218 142878 363454
rect 142518 363134 142878 363218
rect 142518 362898 142580 363134
rect 142816 362898 142878 363134
rect 142518 362866 142878 362898
rect 151290 363454 151638 363486
rect 151290 363218 151346 363454
rect 151582 363218 151638 363454
rect 151290 363134 151638 363218
rect 151290 362898 151346 363134
rect 151582 362898 151638 363134
rect 151290 362866 151638 362898
rect 244994 363454 245342 363486
rect 244994 363218 245050 363454
rect 245286 363218 245342 363454
rect 244994 363134 245342 363218
rect 244994 362898 245050 363134
rect 245286 362898 245342 363134
rect 244994 362866 245342 362898
rect 436666 363454 437014 363486
rect 436666 363218 436722 363454
rect 436958 363218 437014 363454
rect 436666 363134 437014 363218
rect 436666 362898 436722 363134
rect 436958 362898 437014 363134
rect 436666 362866 437014 362898
rect 530370 363454 530718 363486
rect 530370 363218 530426 363454
rect 530662 363218 530718 363454
rect 530370 363134 530718 363218
rect 530370 362898 530426 363134
rect 530662 362898 530718 363134
rect 530370 362866 530718 362898
rect 539566 363454 539926 363486
rect 539566 363218 539628 363454
rect 539864 363218 539926 363454
rect 539566 363134 539926 363218
rect 539566 362898 539628 363134
rect 539864 362898 539926 363134
rect 539566 362866 539926 362898
rect 578300 363454 578660 363486
rect 578300 363218 578362 363454
rect 578598 363218 578660 363454
rect 578300 363134 578660 363218
rect 578300 362898 578362 363134
rect 578598 362898 578660 363134
rect 578300 362866 578660 362898
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95514 313174 96134 348618
rect 100584 345454 100944 345486
rect 100584 345218 100646 345454
rect 100882 345218 100944 345454
rect 100584 345134 100944 345218
rect 100584 344898 100646 345134
rect 100882 344898 100944 345134
rect 100584 344866 100944 344898
rect 141798 345454 142158 345486
rect 141798 345218 141860 345454
rect 142096 345218 142158 345454
rect 141798 345134 142158 345218
rect 141798 344898 141860 345134
rect 142096 344898 142158 345134
rect 141798 344866 142158 344898
rect 150610 345454 150958 345486
rect 150610 345218 150666 345454
rect 150902 345218 150958 345454
rect 150610 345134 150958 345218
rect 150610 344898 150666 345134
rect 150902 344898 150958 345134
rect 150610 344866 150958 344898
rect 245674 345454 246022 345486
rect 245674 345218 245730 345454
rect 245966 345218 246022 345454
rect 245674 345134 246022 345218
rect 245674 344898 245730 345134
rect 245966 344898 246022 345134
rect 245674 344866 246022 344898
rect 435986 345454 436334 345486
rect 435986 345218 436042 345454
rect 436278 345218 436334 345454
rect 435986 345134 436334 345218
rect 435986 344898 436042 345134
rect 436278 344898 436334 345134
rect 435986 344866 436334 344898
rect 531050 345454 531398 345486
rect 531050 345218 531106 345454
rect 531342 345218 531398 345454
rect 531050 345134 531398 345218
rect 531050 344898 531106 345134
rect 531342 344898 531398 345134
rect 531050 344866 531398 344898
rect 540286 345454 540646 345486
rect 540286 345218 540348 345454
rect 540584 345218 540646 345454
rect 540286 345134 540646 345218
rect 540286 344898 540348 345134
rect 540584 344898 540646 345134
rect 540286 344866 540646 344898
rect 579020 345454 579380 345486
rect 579020 345218 579082 345454
rect 579318 345218 579380 345454
rect 579020 345134 579380 345218
rect 579020 344898 579082 345134
rect 579318 344898 579380 345134
rect 579020 344866 579380 344898
rect 101304 327454 101664 327486
rect 101304 327218 101366 327454
rect 101602 327218 101664 327454
rect 101304 327134 101664 327218
rect 101304 326898 101366 327134
rect 101602 326898 101664 327134
rect 101304 326866 101664 326898
rect 142518 327454 142878 327486
rect 142518 327218 142580 327454
rect 142816 327218 142878 327454
rect 142518 327134 142878 327218
rect 142518 326898 142580 327134
rect 142816 326898 142878 327134
rect 142518 326866 142878 326898
rect 151290 327454 151638 327486
rect 151290 327218 151346 327454
rect 151582 327218 151638 327454
rect 151290 327134 151638 327218
rect 151290 326898 151346 327134
rect 151582 326898 151638 327134
rect 151290 326866 151638 326898
rect 244994 327454 245342 327486
rect 244994 327218 245050 327454
rect 245286 327218 245342 327454
rect 244994 327134 245342 327218
rect 244994 326898 245050 327134
rect 245286 326898 245342 327134
rect 244994 326866 245342 326898
rect 436666 327454 437014 327486
rect 436666 327218 436722 327454
rect 436958 327218 437014 327454
rect 436666 327134 437014 327218
rect 436666 326898 436722 327134
rect 436958 326898 437014 327134
rect 436666 326866 437014 326898
rect 530370 327454 530718 327486
rect 530370 327218 530426 327454
rect 530662 327218 530718 327454
rect 530370 327134 530718 327218
rect 530370 326898 530426 327134
rect 530662 326898 530718 327134
rect 530370 326866 530718 326898
rect 539566 327454 539926 327486
rect 539566 327218 539628 327454
rect 539864 327218 539926 327454
rect 539566 327134 539926 327218
rect 539566 326898 539628 327134
rect 539864 326898 539926 327134
rect 539566 326866 539926 326898
rect 578300 327454 578660 327486
rect 578300 327218 578362 327454
rect 578598 327218 578660 327454
rect 578300 327134 578660 327218
rect 578300 326898 578362 327134
rect 578598 326898 578660 327134
rect 578300 326866 578660 326898
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 277174 96134 312618
rect 100584 309454 100944 309486
rect 100584 309218 100646 309454
rect 100882 309218 100944 309454
rect 100584 309134 100944 309218
rect 100584 308898 100646 309134
rect 100882 308898 100944 309134
rect 100584 308866 100944 308898
rect 141798 309454 142158 309486
rect 141798 309218 141860 309454
rect 142096 309218 142158 309454
rect 141798 309134 142158 309218
rect 141798 308898 141860 309134
rect 142096 308898 142158 309134
rect 141798 308866 142158 308898
rect 540286 309454 540646 309486
rect 540286 309218 540348 309454
rect 540584 309218 540646 309454
rect 540286 309134 540646 309218
rect 540286 308898 540348 309134
rect 540584 308898 540646 309134
rect 540286 308866 540646 308898
rect 579020 309454 579380 309486
rect 579020 309218 579082 309454
rect 579318 309218 579380 309454
rect 579020 309134 579380 309218
rect 579020 308898 579082 309134
rect 579318 308898 579380 309134
rect 579020 308866 579380 308898
rect 101304 291454 101664 291486
rect 101304 291218 101366 291454
rect 101602 291218 101664 291454
rect 101304 291134 101664 291218
rect 101304 290898 101366 291134
rect 101602 290898 101664 291134
rect 101304 290866 101664 290898
rect 142518 291454 142878 291486
rect 142518 291218 142580 291454
rect 142816 291218 142878 291454
rect 142518 291134 142878 291218
rect 142518 290898 142580 291134
rect 142816 290898 142878 291134
rect 142518 290866 142878 290898
rect 151290 291454 151638 291486
rect 151290 291218 151346 291454
rect 151582 291218 151638 291454
rect 151290 291134 151638 291218
rect 151290 290898 151346 291134
rect 151582 290898 151638 291134
rect 151290 290866 151638 290898
rect 244994 291454 245342 291486
rect 244994 291218 245050 291454
rect 245286 291218 245342 291454
rect 244994 291134 245342 291218
rect 244994 290898 245050 291134
rect 245286 290898 245342 291134
rect 244994 290866 245342 290898
rect 436666 291454 437014 291486
rect 436666 291218 436722 291454
rect 436958 291218 437014 291454
rect 436666 291134 437014 291218
rect 436666 290898 436722 291134
rect 436958 290898 437014 291134
rect 436666 290866 437014 290898
rect 530370 291454 530718 291486
rect 530370 291218 530426 291454
rect 530662 291218 530718 291454
rect 530370 291134 530718 291218
rect 530370 290898 530426 291134
rect 530662 290898 530718 291134
rect 530370 290866 530718 290898
rect 539566 291454 539926 291486
rect 539566 291218 539628 291454
rect 539864 291218 539926 291454
rect 539566 291134 539926 291218
rect 539566 290898 539628 291134
rect 539864 290898 539926 291134
rect 539566 290866 539926 290898
rect 578300 291454 578660 291486
rect 578300 291218 578362 291454
rect 578598 291218 578660 291454
rect 578300 291134 578660 291218
rect 578300 290898 578362 291134
rect 578598 290898 578660 291134
rect 578300 290866 578660 290898
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 95514 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 96134 277174
rect 95514 276854 96134 276938
rect 95514 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 96134 276854
rect 95514 241174 96134 276618
rect 100584 273454 100944 273486
rect 100584 273218 100646 273454
rect 100882 273218 100944 273454
rect 100584 273134 100944 273218
rect 100584 272898 100646 273134
rect 100882 272898 100944 273134
rect 100584 272866 100944 272898
rect 141798 273454 142158 273486
rect 141798 273218 141860 273454
rect 142096 273218 142158 273454
rect 141798 273134 142158 273218
rect 141798 272898 141860 273134
rect 142096 272898 142158 273134
rect 141798 272866 142158 272898
rect 150610 273454 150958 273486
rect 150610 273218 150666 273454
rect 150902 273218 150958 273454
rect 150610 273134 150958 273218
rect 150610 272898 150666 273134
rect 150902 272898 150958 273134
rect 150610 272866 150958 272898
rect 245674 273454 246022 273486
rect 245674 273218 245730 273454
rect 245966 273218 246022 273454
rect 245674 273134 246022 273218
rect 245674 272898 245730 273134
rect 245966 272898 246022 273134
rect 245674 272866 246022 272898
rect 435986 273454 436334 273486
rect 435986 273218 436042 273454
rect 436278 273218 436334 273454
rect 435986 273134 436334 273218
rect 435986 272898 436042 273134
rect 436278 272898 436334 273134
rect 435986 272866 436334 272898
rect 531050 273454 531398 273486
rect 531050 273218 531106 273454
rect 531342 273218 531398 273454
rect 531050 273134 531398 273218
rect 531050 272898 531106 273134
rect 531342 272898 531398 273134
rect 531050 272866 531398 272898
rect 540286 273454 540646 273486
rect 540286 273218 540348 273454
rect 540584 273218 540646 273454
rect 540286 273134 540646 273218
rect 540286 272898 540348 273134
rect 540584 272898 540646 273134
rect 540286 272866 540646 272898
rect 579020 273454 579380 273486
rect 579020 273218 579082 273454
rect 579318 273218 579380 273454
rect 579020 273134 579380 273218
rect 579020 272898 579082 273134
rect 579318 272898 579380 273134
rect 579020 272866 579380 272898
rect 101304 255454 101664 255486
rect 101304 255218 101366 255454
rect 101602 255218 101664 255454
rect 101304 255134 101664 255218
rect 101304 254898 101366 255134
rect 101602 254898 101664 255134
rect 101304 254866 101664 254898
rect 142518 255454 142878 255486
rect 142518 255218 142580 255454
rect 142816 255218 142878 255454
rect 142518 255134 142878 255218
rect 142518 254898 142580 255134
rect 142816 254898 142878 255134
rect 142518 254866 142878 254898
rect 151290 255454 151638 255486
rect 151290 255218 151346 255454
rect 151582 255218 151638 255454
rect 151290 255134 151638 255218
rect 151290 254898 151346 255134
rect 151582 254898 151638 255134
rect 151290 254866 151638 254898
rect 244994 255454 245342 255486
rect 244994 255218 245050 255454
rect 245286 255218 245342 255454
rect 244994 255134 245342 255218
rect 244994 254898 245050 255134
rect 245286 254898 245342 255134
rect 244994 254866 245342 254898
rect 436666 255454 437014 255486
rect 436666 255218 436722 255454
rect 436958 255218 437014 255454
rect 436666 255134 437014 255218
rect 436666 254898 436722 255134
rect 436958 254898 437014 255134
rect 436666 254866 437014 254898
rect 530370 255454 530718 255486
rect 530370 255218 530426 255454
rect 530662 255218 530718 255454
rect 530370 255134 530718 255218
rect 530370 254898 530426 255134
rect 530662 254898 530718 255134
rect 530370 254866 530718 254898
rect 539566 255454 539926 255486
rect 539566 255218 539628 255454
rect 539864 255218 539926 255454
rect 539566 255134 539926 255218
rect 539566 254898 539628 255134
rect 539864 254898 539926 255134
rect 539566 254866 539926 254898
rect 578300 255454 578660 255486
rect 578300 255218 578362 255454
rect 578598 255218 578660 255454
rect 578300 255134 578660 255218
rect 578300 254898 578362 255134
rect 578598 254898 578660 255134
rect 578300 254866 578660 254898
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 95514 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 96134 241174
rect 95514 240854 96134 240938
rect 95514 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 96134 240854
rect 95514 205174 96134 240618
rect 100584 237454 100944 237486
rect 100584 237218 100646 237454
rect 100882 237218 100944 237454
rect 100584 237134 100944 237218
rect 100584 236898 100646 237134
rect 100882 236898 100944 237134
rect 100584 236866 100944 236898
rect 141798 237454 142158 237486
rect 141798 237218 141860 237454
rect 142096 237218 142158 237454
rect 141798 237134 142158 237218
rect 141798 236898 141860 237134
rect 142096 236898 142158 237134
rect 141798 236866 142158 236898
rect 150610 237454 150958 237486
rect 150610 237218 150666 237454
rect 150902 237218 150958 237454
rect 150610 237134 150958 237218
rect 150610 236898 150666 237134
rect 150902 236898 150958 237134
rect 150610 236866 150958 236898
rect 245674 237454 246022 237486
rect 245674 237218 245730 237454
rect 245966 237218 246022 237454
rect 245674 237134 246022 237218
rect 245674 236898 245730 237134
rect 245966 236898 246022 237134
rect 245674 236866 246022 236898
rect 435986 237454 436334 237486
rect 435986 237218 436042 237454
rect 436278 237218 436334 237454
rect 435986 237134 436334 237218
rect 435986 236898 436042 237134
rect 436278 236898 436334 237134
rect 435986 236866 436334 236898
rect 531050 237454 531398 237486
rect 531050 237218 531106 237454
rect 531342 237218 531398 237454
rect 531050 237134 531398 237218
rect 531050 236898 531106 237134
rect 531342 236898 531398 237134
rect 531050 236866 531398 236898
rect 540286 237454 540646 237486
rect 540286 237218 540348 237454
rect 540584 237218 540646 237454
rect 540286 237134 540646 237218
rect 540286 236898 540348 237134
rect 540584 236898 540646 237134
rect 540286 236866 540646 236898
rect 579020 237454 579380 237486
rect 579020 237218 579082 237454
rect 579318 237218 579380 237454
rect 579020 237134 579380 237218
rect 579020 236898 579082 237134
rect 579318 236898 579380 237134
rect 579020 236866 579380 236898
rect 101304 219454 101664 219486
rect 101304 219218 101366 219454
rect 101602 219218 101664 219454
rect 101304 219134 101664 219218
rect 101304 218898 101366 219134
rect 101602 218898 101664 219134
rect 101304 218866 101664 218898
rect 142518 219454 142878 219486
rect 142518 219218 142580 219454
rect 142816 219218 142878 219454
rect 142518 219134 142878 219218
rect 142518 218898 142580 219134
rect 142816 218898 142878 219134
rect 142518 218866 142878 218898
rect 436666 219454 437014 219486
rect 436666 219218 436722 219454
rect 436958 219218 437014 219454
rect 436666 219134 437014 219218
rect 436666 218898 436722 219134
rect 436958 218898 437014 219134
rect 436666 218866 437014 218898
rect 530370 219454 530718 219486
rect 530370 219218 530426 219454
rect 530662 219218 530718 219454
rect 530370 219134 530718 219218
rect 530370 218898 530426 219134
rect 530662 218898 530718 219134
rect 530370 218866 530718 218898
rect 539566 219454 539926 219486
rect 539566 219218 539628 219454
rect 539864 219218 539926 219454
rect 539566 219134 539926 219218
rect 539566 218898 539628 219134
rect 539864 218898 539926 219134
rect 539566 218866 539926 218898
rect 578300 219454 578660 219486
rect 578300 219218 578362 219454
rect 578598 219218 578660 219454
rect 578300 219134 578660 219218
rect 578300 218898 578362 219134
rect 578598 218898 578660 219134
rect 578300 218866 578660 218898
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 169174 96134 204618
rect 100584 201454 100944 201486
rect 100584 201218 100646 201454
rect 100882 201218 100944 201454
rect 100584 201134 100944 201218
rect 100584 200898 100646 201134
rect 100882 200898 100944 201134
rect 100584 200866 100944 200898
rect 141798 201454 142158 201486
rect 141798 201218 141860 201454
rect 142096 201218 142158 201454
rect 141798 201134 142158 201218
rect 141798 200898 141860 201134
rect 142096 200898 142158 201134
rect 141798 200866 142158 200898
rect 150610 201454 150958 201486
rect 150610 201218 150666 201454
rect 150902 201218 150958 201454
rect 150610 201134 150958 201218
rect 150610 200898 150666 201134
rect 150902 200898 150958 201134
rect 150610 200866 150958 200898
rect 245674 201454 246022 201486
rect 245674 201218 245730 201454
rect 245966 201218 246022 201454
rect 245674 201134 246022 201218
rect 245674 200898 245730 201134
rect 245966 200898 246022 201134
rect 245674 200866 246022 200898
rect 435986 201454 436334 201486
rect 435986 201218 436042 201454
rect 436278 201218 436334 201454
rect 435986 201134 436334 201218
rect 435986 200898 436042 201134
rect 436278 200898 436334 201134
rect 435986 200866 436334 200898
rect 531050 201454 531398 201486
rect 531050 201218 531106 201454
rect 531342 201218 531398 201454
rect 531050 201134 531398 201218
rect 531050 200898 531106 201134
rect 531342 200898 531398 201134
rect 531050 200866 531398 200898
rect 540286 201454 540646 201486
rect 540286 201218 540348 201454
rect 540584 201218 540646 201454
rect 540286 201134 540646 201218
rect 540286 200898 540348 201134
rect 540584 200898 540646 201134
rect 540286 200866 540646 200898
rect 579020 201454 579380 201486
rect 579020 201218 579082 201454
rect 579318 201218 579380 201454
rect 579020 201134 579380 201218
rect 579020 200898 579082 201134
rect 579318 200898 579380 201134
rect 579020 200866 579380 200898
rect 101304 183454 101664 183486
rect 101304 183218 101366 183454
rect 101602 183218 101664 183454
rect 101304 183134 101664 183218
rect 101304 182898 101366 183134
rect 101602 182898 101664 183134
rect 101304 182866 101664 182898
rect 142518 183454 142878 183486
rect 142518 183218 142580 183454
rect 142816 183218 142878 183454
rect 142518 183134 142878 183218
rect 142518 182898 142580 183134
rect 142816 182898 142878 183134
rect 142518 182866 142878 182898
rect 151290 183454 151638 183486
rect 151290 183218 151346 183454
rect 151582 183218 151638 183454
rect 151290 183134 151638 183218
rect 151290 182898 151346 183134
rect 151582 182898 151638 183134
rect 151290 182866 151638 182898
rect 244994 183454 245342 183486
rect 244994 183218 245050 183454
rect 245286 183218 245342 183454
rect 244994 183134 245342 183218
rect 244994 182898 245050 183134
rect 245286 182898 245342 183134
rect 244994 182866 245342 182898
rect 436666 183454 437014 183486
rect 436666 183218 436722 183454
rect 436958 183218 437014 183454
rect 436666 183134 437014 183218
rect 436666 182898 436722 183134
rect 436958 182898 437014 183134
rect 436666 182866 437014 182898
rect 530370 183454 530718 183486
rect 530370 183218 530426 183454
rect 530662 183218 530718 183454
rect 530370 183134 530718 183218
rect 530370 182898 530426 183134
rect 530662 182898 530718 183134
rect 530370 182866 530718 182898
rect 539566 183454 539926 183486
rect 539566 183218 539628 183454
rect 539864 183218 539926 183454
rect 539566 183134 539926 183218
rect 539566 182898 539628 183134
rect 539864 182898 539926 183134
rect 539566 182866 539926 182898
rect 578300 183454 578660 183486
rect 578300 183218 578362 183454
rect 578598 183218 578660 183454
rect 578300 183134 578660 183218
rect 578300 182898 578362 183134
rect 578598 182898 578660 183134
rect 578300 182866 578660 182898
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 95514 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 96134 169174
rect 95514 168854 96134 168938
rect 95514 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 96134 168854
rect 95514 133174 96134 168618
rect 100584 165454 100944 165486
rect 100584 165218 100646 165454
rect 100882 165218 100944 165454
rect 100584 165134 100944 165218
rect 100584 164898 100646 165134
rect 100882 164898 100944 165134
rect 100584 164866 100944 164898
rect 141798 165454 142158 165486
rect 141798 165218 141860 165454
rect 142096 165218 142158 165454
rect 141798 165134 142158 165218
rect 141798 164898 141860 165134
rect 142096 164898 142158 165134
rect 141798 164866 142158 164898
rect 150610 165454 150958 165486
rect 150610 165218 150666 165454
rect 150902 165218 150958 165454
rect 150610 165134 150958 165218
rect 150610 164898 150666 165134
rect 150902 164898 150958 165134
rect 150610 164866 150958 164898
rect 245674 165454 246022 165486
rect 245674 165218 245730 165454
rect 245966 165218 246022 165454
rect 245674 165134 246022 165218
rect 245674 164898 245730 165134
rect 245966 164898 246022 165134
rect 245674 164866 246022 164898
rect 435986 165454 436334 165486
rect 435986 165218 436042 165454
rect 436278 165218 436334 165454
rect 435986 165134 436334 165218
rect 435986 164898 436042 165134
rect 436278 164898 436334 165134
rect 435986 164866 436334 164898
rect 531050 165454 531398 165486
rect 531050 165218 531106 165454
rect 531342 165218 531398 165454
rect 531050 165134 531398 165218
rect 531050 164898 531106 165134
rect 531342 164898 531398 165134
rect 531050 164866 531398 164898
rect 540286 165454 540646 165486
rect 540286 165218 540348 165454
rect 540584 165218 540646 165454
rect 540286 165134 540646 165218
rect 540286 164898 540348 165134
rect 540584 164898 540646 165134
rect 540286 164866 540646 164898
rect 579020 165454 579380 165486
rect 579020 165218 579082 165454
rect 579318 165218 579380 165454
rect 579020 165134 579380 165218
rect 579020 164898 579082 165134
rect 579318 164898 579380 165134
rect 579020 164866 579380 164898
rect 101304 147454 101664 147486
rect 101304 147218 101366 147454
rect 101602 147218 101664 147454
rect 101304 147134 101664 147218
rect 101304 146898 101366 147134
rect 101602 146898 101664 147134
rect 101304 146866 101664 146898
rect 142518 147454 142878 147486
rect 142518 147218 142580 147454
rect 142816 147218 142878 147454
rect 142518 147134 142878 147218
rect 142518 146898 142580 147134
rect 142816 146898 142878 147134
rect 142518 146866 142878 146898
rect 151290 147454 151638 147486
rect 151290 147218 151346 147454
rect 151582 147218 151638 147454
rect 151290 147134 151638 147218
rect 151290 146898 151346 147134
rect 151582 146898 151638 147134
rect 151290 146866 151638 146898
rect 244994 147454 245342 147486
rect 244994 147218 245050 147454
rect 245286 147218 245342 147454
rect 244994 147134 245342 147218
rect 244994 146898 245050 147134
rect 245286 146898 245342 147134
rect 244994 146866 245342 146898
rect 436666 147454 437014 147486
rect 436666 147218 436722 147454
rect 436958 147218 437014 147454
rect 436666 147134 437014 147218
rect 436666 146898 436722 147134
rect 436958 146898 437014 147134
rect 436666 146866 437014 146898
rect 530370 147454 530718 147486
rect 530370 147218 530426 147454
rect 530662 147218 530718 147454
rect 530370 147134 530718 147218
rect 530370 146898 530426 147134
rect 530662 146898 530718 147134
rect 530370 146866 530718 146898
rect 539566 147454 539926 147486
rect 539566 147218 539628 147454
rect 539864 147218 539926 147454
rect 539566 147134 539926 147218
rect 539566 146898 539628 147134
rect 539864 146898 539926 147134
rect 539566 146866 539926 146898
rect 578300 147454 578660 147486
rect 578300 147218 578362 147454
rect 578598 147218 578660 147454
rect 578300 147134 578660 147218
rect 578300 146898 578362 147134
rect 578598 146898 578660 147134
rect 578300 146866 578660 146898
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 95514 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 96134 133174
rect 95514 132854 96134 132938
rect 95514 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 96134 132854
rect 95514 97174 96134 132618
rect 100584 129454 100944 129486
rect 100584 129218 100646 129454
rect 100882 129218 100944 129454
rect 100584 129134 100944 129218
rect 100584 128898 100646 129134
rect 100882 128898 100944 129134
rect 100584 128866 100944 128898
rect 141798 129454 142158 129486
rect 141798 129218 141860 129454
rect 142096 129218 142158 129454
rect 141798 129134 142158 129218
rect 141798 128898 141860 129134
rect 142096 128898 142158 129134
rect 141798 128866 142158 128898
rect 150610 129454 150958 129486
rect 150610 129218 150666 129454
rect 150902 129218 150958 129454
rect 150610 129134 150958 129218
rect 150610 128898 150666 129134
rect 150902 128898 150958 129134
rect 150610 128866 150958 128898
rect 245674 129454 246022 129486
rect 245674 129218 245730 129454
rect 245966 129218 246022 129454
rect 245674 129134 246022 129218
rect 245674 128898 245730 129134
rect 245966 128898 246022 129134
rect 245674 128866 246022 128898
rect 435986 129454 436334 129486
rect 435986 129218 436042 129454
rect 436278 129218 436334 129454
rect 435986 129134 436334 129218
rect 435986 128898 436042 129134
rect 436278 128898 436334 129134
rect 435986 128866 436334 128898
rect 531050 129454 531398 129486
rect 531050 129218 531106 129454
rect 531342 129218 531398 129454
rect 531050 129134 531398 129218
rect 531050 128898 531106 129134
rect 531342 128898 531398 129134
rect 531050 128866 531398 128898
rect 540286 129454 540646 129486
rect 540286 129218 540348 129454
rect 540584 129218 540646 129454
rect 540286 129134 540646 129218
rect 540286 128898 540348 129134
rect 540584 128898 540646 129134
rect 540286 128866 540646 128898
rect 579020 129454 579380 129486
rect 579020 129218 579082 129454
rect 579318 129218 579380 129454
rect 579020 129134 579380 129218
rect 579020 128898 579082 129134
rect 579318 128898 579380 129134
rect 579020 128866 579380 128898
rect 101304 111454 101664 111486
rect 101304 111218 101366 111454
rect 101602 111218 101664 111454
rect 101304 111134 101664 111218
rect 101304 110898 101366 111134
rect 101602 110898 101664 111134
rect 101304 110866 101664 110898
rect 578300 111454 578660 111486
rect 578300 111218 578362 111454
rect 578598 111218 578660 111454
rect 578300 111134 578660 111218
rect 578300 110898 578362 111134
rect 578598 110898 578660 111134
rect 578300 110866 578660 110898
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 95514 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 96134 97174
rect 95514 96854 96134 96938
rect 95514 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 96134 96854
rect 95514 61174 96134 96618
rect 100584 93454 100944 93486
rect 100584 93218 100646 93454
rect 100882 93218 100944 93454
rect 100584 93134 100944 93218
rect 100584 92898 100646 93134
rect 100882 92898 100944 93134
rect 100584 92866 100944 92898
rect 579020 93454 579380 93486
rect 579020 93218 579082 93454
rect 579318 93218 579380 93454
rect 579020 93134 579380 93218
rect 579020 92898 579082 93134
rect 579318 92898 579380 93134
rect 579020 92866 579380 92898
rect 101304 75454 101664 75486
rect 101304 75218 101366 75454
rect 101602 75218 101664 75454
rect 101304 75134 101664 75218
rect 101304 74898 101366 75134
rect 101602 74898 101664 75134
rect 101304 74866 101664 74898
rect 578300 75454 578660 75486
rect 578300 75218 578362 75454
rect 578598 75218 578660 75454
rect 578300 75134 578660 75218
rect 578300 74898 578362 75134
rect 578598 74898 578660 75134
rect 578300 74866 578660 74898
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 100584 57454 100944 57486
rect 100584 57218 100646 57454
rect 100882 57218 100944 57454
rect 100584 57134 100944 57218
rect 100584 56898 100646 57134
rect 100882 56898 100944 57134
rect 100584 56866 100944 56898
rect 579020 57454 579380 57486
rect 579020 57218 579082 57454
rect 579318 57218 579380 57454
rect 579020 57134 579380 57218
rect 579020 56898 579082 57134
rect 579318 56898 579380 57134
rect 579020 56866 579380 56898
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 28894 99854 48000
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 32614 103574 48000
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 39454 110414 48000
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 43174 114134 48000
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 46894 117854 48000
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 14614 121574 48000
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 21454 128414 48000
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 48000
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 28894 135854 48000
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 32614 139574 48000
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 39454 146414 48000
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 43174 150134 48000
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 46894 153854 48000
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 14614 157574 48000
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 21454 164414 48000
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 25174 168134 48000
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 28894 171854 48000
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 32614 175574 48000
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 39454 182414 48000
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 43174 186134 48000
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 46894 189854 48000
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 14614 193574 48000
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 21454 200414 48000
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 48000
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 28894 207854 48000
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 32614 211574 48000
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 39454 218414 48000
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 43174 222134 48000
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 46894 225854 48000
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 14614 229574 48000
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 21454 236414 48000
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 48000
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 28894 243854 48000
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 32614 247574 48000
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 39454 254414 48000
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 43174 258134 48000
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 46894 261854 48000
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 14614 265574 48000
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 21454 272414 48000
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 25174 276134 48000
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 28894 279854 48000
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 32614 283574 48000
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 39454 290414 48000
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 43174 294134 48000
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 46894 297854 48000
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 14614 301574 48000
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 21454 308414 48000
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 25174 312134 48000
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 28894 315854 48000
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 32614 319574 48000
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 39454 326414 48000
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 43174 330134 48000
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 46894 333854 48000
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 14614 337574 48000
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 21454 344414 48000
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 25174 348134 48000
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 28894 351854 48000
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 32614 355574 48000
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 39454 362414 48000
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 43174 366134 48000
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 46894 369854 48000
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 14614 373574 48000
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 21454 380414 48000
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 25174 384134 48000
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 28894 387854 48000
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 32614 391574 48000
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 39454 398414 48000
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 43174 402134 48000
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 46894 405854 48000
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 14614 409574 48000
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 21454 416414 48000
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 25174 420134 48000
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 28894 423854 48000
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 32614 427574 48000
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 39454 434414 48000
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 43174 438134 48000
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 46894 441854 48000
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 14614 445574 48000
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 21454 452414 48000
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 25174 456134 48000
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 28894 459854 48000
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 32614 463574 48000
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 39454 470414 48000
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 43174 474134 48000
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 46894 477854 48000
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 14614 481574 48000
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 21454 488414 48000
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 25174 492134 48000
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 28894 495854 48000
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 32614 499574 48000
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 39454 506414 48000
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 43174 510134 48000
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 46894 513854 48000
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 14614 517574 48000
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 21454 524414 48000
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 25174 528134 48000
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 28894 531854 48000
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 32614 535574 48000
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 39454 542414 48000
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 43174 546134 48000
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 46894 549854 48000
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 14614 553574 48000
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 21454 560414 48000
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 25174 564134 48000
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 28894 567854 48000
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 32614 571574 48000
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 39454 578414 48000
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 43174 582134 48000
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 66986 104378 67222 104614
rect 67306 104378 67542 104614
rect 66986 104058 67222 104294
rect 67306 104058 67542 104294
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 81266 118658 81502 118894
rect 81586 118658 81822 118894
rect 81266 118338 81502 118574
rect 81586 118338 81822 118574
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 84986 122378 85222 122614
rect 85306 122378 85542 122614
rect 84986 122058 85222 122294
rect 85306 122058 85542 122294
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 578362 543218 578598 543454
rect 578362 542898 578598 543134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 100646 525218 100882 525454
rect 100646 524898 100882 525134
rect 579082 525218 579318 525454
rect 579082 524898 579318 525134
rect 101366 507218 101602 507454
rect 101366 506898 101602 507134
rect 578362 507218 578598 507454
rect 578362 506898 578598 507134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 100646 489218 100882 489454
rect 100646 488898 100882 489134
rect 141860 489218 142096 489454
rect 141860 488898 142096 489134
rect 540348 489218 540584 489454
rect 540348 488898 540584 489134
rect 579082 489218 579318 489454
rect 579082 488898 579318 489134
rect 101366 471218 101602 471454
rect 101366 470898 101602 471134
rect 142580 471218 142816 471454
rect 142580 470898 142816 471134
rect 151346 471218 151582 471454
rect 151346 470898 151582 471134
rect 245050 471218 245286 471454
rect 245050 470898 245286 471134
rect 436722 471218 436958 471454
rect 436722 470898 436958 471134
rect 530426 471218 530662 471454
rect 530426 470898 530662 471134
rect 539628 471218 539864 471454
rect 539628 470898 539864 471134
rect 578362 471218 578598 471454
rect 578362 470898 578598 471134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 100646 453218 100882 453454
rect 100646 452898 100882 453134
rect 141860 453218 142096 453454
rect 141860 452898 142096 453134
rect 150666 453218 150902 453454
rect 150666 452898 150902 453134
rect 245730 453218 245966 453454
rect 245730 452898 245966 453134
rect 436042 453218 436278 453454
rect 436042 452898 436278 453134
rect 531106 453218 531342 453454
rect 531106 452898 531342 453134
rect 540348 453218 540584 453454
rect 540348 452898 540584 453134
rect 579082 453218 579318 453454
rect 579082 452898 579318 453134
rect 101366 435218 101602 435454
rect 101366 434898 101602 435134
rect 142580 435218 142816 435454
rect 142580 434898 142816 435134
rect 151346 435218 151582 435454
rect 151346 434898 151582 435134
rect 245050 435218 245286 435454
rect 245050 434898 245286 435134
rect 436722 435218 436958 435454
rect 436722 434898 436958 435134
rect 530426 435218 530662 435454
rect 530426 434898 530662 435134
rect 539628 435218 539864 435454
rect 539628 434898 539864 435134
rect 578362 435218 578598 435454
rect 578362 434898 578598 435134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 100646 417218 100882 417454
rect 100646 416898 100882 417134
rect 141860 417218 142096 417454
rect 141860 416898 142096 417134
rect 150666 417218 150902 417454
rect 150666 416898 150902 417134
rect 245730 417218 245966 417454
rect 245730 416898 245966 417134
rect 436042 417218 436278 417454
rect 436042 416898 436278 417134
rect 531106 417218 531342 417454
rect 531106 416898 531342 417134
rect 540348 417218 540584 417454
rect 540348 416898 540584 417134
rect 579082 417218 579318 417454
rect 579082 416898 579318 417134
rect 101366 399218 101602 399454
rect 101366 398898 101602 399134
rect 142580 399218 142816 399454
rect 142580 398898 142816 399134
rect 539628 399218 539864 399454
rect 539628 398898 539864 399134
rect 578362 399218 578598 399454
rect 578362 398898 578598 399134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 100646 381218 100882 381454
rect 100646 380898 100882 381134
rect 141860 381218 142096 381454
rect 141860 380898 142096 381134
rect 150666 381218 150902 381454
rect 150666 380898 150902 381134
rect 245730 381218 245966 381454
rect 245730 380898 245966 381134
rect 436042 381218 436278 381454
rect 436042 380898 436278 381134
rect 531106 381218 531342 381454
rect 531106 380898 531342 381134
rect 540348 381218 540584 381454
rect 540348 380898 540584 381134
rect 579082 381218 579318 381454
rect 579082 380898 579318 381134
rect 101366 363218 101602 363454
rect 101366 362898 101602 363134
rect 142580 363218 142816 363454
rect 142580 362898 142816 363134
rect 151346 363218 151582 363454
rect 151346 362898 151582 363134
rect 245050 363218 245286 363454
rect 245050 362898 245286 363134
rect 436722 363218 436958 363454
rect 436722 362898 436958 363134
rect 530426 363218 530662 363454
rect 530426 362898 530662 363134
rect 539628 363218 539864 363454
rect 539628 362898 539864 363134
rect 578362 363218 578598 363454
rect 578362 362898 578598 363134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 100646 345218 100882 345454
rect 100646 344898 100882 345134
rect 141860 345218 142096 345454
rect 141860 344898 142096 345134
rect 150666 345218 150902 345454
rect 150666 344898 150902 345134
rect 245730 345218 245966 345454
rect 245730 344898 245966 345134
rect 436042 345218 436278 345454
rect 436042 344898 436278 345134
rect 531106 345218 531342 345454
rect 531106 344898 531342 345134
rect 540348 345218 540584 345454
rect 540348 344898 540584 345134
rect 579082 345218 579318 345454
rect 579082 344898 579318 345134
rect 101366 327218 101602 327454
rect 101366 326898 101602 327134
rect 142580 327218 142816 327454
rect 142580 326898 142816 327134
rect 151346 327218 151582 327454
rect 151346 326898 151582 327134
rect 245050 327218 245286 327454
rect 245050 326898 245286 327134
rect 436722 327218 436958 327454
rect 436722 326898 436958 327134
rect 530426 327218 530662 327454
rect 530426 326898 530662 327134
rect 539628 327218 539864 327454
rect 539628 326898 539864 327134
rect 578362 327218 578598 327454
rect 578362 326898 578598 327134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 100646 309218 100882 309454
rect 100646 308898 100882 309134
rect 141860 309218 142096 309454
rect 141860 308898 142096 309134
rect 540348 309218 540584 309454
rect 540348 308898 540584 309134
rect 579082 309218 579318 309454
rect 579082 308898 579318 309134
rect 101366 291218 101602 291454
rect 101366 290898 101602 291134
rect 142580 291218 142816 291454
rect 142580 290898 142816 291134
rect 151346 291218 151582 291454
rect 151346 290898 151582 291134
rect 245050 291218 245286 291454
rect 245050 290898 245286 291134
rect 436722 291218 436958 291454
rect 436722 290898 436958 291134
rect 530426 291218 530662 291454
rect 530426 290898 530662 291134
rect 539628 291218 539864 291454
rect 539628 290898 539864 291134
rect 578362 291218 578598 291454
rect 578362 290898 578598 291134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 95546 276938 95782 277174
rect 95866 276938 96102 277174
rect 95546 276618 95782 276854
rect 95866 276618 96102 276854
rect 100646 273218 100882 273454
rect 100646 272898 100882 273134
rect 141860 273218 142096 273454
rect 141860 272898 142096 273134
rect 150666 273218 150902 273454
rect 150666 272898 150902 273134
rect 245730 273218 245966 273454
rect 245730 272898 245966 273134
rect 436042 273218 436278 273454
rect 436042 272898 436278 273134
rect 531106 273218 531342 273454
rect 531106 272898 531342 273134
rect 540348 273218 540584 273454
rect 540348 272898 540584 273134
rect 579082 273218 579318 273454
rect 579082 272898 579318 273134
rect 101366 255218 101602 255454
rect 101366 254898 101602 255134
rect 142580 255218 142816 255454
rect 142580 254898 142816 255134
rect 151346 255218 151582 255454
rect 151346 254898 151582 255134
rect 245050 255218 245286 255454
rect 245050 254898 245286 255134
rect 436722 255218 436958 255454
rect 436722 254898 436958 255134
rect 530426 255218 530662 255454
rect 530426 254898 530662 255134
rect 539628 255218 539864 255454
rect 539628 254898 539864 255134
rect 578362 255218 578598 255454
rect 578362 254898 578598 255134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 95546 240938 95782 241174
rect 95866 240938 96102 241174
rect 95546 240618 95782 240854
rect 95866 240618 96102 240854
rect 100646 237218 100882 237454
rect 100646 236898 100882 237134
rect 141860 237218 142096 237454
rect 141860 236898 142096 237134
rect 150666 237218 150902 237454
rect 150666 236898 150902 237134
rect 245730 237218 245966 237454
rect 245730 236898 245966 237134
rect 436042 237218 436278 237454
rect 436042 236898 436278 237134
rect 531106 237218 531342 237454
rect 531106 236898 531342 237134
rect 540348 237218 540584 237454
rect 540348 236898 540584 237134
rect 579082 237218 579318 237454
rect 579082 236898 579318 237134
rect 101366 219218 101602 219454
rect 101366 218898 101602 219134
rect 142580 219218 142816 219454
rect 142580 218898 142816 219134
rect 436722 219218 436958 219454
rect 436722 218898 436958 219134
rect 530426 219218 530662 219454
rect 530426 218898 530662 219134
rect 539628 219218 539864 219454
rect 539628 218898 539864 219134
rect 578362 219218 578598 219454
rect 578362 218898 578598 219134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 100646 201218 100882 201454
rect 100646 200898 100882 201134
rect 141860 201218 142096 201454
rect 141860 200898 142096 201134
rect 150666 201218 150902 201454
rect 150666 200898 150902 201134
rect 245730 201218 245966 201454
rect 245730 200898 245966 201134
rect 436042 201218 436278 201454
rect 436042 200898 436278 201134
rect 531106 201218 531342 201454
rect 531106 200898 531342 201134
rect 540348 201218 540584 201454
rect 540348 200898 540584 201134
rect 579082 201218 579318 201454
rect 579082 200898 579318 201134
rect 101366 183218 101602 183454
rect 101366 182898 101602 183134
rect 142580 183218 142816 183454
rect 142580 182898 142816 183134
rect 151346 183218 151582 183454
rect 151346 182898 151582 183134
rect 245050 183218 245286 183454
rect 245050 182898 245286 183134
rect 436722 183218 436958 183454
rect 436722 182898 436958 183134
rect 530426 183218 530662 183454
rect 530426 182898 530662 183134
rect 539628 183218 539864 183454
rect 539628 182898 539864 183134
rect 578362 183218 578598 183454
rect 578362 182898 578598 183134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 95546 168938 95782 169174
rect 95866 168938 96102 169174
rect 95546 168618 95782 168854
rect 95866 168618 96102 168854
rect 100646 165218 100882 165454
rect 100646 164898 100882 165134
rect 141860 165218 142096 165454
rect 141860 164898 142096 165134
rect 150666 165218 150902 165454
rect 150666 164898 150902 165134
rect 245730 165218 245966 165454
rect 245730 164898 245966 165134
rect 436042 165218 436278 165454
rect 436042 164898 436278 165134
rect 531106 165218 531342 165454
rect 531106 164898 531342 165134
rect 540348 165218 540584 165454
rect 540348 164898 540584 165134
rect 579082 165218 579318 165454
rect 579082 164898 579318 165134
rect 101366 147218 101602 147454
rect 101366 146898 101602 147134
rect 142580 147218 142816 147454
rect 142580 146898 142816 147134
rect 151346 147218 151582 147454
rect 151346 146898 151582 147134
rect 245050 147218 245286 147454
rect 245050 146898 245286 147134
rect 436722 147218 436958 147454
rect 436722 146898 436958 147134
rect 530426 147218 530662 147454
rect 530426 146898 530662 147134
rect 539628 147218 539864 147454
rect 539628 146898 539864 147134
rect 578362 147218 578598 147454
rect 578362 146898 578598 147134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 95546 132938 95782 133174
rect 95866 132938 96102 133174
rect 95546 132618 95782 132854
rect 95866 132618 96102 132854
rect 100646 129218 100882 129454
rect 100646 128898 100882 129134
rect 141860 129218 142096 129454
rect 141860 128898 142096 129134
rect 150666 129218 150902 129454
rect 150666 128898 150902 129134
rect 245730 129218 245966 129454
rect 245730 128898 245966 129134
rect 436042 129218 436278 129454
rect 436042 128898 436278 129134
rect 531106 129218 531342 129454
rect 531106 128898 531342 129134
rect 540348 129218 540584 129454
rect 540348 128898 540584 129134
rect 579082 129218 579318 129454
rect 579082 128898 579318 129134
rect 101366 111218 101602 111454
rect 101366 110898 101602 111134
rect 578362 111218 578598 111454
rect 578362 110898 578598 111134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 95546 96938 95782 97174
rect 95866 96938 96102 97174
rect 95546 96618 95782 96854
rect 95866 96618 96102 96854
rect 100646 93218 100882 93454
rect 100646 92898 100882 93134
rect 579082 93218 579318 93454
rect 579082 92898 579318 93134
rect 101366 75218 101602 75454
rect 101366 74898 101602 75134
rect 578362 75218 578598 75454
rect 578362 74898 578598 75134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 100646 57218 100882 57454
rect 100646 56898 100882 57134
rect 579082 57218 579318 57454
rect 579082 56898 579318 57134
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 578362 543454
rect 578598 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 578362 543134
rect 578598 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 100646 525454
rect 100882 525218 579082 525454
rect 579318 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 100646 525134
rect 100882 524898 579082 525134
rect 579318 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 101366 507454
rect 101602 507218 578362 507454
rect 578598 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 101366 507134
rect 101602 506898 578362 507134
rect 578598 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 100646 489454
rect 100882 489218 141860 489454
rect 142096 489218 540348 489454
rect 540584 489218 579082 489454
rect 579318 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 100646 489134
rect 100882 488898 141860 489134
rect 142096 488898 540348 489134
rect 540584 488898 579082 489134
rect 579318 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 101366 471454
rect 101602 471218 142580 471454
rect 142816 471218 151346 471454
rect 151582 471218 245050 471454
rect 245286 471218 436722 471454
rect 436958 471218 530426 471454
rect 530662 471218 539628 471454
rect 539864 471218 578362 471454
rect 578598 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 101366 471134
rect 101602 470898 142580 471134
rect 142816 470898 151346 471134
rect 151582 470898 245050 471134
rect 245286 470898 436722 471134
rect 436958 470898 530426 471134
rect 530662 470898 539628 471134
rect 539864 470898 578362 471134
rect 578598 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 100646 453454
rect 100882 453218 141860 453454
rect 142096 453218 150666 453454
rect 150902 453218 245730 453454
rect 245966 453218 436042 453454
rect 436278 453218 531106 453454
rect 531342 453218 540348 453454
rect 540584 453218 579082 453454
rect 579318 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 100646 453134
rect 100882 452898 141860 453134
rect 142096 452898 150666 453134
rect 150902 452898 245730 453134
rect 245966 452898 436042 453134
rect 436278 452898 531106 453134
rect 531342 452898 540348 453134
rect 540584 452898 579082 453134
rect 579318 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 101366 435454
rect 101602 435218 142580 435454
rect 142816 435218 151346 435454
rect 151582 435218 245050 435454
rect 245286 435218 436722 435454
rect 436958 435218 530426 435454
rect 530662 435218 539628 435454
rect 539864 435218 578362 435454
rect 578598 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 101366 435134
rect 101602 434898 142580 435134
rect 142816 434898 151346 435134
rect 151582 434898 245050 435134
rect 245286 434898 436722 435134
rect 436958 434898 530426 435134
rect 530662 434898 539628 435134
rect 539864 434898 578362 435134
rect 578598 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 100646 417454
rect 100882 417218 141860 417454
rect 142096 417218 150666 417454
rect 150902 417218 245730 417454
rect 245966 417218 436042 417454
rect 436278 417218 531106 417454
rect 531342 417218 540348 417454
rect 540584 417218 579082 417454
rect 579318 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 100646 417134
rect 100882 416898 141860 417134
rect 142096 416898 150666 417134
rect 150902 416898 245730 417134
rect 245966 416898 436042 417134
rect 436278 416898 531106 417134
rect 531342 416898 540348 417134
rect 540584 416898 579082 417134
rect 579318 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 101366 399454
rect 101602 399218 142580 399454
rect 142816 399218 539628 399454
rect 539864 399218 578362 399454
rect 578598 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 101366 399134
rect 101602 398898 142580 399134
rect 142816 398898 539628 399134
rect 539864 398898 578362 399134
rect 578598 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 100646 381454
rect 100882 381218 141860 381454
rect 142096 381218 150666 381454
rect 150902 381218 245730 381454
rect 245966 381218 436042 381454
rect 436278 381218 531106 381454
rect 531342 381218 540348 381454
rect 540584 381218 579082 381454
rect 579318 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 100646 381134
rect 100882 380898 141860 381134
rect 142096 380898 150666 381134
rect 150902 380898 245730 381134
rect 245966 380898 436042 381134
rect 436278 380898 531106 381134
rect 531342 380898 540348 381134
rect 540584 380898 579082 381134
rect 579318 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 101366 363454
rect 101602 363218 142580 363454
rect 142816 363218 151346 363454
rect 151582 363218 245050 363454
rect 245286 363218 436722 363454
rect 436958 363218 530426 363454
rect 530662 363218 539628 363454
rect 539864 363218 578362 363454
rect 578598 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 101366 363134
rect 101602 362898 142580 363134
rect 142816 362898 151346 363134
rect 151582 362898 245050 363134
rect 245286 362898 436722 363134
rect 436958 362898 530426 363134
rect 530662 362898 539628 363134
rect 539864 362898 578362 363134
rect 578598 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 100646 345454
rect 100882 345218 141860 345454
rect 142096 345218 150666 345454
rect 150902 345218 245730 345454
rect 245966 345218 436042 345454
rect 436278 345218 531106 345454
rect 531342 345218 540348 345454
rect 540584 345218 579082 345454
rect 579318 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 100646 345134
rect 100882 344898 141860 345134
rect 142096 344898 150666 345134
rect 150902 344898 245730 345134
rect 245966 344898 436042 345134
rect 436278 344898 531106 345134
rect 531342 344898 540348 345134
rect 540584 344898 579082 345134
rect 579318 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 101366 327454
rect 101602 327218 142580 327454
rect 142816 327218 151346 327454
rect 151582 327218 245050 327454
rect 245286 327218 436722 327454
rect 436958 327218 530426 327454
rect 530662 327218 539628 327454
rect 539864 327218 578362 327454
rect 578598 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 101366 327134
rect 101602 326898 142580 327134
rect 142816 326898 151346 327134
rect 151582 326898 245050 327134
rect 245286 326898 436722 327134
rect 436958 326898 530426 327134
rect 530662 326898 539628 327134
rect 539864 326898 578362 327134
rect 578598 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 100646 309454
rect 100882 309218 141860 309454
rect 142096 309218 540348 309454
rect 540584 309218 579082 309454
rect 579318 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 100646 309134
rect 100882 308898 141860 309134
rect 142096 308898 540348 309134
rect 540584 308898 579082 309134
rect 579318 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 101366 291454
rect 101602 291218 142580 291454
rect 142816 291218 151346 291454
rect 151582 291218 245050 291454
rect 245286 291218 436722 291454
rect 436958 291218 530426 291454
rect 530662 291218 539628 291454
rect 539864 291218 578362 291454
rect 578598 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 101366 291134
rect 101602 290898 142580 291134
rect 142816 290898 151346 291134
rect 151582 290898 245050 291134
rect 245286 290898 436722 291134
rect 436958 290898 530426 291134
rect 530662 290898 539628 291134
rect 539864 290898 578362 291134
rect 578598 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 100646 273454
rect 100882 273218 141860 273454
rect 142096 273218 150666 273454
rect 150902 273218 245730 273454
rect 245966 273218 436042 273454
rect 436278 273218 531106 273454
rect 531342 273218 540348 273454
rect 540584 273218 579082 273454
rect 579318 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 100646 273134
rect 100882 272898 141860 273134
rect 142096 272898 150666 273134
rect 150902 272898 245730 273134
rect 245966 272898 436042 273134
rect 436278 272898 531106 273134
rect 531342 272898 540348 273134
rect 540584 272898 579082 273134
rect 579318 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 101366 255454
rect 101602 255218 142580 255454
rect 142816 255218 151346 255454
rect 151582 255218 245050 255454
rect 245286 255218 436722 255454
rect 436958 255218 530426 255454
rect 530662 255218 539628 255454
rect 539864 255218 578362 255454
rect 578598 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 101366 255134
rect 101602 254898 142580 255134
rect 142816 254898 151346 255134
rect 151582 254898 245050 255134
rect 245286 254898 436722 255134
rect 436958 254898 530426 255134
rect 530662 254898 539628 255134
rect 539864 254898 578362 255134
rect 578598 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 100646 237454
rect 100882 237218 141860 237454
rect 142096 237218 150666 237454
rect 150902 237218 245730 237454
rect 245966 237218 436042 237454
rect 436278 237218 531106 237454
rect 531342 237218 540348 237454
rect 540584 237218 579082 237454
rect 579318 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 100646 237134
rect 100882 236898 141860 237134
rect 142096 236898 150666 237134
rect 150902 236898 245730 237134
rect 245966 236898 436042 237134
rect 436278 236898 531106 237134
rect 531342 236898 540348 237134
rect 540584 236898 579082 237134
rect 579318 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 101366 219454
rect 101602 219218 142580 219454
rect 142816 219218 436722 219454
rect 436958 219218 530426 219454
rect 530662 219218 539628 219454
rect 539864 219218 578362 219454
rect 578598 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 101366 219134
rect 101602 218898 142580 219134
rect 142816 218898 436722 219134
rect 436958 218898 530426 219134
rect 530662 218898 539628 219134
rect 539864 218898 578362 219134
rect 578598 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 100646 201454
rect 100882 201218 141860 201454
rect 142096 201218 150666 201454
rect 150902 201218 245730 201454
rect 245966 201218 436042 201454
rect 436278 201218 531106 201454
rect 531342 201218 540348 201454
rect 540584 201218 579082 201454
rect 579318 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 100646 201134
rect 100882 200898 141860 201134
rect 142096 200898 150666 201134
rect 150902 200898 245730 201134
rect 245966 200898 436042 201134
rect 436278 200898 531106 201134
rect 531342 200898 540348 201134
rect 540584 200898 579082 201134
rect 579318 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 101366 183454
rect 101602 183218 142580 183454
rect 142816 183218 151346 183454
rect 151582 183218 245050 183454
rect 245286 183218 436722 183454
rect 436958 183218 530426 183454
rect 530662 183218 539628 183454
rect 539864 183218 578362 183454
rect 578598 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 101366 183134
rect 101602 182898 142580 183134
rect 142816 182898 151346 183134
rect 151582 182898 245050 183134
rect 245286 182898 436722 183134
rect 436958 182898 530426 183134
rect 530662 182898 539628 183134
rect 539864 182898 578362 183134
rect 578598 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 100646 165454
rect 100882 165218 141860 165454
rect 142096 165218 150666 165454
rect 150902 165218 245730 165454
rect 245966 165218 436042 165454
rect 436278 165218 531106 165454
rect 531342 165218 540348 165454
rect 540584 165218 579082 165454
rect 579318 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 100646 165134
rect 100882 164898 141860 165134
rect 142096 164898 150666 165134
rect 150902 164898 245730 165134
rect 245966 164898 436042 165134
rect 436278 164898 531106 165134
rect 531342 164898 540348 165134
rect 540584 164898 579082 165134
rect 579318 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 101366 147454
rect 101602 147218 142580 147454
rect 142816 147218 151346 147454
rect 151582 147218 245050 147454
rect 245286 147218 436722 147454
rect 436958 147218 530426 147454
rect 530662 147218 539628 147454
rect 539864 147218 578362 147454
rect 578598 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 101366 147134
rect 101602 146898 142580 147134
rect 142816 146898 151346 147134
rect 151582 146898 245050 147134
rect 245286 146898 436722 147134
rect 436958 146898 530426 147134
rect 530662 146898 539628 147134
rect 539864 146898 578362 147134
rect 578598 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 100646 129454
rect 100882 129218 141860 129454
rect 142096 129218 150666 129454
rect 150902 129218 245730 129454
rect 245966 129218 436042 129454
rect 436278 129218 531106 129454
rect 531342 129218 540348 129454
rect 540584 129218 579082 129454
rect 579318 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 100646 129134
rect 100882 128898 141860 129134
rect 142096 128898 150666 129134
rect 150902 128898 245730 129134
rect 245966 128898 436042 129134
rect 436278 128898 531106 129134
rect 531342 128898 540348 129134
rect 540584 128898 579082 129134
rect 579318 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 101366 111454
rect 101602 111218 578362 111454
rect 578598 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 101366 111134
rect 101602 110898 578362 111134
rect 578598 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 100646 93454
rect 100882 93218 579082 93454
rect 579318 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 100646 93134
rect 100882 92898 579082 93134
rect 579318 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 101366 75454
rect 101602 75218 578362 75454
rect 578598 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 101366 75134
rect 101602 74898 578362 75134
rect 578598 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 100646 57454
rect 100882 57218 579082 57454
rect 579318 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 100646 57134
rect 100882 56898 579082 57134
rect 579318 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use azadi_soc_top_caravel  mprj
timestamp 0
transform 1 0 100000 0 1 50000
box 0 0 479964 500004
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 692052 480 692292 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 598212 480 598452 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 504372 480 504612 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 410532 480 410772 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 316556 480 316796 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 222716 480 222956 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 15 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 16 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 17 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 18 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 19 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 20 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 21 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 23 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 24 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 25 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 26 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 27 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 28 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 29 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 30 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 31 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 32 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 33 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 34 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 35 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 36 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 37 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 38 nsew signal input
rlabel metal3 s -960 668524 480 668764 4 io_in[24]
port 39 nsew signal input
rlabel metal3 s -960 574684 480 574924 4 io_in[25]
port 40 nsew signal input
rlabel metal3 s -960 480844 480 481084 4 io_in[26]
port 41 nsew signal input
rlabel metal3 s -960 387004 480 387244 4 io_in[27]
port 42 nsew signal input
rlabel metal3 s -960 293164 480 293404 4 io_in[28]
port 43 nsew signal input
rlabel metal3 s -960 199324 480 199564 4 io_in[29]
port 44 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 45 nsew signal input
rlabel metal3 s -960 128876 480 129116 4 io_in[30]
port 46 nsew signal input
rlabel metal3 s -960 58564 480 58804 4 io_in[31]
port 47 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 48 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 49 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 50 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 51 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 52 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 53 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 54 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 55 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 56 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 57 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 58 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 59 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 60 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 61 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 62 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 63 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 64 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 65 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 66 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 67 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 68 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 69 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 70 nsew signal tristate
rlabel metal3 s -960 621604 480 621844 4 io_oeb[24]
port 71 nsew signal tristate
rlabel metal3 s -960 527764 480 528004 4 io_oeb[25]
port 72 nsew signal tristate
rlabel metal3 s -960 433924 480 434164 4 io_oeb[26]
port 73 nsew signal tristate
rlabel metal3 s -960 340084 480 340324 4 io_oeb[27]
port 74 nsew signal tristate
rlabel metal3 s -960 246244 480 246484 4 io_oeb[28]
port 75 nsew signal tristate
rlabel metal3 s -960 152404 480 152644 4 io_oeb[29]
port 76 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 77 nsew signal tristate
rlabel metal3 s -960 81956 480 82196 4 io_oeb[30]
port 78 nsew signal tristate
rlabel metal3 s -960 11644 480 11884 4 io_oeb[31]
port 79 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 80 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 81 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 82 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 83 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 84 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 85 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 86 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 87 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 88 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 89 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 90 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 91 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 92 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 93 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 94 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 95 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 96 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 97 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 98 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 99 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 100 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 101 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 102 nsew signal tristate
rlabel metal3 s -960 645132 480 645372 4 io_out[24]
port 103 nsew signal tristate
rlabel metal3 s -960 551292 480 551532 4 io_out[25]
port 104 nsew signal tristate
rlabel metal3 s -960 457452 480 457692 4 io_out[26]
port 105 nsew signal tristate
rlabel metal3 s -960 363612 480 363852 4 io_out[27]
port 106 nsew signal tristate
rlabel metal3 s -960 269636 480 269876 4 io_out[28]
port 107 nsew signal tristate
rlabel metal3 s -960 175796 480 176036 4 io_out[29]
port 108 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 109 nsew signal tristate
rlabel metal3 s -960 105484 480 105724 4 io_out[30]
port 110 nsew signal tristate
rlabel metal3 s -960 35036 480 35276 4 io_out[31]
port 111 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 112 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 113 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 114 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 115 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 116 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 117 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 118 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 119 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 120 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 121 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 122 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 123 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 124 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 125 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 126 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 127 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 128 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 129 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 130 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 131 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 132 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 133 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 134 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 135 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 136 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 137 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 138 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 139 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 140 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 141 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 142 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 143 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 144 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 145 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 146 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 147 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 148 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 149 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 150 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 151 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 152 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 153 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 154 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 155 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 156 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 157 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 158 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 159 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 160 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 161 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 162 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 163 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 164 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 165 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 166 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 167 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 168 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 169 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 170 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 171 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 172 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 173 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 174 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 175 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 176 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 177 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 178 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 179 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 180 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 181 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 182 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 183 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 184 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 185 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 186 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 187 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 188 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 189 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 190 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 191 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 192 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 193 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 194 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 195 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 196 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 197 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 198 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 199 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 200 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 201 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 202 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 203 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 204 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 205 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 206 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 207 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 208 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 209 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 210 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 211 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 212 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 213 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 214 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 215 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 216 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 217 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 218 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 219 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 220 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 221 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 222 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 223 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 224 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 225 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 226 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 227 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 228 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 229 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 230 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 231 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 232 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 233 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 234 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 235 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 236 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 237 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 238 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 239 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 240 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 241 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 242 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 243 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 244 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 245 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 246 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 247 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 248 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 249 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 250 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 251 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 252 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 253 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 254 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 255 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 256 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 257 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 258 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 259 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 260 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 261 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 262 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 263 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 264 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 265 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 266 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 267 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 268 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 269 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 270 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 271 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 272 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 273 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 274 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 275 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 276 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 277 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 278 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 279 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 280 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 281 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 282 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 283 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 284 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 285 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 286 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 287 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 288 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 289 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 290 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 291 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 292 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 293 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 294 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 295 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 296 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 297 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 298 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 299 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 300 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 301 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 302 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 303 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 304 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 305 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 306 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 307 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 308 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 309 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 310 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 311 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 312 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 313 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 314 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 315 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 316 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 317 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 318 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 319 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 320 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 321 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 322 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 323 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 324 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 325 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 326 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 327 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 328 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 329 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 330 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 331 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 332 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 333 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 334 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 335 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 336 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 337 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 338 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 339 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 340 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 341 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 342 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 343 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 344 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 345 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 346 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 347 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 348 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 349 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 350 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 351 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 352 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 353 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 354 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 355 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 356 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 357 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 358 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 359 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 360 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 361 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 362 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 363 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 364 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 365 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 366 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 367 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 368 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 369 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 370 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 371 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 372 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 373 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 374 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 375 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 376 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 377 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 378 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 379 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 380 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 381 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 382 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 383 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 384 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 385 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 386 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 387 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 388 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 389 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 390 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 391 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 392 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 393 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 394 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 395 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 396 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 397 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 398 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 399 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 400 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 401 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 402 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 403 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 404 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 405 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 406 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 407 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 408 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 409 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 410 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 411 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 412 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 413 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 414 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 415 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 416 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 417 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 418 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 419 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 420 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 421 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 422 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 423 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 424 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 425 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 426 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 427 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 428 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 429 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 430 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 431 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 432 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 433 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 434 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 435 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 436 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 437 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 438 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 439 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 440 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 441 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 442 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 443 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 444 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 445 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 446 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 447 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 448 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 449 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 450 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 451 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 452 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 453 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 454 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 455 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 456 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 457 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 458 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 459 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 460 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 461 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 462 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 463 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 464 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 465 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 466 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 467 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 468 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 469 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 470 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 471 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 472 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 473 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 474 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 475 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 476 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 477 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 478 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 479 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 480 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 481 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 482 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 483 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 484 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 485 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 486 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 487 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 488 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 489 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 490 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 491 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 492 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 493 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 494 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 495 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 496 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 497 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 498 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 499 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 500 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 501 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 502 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 503 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 504 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 505 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 506 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 507 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 507 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 507 nsew power input
rlabel metal4 s 109794 -1894 110414 48000 6 vccd1
port 507 nsew power input
rlabel metal4 s 145794 -1894 146414 48000 6 vccd1
port 507 nsew power input
rlabel metal4 s 181794 -1894 182414 48000 6 vccd1
port 507 nsew power input
rlabel metal4 s 217794 -1894 218414 48000 6 vccd1
port 507 nsew power input
rlabel metal4 s 253794 -1894 254414 48000 6 vccd1
port 507 nsew power input
rlabel metal4 s 289794 -1894 290414 48000 6 vccd1
port 507 nsew power input
rlabel metal4 s 325794 -1894 326414 48000 6 vccd1
port 507 nsew power input
rlabel metal4 s 361794 -1894 362414 48000 6 vccd1
port 507 nsew power input
rlabel metal4 s 397794 -1894 398414 48000 6 vccd1
port 507 nsew power input
rlabel metal4 s 433794 -1894 434414 48000 6 vccd1
port 507 nsew power input
rlabel metal4 s 469794 -1894 470414 48000 6 vccd1
port 507 nsew power input
rlabel metal4 s 505794 -1894 506414 48000 6 vccd1
port 507 nsew power input
rlabel metal4 s 541794 -1894 542414 48000 6 vccd1
port 507 nsew power input
rlabel metal4 s 577794 -1894 578414 48000 6 vccd1
port 507 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 507 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 507 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 73794 -1894 74414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 109794 552004 110414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 145794 552004 146414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 181794 552004 182414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 217794 552004 218414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 253794 552004 254414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 289794 552004 290414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 325794 552004 326414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 361794 552004 362414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 397794 552004 398414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 433794 552004 434414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 469794 552004 470414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 505794 552004 506414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 541794 552004 542414 705830 6 vccd1
port 507 nsew power input
rlabel metal4 s 577794 552004 578414 705830 6 vccd1
port 507 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 508 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 508 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 508 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 508 nsew power input
rlabel metal4 s 113514 -3814 114134 48000 6 vccd2
port 508 nsew power input
rlabel metal4 s 149514 -3814 150134 48000 6 vccd2
port 508 nsew power input
rlabel metal4 s 185514 -3814 186134 48000 6 vccd2
port 508 nsew power input
rlabel metal4 s 221514 -3814 222134 48000 6 vccd2
port 508 nsew power input
rlabel metal4 s 257514 -3814 258134 48000 6 vccd2
port 508 nsew power input
rlabel metal4 s 293514 -3814 294134 48000 6 vccd2
port 508 nsew power input
rlabel metal4 s 329514 -3814 330134 48000 6 vccd2
port 508 nsew power input
rlabel metal4 s 365514 -3814 366134 48000 6 vccd2
port 508 nsew power input
rlabel metal4 s 401514 -3814 402134 48000 6 vccd2
port 508 nsew power input
rlabel metal4 s 437514 -3814 438134 48000 6 vccd2
port 508 nsew power input
rlabel metal4 s 473514 -3814 474134 48000 6 vccd2
port 508 nsew power input
rlabel metal4 s 509514 -3814 510134 48000 6 vccd2
port 508 nsew power input
rlabel metal4 s 545514 -3814 546134 48000 6 vccd2
port 508 nsew power input
rlabel metal4 s 581514 -3814 582134 48000 6 vccd2
port 508 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 508 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 508 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 77514 -3814 78134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 113514 552004 114134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 149514 552004 150134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 185514 552004 186134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 221514 552004 222134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 257514 552004 258134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 293514 552004 294134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 329514 552004 330134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 365514 552004 366134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 401514 552004 402134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 437514 552004 438134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 473514 552004 474134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 509514 552004 510134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 545514 552004 546134 707750 6 vccd2
port 508 nsew power input
rlabel metal4 s 581514 552004 582134 707750 6 vccd2
port 508 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 509 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 509 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 509 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 509 nsew power input
rlabel metal4 s 117234 -5734 117854 48000 6 vdda1
port 509 nsew power input
rlabel metal4 s 153234 -5734 153854 48000 6 vdda1
port 509 nsew power input
rlabel metal4 s 189234 -5734 189854 48000 6 vdda1
port 509 nsew power input
rlabel metal4 s 225234 -5734 225854 48000 6 vdda1
port 509 nsew power input
rlabel metal4 s 261234 -5734 261854 48000 6 vdda1
port 509 nsew power input
rlabel metal4 s 297234 -5734 297854 48000 6 vdda1
port 509 nsew power input
rlabel metal4 s 333234 -5734 333854 48000 6 vdda1
port 509 nsew power input
rlabel metal4 s 369234 -5734 369854 48000 6 vdda1
port 509 nsew power input
rlabel metal4 s 405234 -5734 405854 48000 6 vdda1
port 509 nsew power input
rlabel metal4 s 441234 -5734 441854 48000 6 vdda1
port 509 nsew power input
rlabel metal4 s 477234 -5734 477854 48000 6 vdda1
port 509 nsew power input
rlabel metal4 s 513234 -5734 513854 48000 6 vdda1
port 509 nsew power input
rlabel metal4 s 549234 -5734 549854 48000 6 vdda1
port 509 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 509 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 509 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 81234 -5734 81854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 117234 552004 117854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 153234 552004 153854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 189234 552004 189854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 225234 552004 225854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 261234 552004 261854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 297234 552004 297854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 333234 552004 333854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 369234 552004 369854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 405234 552004 405854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 441234 552004 441854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 477234 552004 477854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 513234 552004 513854 709670 6 vdda1
port 509 nsew power input
rlabel metal4 s 549234 552004 549854 709670 6 vdda1
port 509 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 510 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 510 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 510 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 510 nsew power input
rlabel metal4 s 120954 -7654 121574 48000 6 vdda2
port 510 nsew power input
rlabel metal4 s 156954 -7654 157574 48000 6 vdda2
port 510 nsew power input
rlabel metal4 s 192954 -7654 193574 48000 6 vdda2
port 510 nsew power input
rlabel metal4 s 228954 -7654 229574 48000 6 vdda2
port 510 nsew power input
rlabel metal4 s 264954 -7654 265574 48000 6 vdda2
port 510 nsew power input
rlabel metal4 s 300954 -7654 301574 48000 6 vdda2
port 510 nsew power input
rlabel metal4 s 336954 -7654 337574 48000 6 vdda2
port 510 nsew power input
rlabel metal4 s 372954 -7654 373574 48000 6 vdda2
port 510 nsew power input
rlabel metal4 s 408954 -7654 409574 48000 6 vdda2
port 510 nsew power input
rlabel metal4 s 444954 -7654 445574 48000 6 vdda2
port 510 nsew power input
rlabel metal4 s 480954 -7654 481574 48000 6 vdda2
port 510 nsew power input
rlabel metal4 s 516954 -7654 517574 48000 6 vdda2
port 510 nsew power input
rlabel metal4 s 552954 -7654 553574 48000 6 vdda2
port 510 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 510 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 510 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 84954 -7654 85574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 120954 552004 121574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 156954 552004 157574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 192954 552004 193574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 228954 552004 229574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 264954 552004 265574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 300954 552004 301574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 336954 552004 337574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 372954 552004 373574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 408954 552004 409574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 444954 552004 445574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 480954 552004 481574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 516954 552004 517574 711590 6 vdda2
port 510 nsew power input
rlabel metal4 s 552954 552004 553574 711590 6 vdda2
port 510 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 511 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 99234 -5734 99854 48000 6 vssa1
port 511 nsew ground input
rlabel metal4 s 135234 -5734 135854 48000 6 vssa1
port 511 nsew ground input
rlabel metal4 s 171234 -5734 171854 48000 6 vssa1
port 511 nsew ground input
rlabel metal4 s 207234 -5734 207854 48000 6 vssa1
port 511 nsew ground input
rlabel metal4 s 243234 -5734 243854 48000 6 vssa1
port 511 nsew ground input
rlabel metal4 s 279234 -5734 279854 48000 6 vssa1
port 511 nsew ground input
rlabel metal4 s 315234 -5734 315854 48000 6 vssa1
port 511 nsew ground input
rlabel metal4 s 351234 -5734 351854 48000 6 vssa1
port 511 nsew ground input
rlabel metal4 s 387234 -5734 387854 48000 6 vssa1
port 511 nsew ground input
rlabel metal4 s 423234 -5734 423854 48000 6 vssa1
port 511 nsew ground input
rlabel metal4 s 459234 -5734 459854 48000 6 vssa1
port 511 nsew ground input
rlabel metal4 s 495234 -5734 495854 48000 6 vssa1
port 511 nsew ground input
rlabel metal4 s 531234 -5734 531854 48000 6 vssa1
port 511 nsew ground input
rlabel metal4 s 567234 -5734 567854 48000 6 vssa1
port 511 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 511 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 99234 552004 99854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 135234 552004 135854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 171234 552004 171854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 207234 552004 207854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 243234 552004 243854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 279234 552004 279854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 315234 552004 315854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 351234 552004 351854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 387234 552004 387854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 423234 552004 423854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 459234 552004 459854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 495234 552004 495854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 531234 552004 531854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 567234 552004 567854 709670 6 vssa1
port 511 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 511 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 512 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 102954 -7654 103574 48000 6 vssa2
port 512 nsew ground input
rlabel metal4 s 138954 -7654 139574 48000 6 vssa2
port 512 nsew ground input
rlabel metal4 s 174954 -7654 175574 48000 6 vssa2
port 512 nsew ground input
rlabel metal4 s 210954 -7654 211574 48000 6 vssa2
port 512 nsew ground input
rlabel metal4 s 246954 -7654 247574 48000 6 vssa2
port 512 nsew ground input
rlabel metal4 s 282954 -7654 283574 48000 6 vssa2
port 512 nsew ground input
rlabel metal4 s 318954 -7654 319574 48000 6 vssa2
port 512 nsew ground input
rlabel metal4 s 354954 -7654 355574 48000 6 vssa2
port 512 nsew ground input
rlabel metal4 s 390954 -7654 391574 48000 6 vssa2
port 512 nsew ground input
rlabel metal4 s 426954 -7654 427574 48000 6 vssa2
port 512 nsew ground input
rlabel metal4 s 462954 -7654 463574 48000 6 vssa2
port 512 nsew ground input
rlabel metal4 s 498954 -7654 499574 48000 6 vssa2
port 512 nsew ground input
rlabel metal4 s 534954 -7654 535574 48000 6 vssa2
port 512 nsew ground input
rlabel metal4 s 570954 -7654 571574 48000 6 vssa2
port 512 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 512 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 66954 -7654 67574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 102954 552004 103574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 138954 552004 139574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 174954 552004 175574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 210954 552004 211574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 246954 552004 247574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 282954 552004 283574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 318954 552004 319574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 354954 552004 355574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 390954 552004 391574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 426954 552004 427574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 462954 552004 463574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 498954 552004 499574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 534954 552004 535574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 570954 552004 571574 711590 6 vssa2
port 512 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 512 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 513 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 127794 -1894 128414 48000 6 vssd1
port 513 nsew ground input
rlabel metal4 s 163794 -1894 164414 48000 6 vssd1
port 513 nsew ground input
rlabel metal4 s 199794 -1894 200414 48000 6 vssd1
port 513 nsew ground input
rlabel metal4 s 235794 -1894 236414 48000 6 vssd1
port 513 nsew ground input
rlabel metal4 s 271794 -1894 272414 48000 6 vssd1
port 513 nsew ground input
rlabel metal4 s 307794 -1894 308414 48000 6 vssd1
port 513 nsew ground input
rlabel metal4 s 343794 -1894 344414 48000 6 vssd1
port 513 nsew ground input
rlabel metal4 s 379794 -1894 380414 48000 6 vssd1
port 513 nsew ground input
rlabel metal4 s 415794 -1894 416414 48000 6 vssd1
port 513 nsew ground input
rlabel metal4 s 451794 -1894 452414 48000 6 vssd1
port 513 nsew ground input
rlabel metal4 s 487794 -1894 488414 48000 6 vssd1
port 513 nsew ground input
rlabel metal4 s 523794 -1894 524414 48000 6 vssd1
port 513 nsew ground input
rlabel metal4 s 559794 -1894 560414 48000 6 vssd1
port 513 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 513 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 91794 -1894 92414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 127794 552004 128414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 163794 552004 164414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 199794 552004 200414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 235794 552004 236414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 271794 552004 272414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 307794 552004 308414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 343794 552004 344414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 379794 552004 380414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 415794 552004 416414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 451794 552004 452414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 487794 552004 488414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 523794 552004 524414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 559794 552004 560414 705830 6 vssd1
port 513 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 513 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 514 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 131514 -3814 132134 48000 6 vssd2
port 514 nsew ground input
rlabel metal4 s 167514 -3814 168134 48000 6 vssd2
port 514 nsew ground input
rlabel metal4 s 203514 -3814 204134 48000 6 vssd2
port 514 nsew ground input
rlabel metal4 s 239514 -3814 240134 48000 6 vssd2
port 514 nsew ground input
rlabel metal4 s 275514 -3814 276134 48000 6 vssd2
port 514 nsew ground input
rlabel metal4 s 311514 -3814 312134 48000 6 vssd2
port 514 nsew ground input
rlabel metal4 s 347514 -3814 348134 48000 6 vssd2
port 514 nsew ground input
rlabel metal4 s 383514 -3814 384134 48000 6 vssd2
port 514 nsew ground input
rlabel metal4 s 419514 -3814 420134 48000 6 vssd2
port 514 nsew ground input
rlabel metal4 s 455514 -3814 456134 48000 6 vssd2
port 514 nsew ground input
rlabel metal4 s 491514 -3814 492134 48000 6 vssd2
port 514 nsew ground input
rlabel metal4 s 527514 -3814 528134 48000 6 vssd2
port 514 nsew ground input
rlabel metal4 s 563514 -3814 564134 48000 6 vssd2
port 514 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 514 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 95514 -3814 96134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 131514 552004 132134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 167514 552004 168134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 203514 552004 204134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 239514 552004 240134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 275514 552004 276134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 311514 552004 312134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 347514 552004 348134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 383514 552004 384134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 419514 552004 420134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 455514 552004 456134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 491514 552004 492134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 527514 552004 528134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 563514 552004 564134 707750 6 vssd2
port 514 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 514 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 515 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 516 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 517 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 518 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 519 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 520 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 521 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 522 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 523 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 524 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 525 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 526 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 527 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 528 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 529 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 530 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 531 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 532 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 533 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 534 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 535 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 536 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 537 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 538 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 539 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 540 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 541 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 542 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 543 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 544 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 545 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 546 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 547 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 548 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 549 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 550 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 551 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 552 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 553 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 554 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 555 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 556 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 557 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 558 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 559 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 560 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 561 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 562 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 563 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 564 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 565 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 566 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 567 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 568 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 569 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 570 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 571 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 572 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 573 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 574 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 575 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 576 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 577 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 578 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 579 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 580 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 581 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 582 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 583 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 584 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 585 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 586 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 587 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 588 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 589 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 590 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 591 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 592 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 593 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 594 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 595 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 596 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 597 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 598 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 599 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 600 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 601 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 602 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 603 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 604 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 605 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 606 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 607 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 608 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 609 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 610 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 611 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 612 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 613 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 614 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 615 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 616 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 617 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 618 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 619 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 620 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
