magic
tech sky130A
magscale 1 2
timestamp 1654458627
<< metal1 >>
rect 1394 386384 1400 386436
rect 1452 386424 1458 386436
rect 57606 386424 57612 386436
rect 1452 386396 57612 386424
rect 1452 386384 1458 386396
rect 57606 386384 57612 386396
rect 57664 386384 57670 386436
rect 372154 59780 372160 59832
rect 372212 59820 372218 59832
rect 373718 59820 373724 59832
rect 372212 59792 373724 59820
rect 372212 59780 372218 59792
rect 373718 59780 373724 59792
rect 373776 59780 373782 59832
rect 430114 59780 430120 59832
rect 430172 59820 430178 59832
rect 431494 59820 431500 59832
rect 430172 59792 431500 59820
rect 430172 59780 430178 59792
rect 431494 59780 431500 59792
rect 431552 59780 431558 59832
rect 488074 59780 488080 59832
rect 488132 59820 488138 59832
rect 489362 59820 489368 59832
rect 488132 59792 489368 59820
rect 488132 59780 488138 59792
rect 489362 59780 489368 59792
rect 489420 59780 489426 59832
rect 498470 59780 498476 59832
rect 498528 59820 498534 59832
rect 499482 59820 499488 59832
rect 498528 59792 499488 59820
rect 498528 59780 498534 59792
rect 499482 59780 499488 59792
rect 499540 59780 499546 59832
rect 516962 59780 516968 59832
rect 517020 59820 517026 59832
rect 518342 59820 518348 59832
rect 517020 59792 518348 59820
rect 517020 59780 517026 59792
rect 518342 59780 518348 59792
rect 518400 59780 518406 59832
rect 73062 59712 73068 59764
rect 73120 59752 73126 59764
rect 74718 59752 74724 59764
rect 73120 59724 74724 59752
rect 73120 59712 73126 59724
rect 74718 59712 74724 59724
rect 74776 59712 74782 59764
rect 77938 59712 77944 59764
rect 77996 59752 78002 59764
rect 79870 59752 79876 59764
rect 77996 59724 79876 59752
rect 77996 59712 78002 59724
rect 79870 59712 79876 59724
rect 79928 59712 79934 59764
rect 80698 59712 80704 59764
rect 80756 59752 80762 59764
rect 82998 59752 83004 59764
rect 80756 59724 83004 59752
rect 80756 59712 80762 59724
rect 82998 59712 83004 59724
rect 83056 59712 83062 59764
rect 86218 59712 86224 59764
rect 86276 59752 86282 59764
rect 87414 59752 87420 59764
rect 86276 59724 87420 59752
rect 86276 59712 86282 59724
rect 87414 59712 87420 59724
rect 87472 59712 87478 59764
rect 118602 59712 118608 59764
rect 118660 59752 118666 59764
rect 120258 59752 120264 59764
rect 118660 59724 120264 59752
rect 118660 59712 118666 59724
rect 120258 59712 120264 59724
rect 120316 59712 120322 59764
rect 128998 59712 129004 59764
rect 129056 59752 129062 59764
rect 131574 59752 131580 59764
rect 129056 59724 131580 59752
rect 129056 59712 129062 59724
rect 131574 59712 131580 59724
rect 131632 59712 131638 59764
rect 131758 59712 131764 59764
rect 131816 59752 131822 59764
rect 132586 59752 132592 59764
rect 131816 59724 132592 59752
rect 131816 59712 131822 59724
rect 132586 59712 132592 59724
rect 132644 59712 132650 59764
rect 136542 59712 136548 59764
rect 136600 59752 136606 59764
rect 137830 59752 137836 59764
rect 136600 59724 137836 59752
rect 136600 59712 136606 59724
rect 137830 59712 137836 59724
rect 137888 59712 137894 59764
rect 140038 59712 140044 59764
rect 140096 59752 140102 59764
rect 141970 59752 141976 59764
rect 140096 59724 141976 59752
rect 140096 59712 140102 59724
rect 141970 59712 141976 59724
rect 142028 59712 142034 59764
rect 142798 59712 142804 59764
rect 142856 59752 142862 59764
rect 145006 59752 145012 59764
rect 142856 59724 145012 59752
rect 142856 59712 142862 59724
rect 145006 59712 145012 59724
rect 145064 59712 145070 59764
rect 145742 59712 145748 59764
rect 145800 59752 145806 59764
rect 148134 59752 148140 59764
rect 145800 59724 148140 59752
rect 145800 59712 145806 59724
rect 148134 59712 148140 59724
rect 148192 59712 148198 59764
rect 150342 59712 150348 59764
rect 150400 59752 150406 59764
rect 152274 59752 152280 59764
rect 150400 59724 152280 59752
rect 150400 59712 150406 59724
rect 152274 59712 152280 59724
rect 152332 59712 152338 59764
rect 153838 59712 153844 59764
rect 153896 59752 153902 59764
rect 156598 59752 156604 59764
rect 153896 59724 156604 59752
rect 153896 59712 153902 59724
rect 156598 59712 156604 59724
rect 156656 59712 156662 59764
rect 160738 59712 160744 59764
rect 160796 59752 160802 59764
rect 162578 59752 162584 59764
rect 160796 59724 162584 59752
rect 160796 59712 160802 59724
rect 162578 59712 162584 59724
rect 162636 59712 162642 59764
rect 179230 59712 179236 59764
rect 179288 59752 179294 59764
rect 181254 59752 181260 59764
rect 179288 59724 181260 59752
rect 179288 59712 179294 59724
rect 181254 59712 181260 59724
rect 181312 59712 181318 59764
rect 188890 59712 188896 59764
rect 188948 59752 188954 59764
rect 190546 59752 190552 59764
rect 188948 59724 190552 59752
rect 188948 59712 188954 59724
rect 190546 59712 190552 59724
rect 190604 59712 190610 59764
rect 194502 59712 194508 59764
rect 194560 59752 194566 59764
rect 195790 59752 195796 59764
rect 194560 59724 195796 59752
rect 194560 59712 194566 59724
rect 195790 59712 195796 59724
rect 195848 59712 195854 59764
rect 206922 59712 206928 59764
rect 206980 59752 206986 59764
rect 208118 59752 208124 59764
rect 206980 59724 208124 59752
rect 206980 59712 206986 59724
rect 208118 59712 208124 59724
rect 208176 59712 208182 59764
rect 220446 59712 220452 59764
rect 220504 59752 220510 59764
rect 222562 59752 222568 59764
rect 220504 59724 222568 59752
rect 220504 59712 220510 59724
rect 222562 59712 222568 59724
rect 222620 59712 222626 59764
rect 242802 59712 242808 59764
rect 242860 59752 242866 59764
rect 244274 59752 244280 59764
rect 242860 59724 244280 59752
rect 242860 59712 242866 59724
rect 244274 59712 244280 59724
rect 244332 59712 244338 59764
rect 257890 59712 257896 59764
rect 257948 59752 257954 59764
rect 259822 59752 259828 59764
rect 257948 59724 259828 59752
rect 257948 59712 257954 59724
rect 259822 59712 259828 59724
rect 259880 59712 259886 59764
rect 266262 59712 266268 59764
rect 266320 59752 266326 59764
rect 268102 59752 268108 59764
rect 266320 59724 268108 59752
rect 266320 59712 266326 59724
rect 268102 59712 268108 59724
rect 268160 59712 268166 59764
rect 279418 59712 279424 59764
rect 279476 59752 279482 59764
rect 280614 59752 280620 59764
rect 279476 59724 280620 59752
rect 279476 59712 279482 59724
rect 280614 59712 280620 59724
rect 280672 59712 280678 59764
rect 287698 59712 287704 59764
rect 287756 59752 287762 59764
rect 289814 59752 289820 59764
rect 287756 59724 289820 59752
rect 287756 59712 287762 59724
rect 289814 59712 289820 59724
rect 289872 59712 289878 59764
rect 290642 59712 290648 59764
rect 290700 59752 290706 59764
rect 292942 59752 292948 59764
rect 290700 59724 292948 59752
rect 290700 59712 290706 59724
rect 292942 59712 292948 59724
rect 293000 59712 293006 59764
rect 294598 59712 294604 59764
rect 294656 59752 294662 59764
rect 297082 59752 297088 59764
rect 294656 59724 297088 59752
rect 294656 59712 294662 59724
rect 297082 59712 297088 59724
rect 297140 59712 297146 59764
rect 300118 59712 300124 59764
rect 300176 59752 300182 59764
rect 302234 59752 302240 59764
rect 300176 59724 302240 59752
rect 300176 59712 300182 59724
rect 302234 59712 302240 59724
rect 302292 59712 302298 59764
rect 309042 59712 309048 59764
rect 309100 59752 309106 59764
rect 310514 59752 310520 59764
rect 309100 59724 310520 59752
rect 309100 59712 309106 59724
rect 310514 59712 310520 59724
rect 310572 59712 310578 59764
rect 326706 59712 326712 59764
rect 326764 59752 326770 59764
rect 329282 59752 329288 59764
rect 326764 59724 329288 59752
rect 326764 59712 326770 59724
rect 329282 59712 329288 59724
rect 329340 59712 329346 59764
rect 338022 59712 338028 59764
rect 338080 59752 338086 59764
rect 339494 59752 339500 59764
rect 338080 59724 339500 59752
rect 338080 59712 338086 59724
rect 339494 59712 339500 59724
rect 339552 59712 339558 59764
rect 342162 59712 342168 59764
rect 342220 59752 342226 59764
rect 344278 59752 344284 59764
rect 342220 59724 344284 59752
rect 342220 59712 342226 59724
rect 344278 59712 344284 59724
rect 344336 59712 344342 59764
rect 354674 59712 354680 59764
rect 354732 59752 354738 59764
rect 356698 59752 356704 59764
rect 354732 59724 356704 59752
rect 354732 59712 354738 59724
rect 356698 59712 356704 59724
rect 356756 59712 356762 59764
rect 392854 59712 392860 59764
rect 392912 59752 392918 59764
rect 394878 59752 394884 59764
rect 392912 59724 394884 59752
rect 392912 59712 392918 59724
rect 394878 59712 394884 59724
rect 394936 59712 394942 59764
rect 400122 59712 400128 59764
rect 400180 59752 400186 59764
rect 401594 59752 401600 59764
rect 400180 59724 401600 59752
rect 400180 59712 400186 59724
rect 401594 59712 401600 59724
rect 401652 59712 401658 59764
rect 409506 59712 409512 59764
rect 409564 59752 409570 59764
rect 411622 59752 411628 59764
rect 409564 59724 411628 59752
rect 409564 59712 409570 59724
rect 411622 59712 411628 59724
rect 411680 59712 411686 59764
rect 412634 59712 412640 59764
rect 412692 59752 412698 59764
rect 414106 59752 414112 59764
rect 412692 59724 414112 59752
rect 412692 59712 412698 59724
rect 414106 59712 414112 59724
rect 414164 59712 414170 59764
rect 418706 59712 418712 59764
rect 418764 59752 418770 59764
rect 419810 59752 419816 59764
rect 418764 59724 419816 59752
rect 418764 59712 418770 59724
rect 419810 59712 419816 59724
rect 419868 59712 419874 59764
rect 446674 59712 446680 59764
rect 446732 59752 446738 59764
rect 449342 59752 449348 59764
rect 446732 59724 449348 59752
rect 446732 59712 446738 59724
rect 449342 59712 449348 59724
rect 449400 59712 449406 59764
rect 454954 59712 454960 59764
rect 455012 59752 455018 59764
rect 457622 59752 457628 59764
rect 455012 59724 457628 59752
rect 455012 59712 455018 59724
rect 457622 59712 457628 59724
rect 457680 59712 457686 59764
rect 467282 59712 467288 59764
rect 467340 59752 467346 59764
rect 468478 59752 468484 59764
rect 467340 59724 468484 59752
rect 467340 59712 467346 59724
rect 468478 59712 468484 59724
rect 468536 59712 468542 59764
rect 512822 59712 512828 59764
rect 512880 59752 512886 59764
rect 514846 59752 514852 59764
rect 512880 59724 514852 59752
rect 512880 59712 512886 59724
rect 514846 59712 514852 59724
rect 514904 59712 514910 59764
rect 525242 59712 525248 59764
rect 525300 59752 525306 59764
rect 527358 59752 527364 59764
rect 525300 59724 527364 59752
rect 525300 59712 525306 59724
rect 527358 59712 527364 59724
rect 527416 59712 527422 59764
rect 533706 59712 533712 59764
rect 533764 59752 533770 59764
rect 535638 59752 535644 59764
rect 533764 59724 535644 59752
rect 533764 59712 533770 59724
rect 535638 59712 535644 59724
rect 535696 59712 535702 59764
rect 537662 59712 537668 59764
rect 537720 59752 537726 59764
rect 539778 59752 539784 59764
rect 537720 59724 539784 59752
rect 537720 59712 537726 59724
rect 539778 59712 539784 59724
rect 539836 59712 539842 59764
rect 554314 59712 554320 59764
rect 554372 59752 554378 59764
rect 556338 59752 556344 59764
rect 554372 59724 556344 59752
rect 554372 59712 554378 59724
rect 556338 59712 556344 59724
rect 556396 59712 556402 59764
rect 560386 59712 560392 59764
rect 560444 59752 560450 59764
rect 561766 59752 561772 59764
rect 560444 59724 561772 59752
rect 560444 59712 560450 59724
rect 561766 59712 561772 59724
rect 561824 59712 561830 59764
rect 24854 59576 24860 59628
rect 24912 59616 24918 59628
rect 60550 59616 60556 59628
rect 24912 59588 60556 59616
rect 24912 59576 24918 59588
rect 60550 59576 60556 59588
rect 60608 59576 60614 59628
rect 89162 59576 89168 59628
rect 89220 59616 89226 59628
rect 91278 59616 91284 59628
rect 89220 59588 91284 59616
rect 89220 59576 89226 59588
rect 91278 59576 91284 59588
rect 91336 59576 91342 59628
rect 116578 59576 116584 59628
rect 116636 59616 116642 59628
rect 118142 59616 118148 59628
rect 116636 59588 118148 59616
rect 116636 59576 116642 59588
rect 118142 59576 118148 59588
rect 118200 59576 118206 59628
rect 123478 59576 123484 59628
rect 123536 59616 123542 59628
rect 125410 59616 125416 59628
rect 123536 59588 125416 59616
rect 123536 59576 123542 59588
rect 125410 59576 125416 59588
rect 125468 59576 125474 59628
rect 284938 59576 284944 59628
rect 284996 59616 285002 59628
rect 286686 59616 286692 59628
rect 284996 59588 286692 59616
rect 284996 59576 285002 59588
rect 286686 59576 286692 59588
rect 286744 59576 286750 59628
rect 322198 59576 322204 59628
rect 322256 59616 322262 59628
rect 325142 59616 325148 59628
rect 322256 59588 325148 59616
rect 322256 59576 322262 59588
rect 325142 59576 325148 59588
rect 325200 59576 325206 59628
rect 328730 59576 328736 59628
rect 328788 59616 328794 59628
rect 330478 59616 330484 59628
rect 328788 59588 330484 59616
rect 328788 59576 328794 59588
rect 330478 59576 330484 59588
rect 330536 59576 330542 59628
rect 345290 59576 345296 59628
rect 345348 59616 345354 59628
rect 347038 59616 347044 59628
rect 345348 59588 347044 59616
rect 345348 59576 345354 59588
rect 347038 59576 347044 59588
rect 347096 59576 347102 59628
rect 461118 59576 461124 59628
rect 461176 59616 461182 59628
rect 462958 59616 462964 59628
rect 461176 59588 462964 59616
rect 461176 59576 461182 59588
rect 462958 59576 462964 59588
rect 463016 59576 463022 59628
rect 541802 59576 541808 59628
rect 541860 59616 541866 59628
rect 544010 59616 544016 59628
rect 541860 59588 544016 59616
rect 541860 59576 541866 59588
rect 544010 59576 544016 59588
rect 544068 59576 544074 59628
rect 561490 59576 561496 59628
rect 561548 59616 561554 59628
rect 563054 59616 563060 59628
rect 561548 59588 563060 59616
rect 561548 59576 561554 59588
rect 563054 59576 563060 59588
rect 563112 59576 563118 59628
rect 19334 59508 19340 59560
rect 19392 59548 19398 59560
rect 62298 59548 62304 59560
rect 19392 59520 62304 59548
rect 19392 59508 19398 59520
rect 62298 59508 62304 59520
rect 62356 59508 62362 59560
rect 5534 59440 5540 59492
rect 5592 59480 5598 59492
rect 57790 59480 57796 59492
rect 5592 59452 57796 59480
rect 5592 59440 5598 59452
rect 57790 59440 57796 59452
rect 57848 59440 57854 59492
rect 114002 59440 114008 59492
rect 114060 59480 114066 59492
rect 116118 59480 116124 59492
rect 114060 59452 116124 59480
rect 114060 59440 114066 59452
rect 116118 59440 116124 59452
rect 116176 59440 116182 59492
rect 175090 59440 175096 59492
rect 175148 59480 175154 59492
rect 177114 59480 177120 59492
rect 175148 59452 177120 59480
rect 175148 59440 175154 59452
rect 177114 59440 177120 59452
rect 177172 59440 177178 59492
rect 191742 59440 191748 59492
rect 191800 59480 191806 59492
rect 193674 59480 193680 59492
rect 191800 59452 193680 59480
rect 191800 59440 191806 59452
rect 193674 59440 193680 59452
rect 193732 59440 193738 59492
rect 203886 59440 203892 59492
rect 203944 59480 203950 59492
rect 206094 59480 206100 59492
rect 203944 59452 206100 59480
rect 203944 59440 203950 59452
rect 206094 59440 206100 59452
rect 206152 59440 206158 59492
rect 224862 59440 224868 59492
rect 224920 59480 224926 59492
rect 226702 59480 226708 59492
rect 224920 59452 226708 59480
rect 224920 59440 224926 59452
rect 226702 59440 226708 59452
rect 226760 59440 226766 59492
rect 233050 59440 233056 59492
rect 233108 59480 233114 59492
rect 234982 59480 234988 59492
rect 233108 59452 234988 59480
rect 233108 59440 233114 59452
rect 234982 59440 234988 59452
rect 235040 59440 235046 59492
rect 249702 59440 249708 59492
rect 249760 59480 249766 59492
rect 251542 59480 251548 59492
rect 249760 59452 251548 59480
rect 249760 59440 249766 59452
rect 251542 59440 251548 59452
rect 251600 59440 251606 59492
rect 253750 59440 253756 59492
rect 253808 59480 253814 59492
rect 255682 59480 255688 59492
rect 253808 59452 255688 59480
rect 253808 59440 253814 59452
rect 255682 59440 255688 59452
rect 255740 59440 255746 59492
rect 256602 59440 256608 59492
rect 256660 59480 256666 59492
rect 257798 59480 257804 59492
rect 256660 59452 257804 59480
rect 256660 59440 256666 59452
rect 257798 59440 257804 59452
rect 257856 59440 257862 59492
rect 282178 59440 282184 59492
rect 282236 59480 282242 59492
rect 284662 59480 284668 59492
rect 282236 59452 284668 59480
rect 282236 59440 282242 59452
rect 284662 59440 284668 59452
rect 284720 59440 284726 59492
rect 405274 59440 405280 59492
rect 405332 59480 405338 59492
rect 407298 59480 407304 59492
rect 405332 59452 407304 59480
rect 405332 59440 405338 59452
rect 407298 59440 407304 59452
rect 407356 59440 407362 59492
rect 420822 59440 420828 59492
rect 420880 59480 420886 59492
rect 422386 59480 422392 59492
rect 420880 59452 422392 59480
rect 420880 59440 420886 59452
rect 422386 59440 422392 59452
rect 422444 59440 422450 59492
rect 443546 59440 443552 59492
rect 443604 59480 443610 59492
rect 444374 59480 444380 59492
rect 443604 59452 444380 59480
rect 443604 59440 443610 59452
rect 444374 59440 444380 59452
rect 444432 59440 444438 59492
rect 492122 59440 492128 59492
rect 492180 59480 492186 59492
rect 494238 59480 494244 59492
rect 492180 59452 494244 59480
rect 492180 59440 492186 59452
rect 494238 59440 494244 59452
rect 494296 59440 494302 59492
rect 504542 59440 504548 59492
rect 504600 59480 504606 59492
rect 506658 59480 506664 59492
rect 504600 59452 506664 59480
rect 504600 59440 504606 59452
rect 506658 59440 506664 59452
rect 506716 59440 506722 59492
rect 4154 59372 4160 59424
rect 4212 59412 4218 59424
rect 58158 59412 58164 59424
rect 4212 59384 58164 59412
rect 4212 59372 4218 59384
rect 58158 59372 58164 59384
rect 58216 59372 58222 59424
rect 365806 59372 365812 59424
rect 365864 59412 365870 59424
rect 366542 59412 366548 59424
rect 365864 59384 366548 59412
rect 365864 59372 365870 59384
rect 366542 59372 366548 59384
rect 366600 59372 366606 59424
rect 384482 59372 384488 59424
rect 384540 59412 384546 59424
rect 385218 59412 385224 59424
rect 384540 59384 385224 59412
rect 384540 59372 384546 59384
rect 385218 59372 385224 59384
rect 385276 59372 385282 59424
rect 101950 59304 101956 59356
rect 102008 59344 102014 59356
rect 103422 59344 103428 59356
rect 102008 59316 103428 59344
rect 102008 59304 102014 59316
rect 103422 59304 103428 59316
rect 103480 59304 103486 59356
rect 262214 59304 262220 59356
rect 262272 59344 262278 59356
rect 263962 59344 263968 59356
rect 262272 59316 263968 59344
rect 262272 59304 262278 59316
rect 263962 59304 263968 59316
rect 264020 59304 264026 59356
rect 362218 59032 362224 59084
rect 362276 59072 362282 59084
rect 389174 59072 389180 59084
rect 362276 59044 389180 59072
rect 362276 59032 362282 59044
rect 389174 59032 389180 59044
rect 389232 59032 389238 59084
rect 328454 58964 328460 59016
rect 328512 59004 328518 59016
rect 376754 59004 376760 59016
rect 328512 58976 376760 59004
rect 328512 58964 328518 58976
rect 376754 58964 376760 58976
rect 376812 58964 376818 59016
rect 217962 58896 217968 58948
rect 218020 58936 218026 58948
rect 425054 58936 425060 58948
rect 218020 58908 425060 58936
rect 218020 58896 218026 58908
rect 425054 58896 425060 58908
rect 425112 58896 425118 58948
rect 449710 58896 449716 58948
rect 449768 58936 449774 58948
rect 536834 58936 536840 58948
rect 449768 58908 536840 58936
rect 449768 58896 449774 58908
rect 536834 58896 536840 58908
rect 536892 58896 536898 58948
rect 306190 58828 306196 58880
rect 306248 58868 306254 58880
rect 572714 58868 572720 58880
rect 306248 58840 572720 58868
rect 306248 58828 306254 58840
rect 572714 58828 572720 58840
rect 572772 58828 572778 58880
rect 259454 58760 259460 58812
rect 259512 58800 259518 58812
rect 529014 58800 529020 58812
rect 259512 58772 529020 58800
rect 259512 58760 259518 58772
rect 529014 58760 529020 58772
rect 529072 58760 529078 58812
rect 53834 58692 53840 58744
rect 53892 58732 53898 58744
rect 150342 58732 150348 58744
rect 53892 58704 150348 58732
rect 53892 58692 53898 58704
rect 150342 58692 150348 58704
rect 150400 58692 150406 58744
rect 188982 58692 188988 58744
rect 189040 58732 189046 58744
rect 524414 58732 524420 58744
rect 189040 58704 524420 58732
rect 189040 58692 189046 58704
rect 524414 58692 524420 58704
rect 524472 58692 524478 58744
rect 49694 58624 49700 58676
rect 49752 58664 49758 58676
rect 85482 58664 85488 58676
rect 49752 58636 85488 58664
rect 49752 58624 49758 58636
rect 85482 58624 85488 58636
rect 85540 58624 85546 58676
rect 109862 58624 109868 58676
rect 109920 58664 109926 58676
rect 110874 58664 110880 58676
rect 109920 58636 110880 58664
rect 109920 58624 109926 58636
rect 110874 58624 110880 58636
rect 110932 58624 110938 58676
rect 146294 58624 146300 58676
rect 146352 58664 146358 58676
rect 561858 58664 561864 58676
rect 146352 58636 561864 58664
rect 146352 58624 146358 58636
rect 561858 58624 561864 58636
rect 561916 58624 561922 58676
rect 246942 58556 246948 58608
rect 247000 58596 247006 58608
rect 248414 58596 248420 58608
rect 247000 58568 248420 58596
rect 247000 58556 247006 58568
rect 248414 58556 248420 58568
rect 248472 58556 248478 58608
rect 322106 58488 322112 58540
rect 322164 58528 322170 58540
rect 323578 58528 323584 58540
rect 322164 58500 323584 58528
rect 322164 58488 322170 58500
rect 323578 58488 323584 58500
rect 323636 58488 323642 58540
rect 245286 58352 245292 58404
rect 245344 58392 245350 58404
rect 246758 58392 246764 58404
rect 245344 58364 246764 58392
rect 245344 58352 245350 58364
rect 246758 58352 246764 58364
rect 246816 58352 246822 58404
rect 320450 58352 320456 58404
rect 320508 58392 320514 58404
rect 322198 58392 322204 58404
rect 320508 58364 322204 58392
rect 320508 58352 320514 58364
rect 322198 58352 322204 58364
rect 322256 58352 322262 58404
rect 384114 58352 384120 58404
rect 384172 58392 384178 58404
rect 385034 58392 385040 58404
rect 384172 58364 385040 58392
rect 384172 58352 384178 58364
rect 385034 58352 385040 58364
rect 385092 58352 385098 58404
rect 342254 57536 342260 57588
rect 342312 57576 342318 57588
rect 373994 57576 374000 57588
rect 342312 57548 374000 57576
rect 342312 57536 342318 57548
rect 373994 57536 374000 57548
rect 374052 57536 374058 57588
rect 242710 57468 242716 57520
rect 242768 57508 242774 57520
rect 340874 57508 340880 57520
rect 242768 57480 340880 57508
rect 242768 57468 242774 57480
rect 340874 57468 340880 57480
rect 340932 57468 340938 57520
rect 374086 57468 374092 57520
rect 374144 57508 374150 57520
rect 495618 57508 495624 57520
rect 374144 57480 495624 57508
rect 374144 57468 374150 57480
rect 495618 57468 495624 57480
rect 495676 57468 495682 57520
rect 251174 57400 251180 57452
rect 251232 57440 251238 57452
rect 266078 57440 266084 57452
rect 251232 57412 266084 57440
rect 251232 57400 251238 57412
rect 266078 57400 266084 57412
rect 266136 57400 266142 57452
rect 339494 57400 339500 57452
rect 339552 57440 339558 57452
rect 466454 57440 466460 57452
rect 339552 57412 466460 57440
rect 339552 57400 339558 57412
rect 466454 57400 466460 57412
rect 466512 57400 466518 57452
rect 204254 57332 204260 57384
rect 204312 57372 204318 57384
rect 413186 57372 413192 57384
rect 204312 57344 413192 57372
rect 204312 57332 204318 57344
rect 413186 57332 413192 57344
rect 413244 57332 413250 57384
rect 161474 57264 161480 57316
rect 161532 57304 161538 57316
rect 425330 57304 425336 57316
rect 161532 57276 425336 57304
rect 161532 57264 161538 57276
rect 425330 57264 425336 57276
rect 425388 57264 425394 57316
rect 444558 57264 444564 57316
rect 444616 57304 444622 57316
rect 557534 57304 557540 57316
rect 444616 57276 557540 57304
rect 444616 57264 444622 57276
rect 557534 57264 557540 57276
rect 557592 57264 557598 57316
rect 7558 57196 7564 57248
rect 7616 57236 7622 57248
rect 164142 57236 164148 57248
rect 7616 57208 164148 57236
rect 7616 57196 7622 57208
rect 164142 57196 164148 57208
rect 164200 57196 164206 57248
rect 263594 57196 263600 57248
rect 263652 57236 263658 57248
rect 528646 57236 528652 57248
rect 263652 57208 528652 57236
rect 263652 57196 263658 57208
rect 528646 57196 528652 57208
rect 528704 57196 528710 57248
rect 353294 56176 353300 56228
rect 353352 56216 353358 56228
rect 420914 56216 420920 56228
rect 353352 56188 420920 56216
rect 353352 56176 353358 56188
rect 420914 56176 420920 56188
rect 420972 56176 420978 56228
rect 430574 56176 430580 56228
rect 430632 56216 430638 56228
rect 481634 56216 481640 56228
rect 430632 56188 481640 56216
rect 430632 56176 430638 56188
rect 481634 56176 481640 56188
rect 481692 56176 481698 56228
rect 267734 56108 267740 56160
rect 267792 56148 267798 56160
rect 394694 56148 394700 56160
rect 267792 56120 394700 56148
rect 267792 56108 267798 56120
rect 394694 56108 394700 56120
rect 394752 56108 394758 56160
rect 248414 56040 248420 56092
rect 248472 56080 248478 56092
rect 266262 56080 266268 56092
rect 248472 56052 266268 56080
rect 248472 56040 248478 56052
rect 266262 56040 266268 56052
rect 266320 56040 266326 56092
rect 335354 56040 335360 56092
rect 335412 56080 335418 56092
rect 481634 56080 481640 56092
rect 335412 56052 481640 56080
rect 335412 56040 335418 56052
rect 481634 56040 481640 56052
rect 481692 56040 481698 56092
rect 229002 55972 229008 56024
rect 229060 56012 229066 56024
rect 379514 56012 379520 56024
rect 229060 55984 379520 56012
rect 229060 55972 229066 55984
rect 379514 55972 379520 55984
rect 379572 55972 379578 56024
rect 103514 55904 103520 55956
rect 103572 55944 103578 55956
rect 136542 55944 136548 55956
rect 103572 55916 136548 55944
rect 103572 55904 103578 55916
rect 136542 55904 136548 55916
rect 136600 55904 136606 55956
rect 168374 55904 168380 55956
rect 168432 55944 168438 55956
rect 423674 55944 423680 55956
rect 168432 55916 423680 55944
rect 168432 55904 168438 55916
rect 423674 55904 423680 55916
rect 423732 55904 423738 55956
rect 444374 55904 444380 55956
rect 444432 55944 444438 55956
rect 561674 55944 561680 55956
rect 444432 55916 561680 55944
rect 444432 55904 444438 55916
rect 561674 55904 561680 55916
rect 561732 55904 561738 55956
rect 48314 55836 48320 55888
rect 48372 55876 48378 55888
rect 118602 55876 118608 55888
rect 48372 55848 118608 55876
rect 48372 55836 48378 55848
rect 118602 55836 118608 55848
rect 118660 55836 118666 55888
rect 135254 55836 135260 55888
rect 135312 55876 135318 55888
rect 567286 55876 567292 55888
rect 135312 55848 567292 55876
rect 135312 55836 135318 55848
rect 567286 55836 567292 55848
rect 567344 55836 567350 55888
rect 261938 54952 261944 55004
rect 261996 54992 262002 55004
rect 266354 54992 266360 55004
rect 261996 54964 266360 54992
rect 261996 54952 262002 54964
rect 266354 54952 266360 54964
rect 266412 54952 266418 55004
rect 303614 54816 303620 54868
rect 303672 54856 303678 54868
rect 386414 54856 386420 54868
rect 303672 54828 386420 54856
rect 303672 54816 303678 54828
rect 386414 54816 386420 54828
rect 386472 54816 386478 54868
rect 233050 54748 233056 54800
rect 233108 54788 233114 54800
rect 361574 54788 361580 54800
rect 233108 54760 361580 54788
rect 233108 54748 233114 54760
rect 361574 54748 361580 54760
rect 361632 54748 361638 54800
rect 362126 54748 362132 54800
rect 362184 54788 362190 54800
rect 391934 54788 391940 54800
rect 362184 54760 391940 54788
rect 362184 54748 362190 54760
rect 391934 54748 391940 54760
rect 391992 54748 391998 54800
rect 216490 54680 216496 54732
rect 216548 54720 216554 54732
rect 418154 54720 418160 54732
rect 216548 54692 418160 54720
rect 216548 54680 216554 54692
rect 418154 54680 418160 54692
rect 418212 54680 418218 54732
rect 458174 54680 458180 54732
rect 458232 54720 458238 54732
rect 473354 54720 473360 54732
rect 458232 54692 473360 54720
rect 458232 54680 458238 54692
rect 473354 54680 473360 54692
rect 473412 54680 473418 54732
rect 162854 54612 162860 54664
rect 162912 54652 162918 54664
rect 290642 54652 290648 54664
rect 162912 54624 290648 54652
rect 162912 54612 162918 54624
rect 290642 54612 290648 54624
rect 290700 54612 290706 54664
rect 309042 54612 309048 54664
rect 309100 54652 309106 54664
rect 556154 54652 556160 54664
rect 309100 54624 556160 54652
rect 309100 54612 309106 54624
rect 556154 54612 556160 54624
rect 556212 54612 556218 54664
rect 274634 54544 274640 54596
rect 274692 54584 274698 54596
rect 527174 54584 527180 54596
rect 274692 54556 527180 54584
rect 274692 54544 274698 54556
rect 527174 54544 527180 54556
rect 527232 54544 527238 54596
rect 10318 54476 10324 54528
rect 10376 54516 10382 54528
rect 162578 54516 162584 54528
rect 10376 54488 162584 54516
rect 10376 54476 10382 54488
rect 162578 54476 162584 54488
rect 162636 54476 162642 54528
rect 168466 54476 168472 54528
rect 168524 54516 168530 54528
rect 556614 54516 556620 54528
rect 168524 54488 556620 54516
rect 168524 54476 168530 54488
rect 556614 54476 556620 54488
rect 556672 54476 556678 54528
rect 311618 53320 311624 53372
rect 311676 53360 311682 53372
rect 545206 53360 545212 53372
rect 311676 53332 545212 53360
rect 311676 53320 311682 53332
rect 545206 53320 545212 53332
rect 545264 53320 545270 53372
rect 288434 53252 288440 53304
rect 288492 53292 288498 53304
rect 523034 53292 523040 53304
rect 288492 53264 523040 53292
rect 288492 53252 288498 53264
rect 523034 53252 523040 53264
rect 523092 53252 523098 53304
rect 140774 53184 140780 53236
rect 140832 53224 140838 53236
rect 434714 53224 434720 53236
rect 140832 53196 434720 53224
rect 140832 53184 140838 53196
rect 434714 53184 434720 53196
rect 434772 53184 434778 53236
rect 469214 53184 469220 53236
rect 469272 53224 469278 53236
rect 476114 53224 476120 53236
rect 469272 53196 476120 53224
rect 469272 53184 469278 53196
rect 476114 53184 476120 53196
rect 476172 53184 476178 53236
rect 183462 53116 183468 53168
rect 183520 53156 183526 53168
rect 530578 53156 530584 53168
rect 183520 53128 530584 53156
rect 183520 53116 183526 53128
rect 530578 53116 530584 53128
rect 530636 53116 530642 53168
rect 57974 53048 57980 53100
rect 58032 53088 58038 53100
rect 149698 53088 149704 53100
rect 58032 53060 149704 53088
rect 58032 53048 58038 53060
rect 149698 53048 149704 53060
rect 149756 53048 149762 53100
rect 200114 53048 200120 53100
rect 200172 53088 200178 53100
rect 549254 53088 549260 53100
rect 200172 53060 549260 53088
rect 200172 53048 200178 53060
rect 549254 53048 549260 53060
rect 549312 53048 549318 53100
rect 332594 51960 332600 52012
rect 332652 52000 332658 52012
rect 488534 52000 488540 52012
rect 332652 51972 488540 52000
rect 332652 51960 332658 51972
rect 488534 51960 488540 51972
rect 488592 51960 488598 52012
rect 313274 51892 313280 51944
rect 313332 51932 313338 51944
rect 516134 51932 516140 51944
rect 313332 51904 516140 51932
rect 313332 51892 313338 51904
rect 516134 51892 516140 51904
rect 516192 51892 516198 51944
rect 133874 51824 133880 51876
rect 133932 51864 133938 51876
rect 436186 51864 436192 51876
rect 133932 51836 436192 51864
rect 133932 51824 133938 51836
rect 436186 51824 436192 51836
rect 436244 51824 436250 51876
rect 188890 51756 188896 51808
rect 188948 51796 188954 51808
rect 514754 51796 514760 51808
rect 188948 51768 514760 51796
rect 188948 51756 188954 51768
rect 514754 51756 514760 51768
rect 514812 51756 514818 51808
rect 44174 51688 44180 51740
rect 44232 51728 44238 51740
rect 154022 51728 154028 51740
rect 44232 51700 154028 51728
rect 44232 51688 44238 51700
rect 154022 51688 154028 51700
rect 154080 51688 154086 51740
rect 213914 51688 213920 51740
rect 213972 51728 213978 51740
rect 545114 51728 545120 51740
rect 213972 51700 545120 51728
rect 213972 51688 213978 51700
rect 545114 51688 545120 51700
rect 545172 51688 545178 51740
rect 355318 50668 355324 50720
rect 355376 50708 355382 50720
rect 414014 50708 414020 50720
rect 355376 50680 414020 50708
rect 355376 50668 355382 50680
rect 414014 50668 414020 50680
rect 414072 50668 414078 50720
rect 292574 50600 292580 50652
rect 292632 50640 292638 50652
rect 390646 50640 390652 50652
rect 292632 50612 390652 50640
rect 292632 50600 292638 50612
rect 390646 50600 390652 50612
rect 390704 50600 390710 50652
rect 321002 50532 321008 50584
rect 321060 50572 321066 50584
rect 531406 50572 531412 50584
rect 321060 50544 531412 50572
rect 321060 50532 321066 50544
rect 531406 50532 531412 50544
rect 531464 50532 531470 50584
rect 218054 50464 218060 50516
rect 218112 50504 218118 50516
rect 543826 50504 543832 50516
rect 218112 50476 543832 50504
rect 218112 50464 218118 50476
rect 543826 50464 543832 50476
rect 543884 50464 543890 50516
rect 40034 50396 40040 50448
rect 40092 50436 40098 50448
rect 153838 50436 153844 50448
rect 40092 50408 153844 50436
rect 40092 50396 40098 50408
rect 153838 50396 153844 50408
rect 153896 50396 153902 50448
rect 179230 50396 179236 50448
rect 179288 50436 179294 50448
rect 546586 50436 546592 50448
rect 179288 50408 546592 50436
rect 179288 50396 179294 50408
rect 546586 50396 546592 50408
rect 546644 50396 546650 50448
rect 139394 50328 139400 50380
rect 139452 50368 139458 50380
rect 567194 50368 567200 50380
rect 139452 50340 567200 50368
rect 139452 50328 139458 50340
rect 567194 50328 567200 50340
rect 567252 50328 567258 50380
rect 258074 49240 258080 49292
rect 258132 49280 258138 49292
rect 400214 49280 400220 49292
rect 258132 49252 400220 49280
rect 258132 49240 258138 49252
rect 400214 49240 400220 49252
rect 400272 49240 400278 49292
rect 325142 49172 325148 49224
rect 325200 49212 325206 49224
rect 520274 49212 520280 49224
rect 325200 49184 520280 49212
rect 325200 49172 325206 49184
rect 520274 49172 520280 49184
rect 520332 49172 520338 49224
rect 151814 49104 151820 49156
rect 151872 49144 151878 49156
rect 294782 49144 294788 49156
rect 151872 49116 294788 49144
rect 151872 49104 151878 49116
rect 294782 49104 294788 49116
rect 294840 49104 294846 49156
rect 316034 49104 316040 49156
rect 316092 49144 316098 49156
rect 515030 49144 515036 49156
rect 316092 49116 515036 49144
rect 316092 49104 316098 49116
rect 515030 49104 515036 49116
rect 515088 49104 515094 49156
rect 110506 49036 110512 49088
rect 110564 49076 110570 49088
rect 133322 49076 133328 49088
rect 110564 49048 133328 49076
rect 110564 49036 110570 49048
rect 133322 49036 133328 49048
rect 133380 49036 133386 49088
rect 143534 49036 143540 49088
rect 143592 49076 143598 49088
rect 433334 49076 433340 49088
rect 143592 49048 433340 49076
rect 143592 49036 143598 49048
rect 433334 49036 433340 49048
rect 433392 49036 433398 49088
rect 52454 48968 52460 49020
rect 52512 49008 52518 49020
rect 117958 49008 117964 49020
rect 52512 48980 117964 49008
rect 52512 48968 52518 48980
rect 117958 48968 117964 48980
rect 118016 48968 118022 49020
rect 209774 48968 209780 49020
rect 209832 49008 209838 49020
rect 546494 49008 546500 49020
rect 209832 48980 546500 49008
rect 209832 48968 209838 48980
rect 546494 48968 546500 48980
rect 546552 48968 546558 49020
rect 276014 47880 276020 47932
rect 276072 47920 276078 47932
rect 394786 47920 394792 47932
rect 276072 47892 394792 47920
rect 276072 47880 276078 47892
rect 394786 47880 394792 47892
rect 394844 47880 394850 47932
rect 341702 47812 341708 47864
rect 341760 47852 341766 47864
rect 463694 47852 463700 47864
rect 341760 47824 463700 47852
rect 341760 47812 341766 47824
rect 463694 47812 463700 47824
rect 463752 47812 463758 47864
rect 219342 47744 219348 47796
rect 219400 47784 219406 47796
rect 411254 47784 411260 47796
rect 219400 47756 411260 47784
rect 219400 47744 219406 47756
rect 411254 47744 411260 47756
rect 411312 47744 411318 47796
rect 201494 47676 201500 47728
rect 201552 47716 201558 47728
rect 279418 47716 279424 47728
rect 201552 47688 279424 47716
rect 201552 47676 201558 47688
rect 279418 47676 279424 47688
rect 279476 47676 279482 47728
rect 323578 47676 323584 47728
rect 323636 47716 323642 47728
rect 523034 47716 523040 47728
rect 323636 47688 523040 47716
rect 323636 47676 323642 47688
rect 523034 47676 523040 47688
rect 523092 47676 523098 47728
rect 93854 47608 93860 47660
rect 93912 47648 93918 47660
rect 138658 47648 138664 47660
rect 93912 47620 138664 47648
rect 93912 47608 93918 47620
rect 138658 47608 138664 47620
rect 138716 47608 138722 47660
rect 207014 47608 207020 47660
rect 207072 47648 207078 47660
rect 547874 47648 547880 47660
rect 207072 47620 547880 47648
rect 207072 47608 207078 47620
rect 547874 47608 547880 47620
rect 547932 47608 547938 47660
rect 11698 47540 11704 47592
rect 11756 47580 11762 47592
rect 95878 47580 95884 47592
rect 11756 47552 95884 47580
rect 11756 47540 11762 47552
rect 95878 47540 95884 47552
rect 95936 47540 95942 47592
rect 143626 47540 143632 47592
rect 143684 47580 143690 47592
rect 565814 47580 565820 47592
rect 143684 47552 565820 47580
rect 143684 47540 143690 47552
rect 565814 47540 565820 47552
rect 565872 47540 565878 47592
rect 364334 47064 364340 47116
rect 364392 47104 364398 47116
rect 369946 47104 369952 47116
rect 364392 47076 369952 47104
rect 364392 47064 364398 47076
rect 369946 47064 369952 47076
rect 370004 47064 370010 47116
rect 338114 46520 338120 46572
rect 338172 46560 338178 46572
rect 509234 46560 509240 46572
rect 338172 46532 509240 46560
rect 338172 46520 338178 46532
rect 509234 46520 509240 46532
rect 509292 46520 509298 46572
rect 222102 46452 222108 46504
rect 222160 46492 222166 46504
rect 400214 46492 400220 46504
rect 222160 46464 400220 46492
rect 222160 46452 222166 46464
rect 400214 46452 400220 46464
rect 400272 46452 400278 46504
rect 325694 46384 325700 46436
rect 325752 46424 325758 46436
rect 513374 46424 513380 46436
rect 325752 46396 513380 46424
rect 325752 46384 325758 46396
rect 513374 46384 513380 46396
rect 513432 46384 513438 46436
rect 208394 46316 208400 46368
rect 208452 46356 208458 46368
rect 415578 46356 415584 46368
rect 208452 46328 415584 46356
rect 208452 46316 208458 46328
rect 415578 46316 415584 46328
rect 415636 46316 415642 46368
rect 469858 46316 469864 46368
rect 469916 46356 469922 46368
rect 473354 46356 473360 46368
rect 469916 46328 473360 46356
rect 469916 46316 469922 46328
rect 473354 46316 473360 46328
rect 473412 46316 473418 46368
rect 198642 46248 198648 46300
rect 198700 46288 198706 46300
rect 481726 46288 481732 46300
rect 198700 46260 481732 46288
rect 198700 46248 198706 46260
rect 481726 46248 481732 46260
rect 481784 46248 481790 46300
rect 3418 46180 3424 46232
rect 3476 46220 3482 46232
rect 164878 46220 164884 46232
rect 3476 46192 164884 46220
rect 3476 46180 3482 46192
rect 164878 46180 164884 46192
rect 164936 46180 164942 46232
rect 195974 46180 195980 46232
rect 196032 46220 196038 46232
rect 550634 46220 550640 46232
rect 196032 46192 550640 46220
rect 196032 46180 196038 46192
rect 550634 46180 550640 46192
rect 550692 46180 550698 46232
rect 337562 45160 337568 45212
rect 337620 45200 337626 45212
rect 473446 45200 473452 45212
rect 337620 45172 473452 45200
rect 337620 45160 337626 45172
rect 473446 45160 473452 45172
rect 473504 45160 473510 45212
rect 244182 45092 244188 45144
rect 244240 45132 244246 45144
rect 325694 45132 325700 45144
rect 244240 45104 325700 45132
rect 244240 45092 244246 45104
rect 325694 45092 325700 45104
rect 325752 45092 325758 45144
rect 334618 45092 334624 45144
rect 334676 45132 334682 45144
rect 484394 45132 484400 45144
rect 334676 45104 484400 45132
rect 334676 45092 334682 45104
rect 484394 45092 484400 45104
rect 484452 45092 484458 45144
rect 138014 45024 138020 45076
rect 138072 45064 138078 45076
rect 298922 45064 298928 45076
rect 138072 45036 298928 45064
rect 138072 45024 138078 45036
rect 298922 45024 298928 45036
rect 298980 45024 298986 45076
rect 349154 45024 349160 45076
rect 349212 45064 349218 45076
rect 506658 45064 506664 45076
rect 349212 45036 506664 45064
rect 349212 45024 349218 45036
rect 506658 45024 506664 45036
rect 506716 45024 506722 45076
rect 193214 44956 193220 45008
rect 193272 44996 193278 45008
rect 419626 44996 419632 45008
rect 193272 44968 419632 44996
rect 193272 44956 193278 44968
rect 419626 44956 419632 44968
rect 419684 44956 419690 45008
rect 211062 44888 211068 44940
rect 211120 44928 211126 44940
rect 440234 44928 440240 44940
rect 211120 44900 440240 44928
rect 211120 44888 211126 44900
rect 440234 44888 440240 44900
rect 440292 44888 440298 44940
rect 62114 44820 62120 44872
rect 62172 44860 62178 44872
rect 114002 44860 114008 44872
rect 62172 44832 114008 44860
rect 62172 44820 62178 44832
rect 114002 44820 114008 44832
rect 114060 44820 114066 44872
rect 128354 44820 128360 44872
rect 128412 44860 128418 44872
rect 569954 44860 569960 44872
rect 128412 44832 569960 44860
rect 128412 44820 128418 44832
rect 569954 44820 569960 44832
rect 570012 44820 570018 44872
rect 338758 43732 338764 43784
rect 338816 43772 338822 43784
rect 470594 43772 470600 43784
rect 338816 43744 470600 43772
rect 338816 43732 338822 43744
rect 470594 43732 470600 43744
rect 470652 43732 470658 43784
rect 233234 43664 233240 43716
rect 233292 43704 233298 43716
rect 407114 43704 407120 43716
rect 233292 43676 407120 43704
rect 233292 43664 233298 43676
rect 407114 43664 407120 43676
rect 407172 43664 407178 43716
rect 331214 43596 331220 43648
rect 331272 43636 331278 43648
rect 510706 43636 510712 43648
rect 331272 43608 510712 43636
rect 331272 43596 331278 43608
rect 510706 43596 510712 43608
rect 510764 43596 510770 43648
rect 324958 43528 324964 43580
rect 325016 43568 325022 43580
rect 516134 43568 516140 43580
rect 325016 43540 516140 43568
rect 325016 43528 325022 43540
rect 516134 43528 516140 43540
rect 516192 43528 516198 43580
rect 193306 43460 193312 43512
rect 193364 43500 193370 43512
rect 552106 43500 552112 43512
rect 193364 43472 552112 43500
rect 193364 43460 193370 43472
rect 552106 43460 552112 43472
rect 552164 43460 552170 43512
rect 46934 43392 46940 43444
rect 46992 43432 46998 43444
rect 152458 43432 152464 43444
rect 46992 43404 152464 43432
rect 46992 43392 46998 43404
rect 152458 43392 152464 43404
rect 152516 43392 152522 43444
rect 173802 43392 173808 43444
rect 173860 43432 173866 43444
rect 566458 43432 566464 43444
rect 173860 43404 566464 43432
rect 173860 43392 173866 43404
rect 566458 43392 566464 43404
rect 566516 43392 566522 43444
rect 226242 42372 226248 42424
rect 226300 42412 226306 42424
rect 386414 42412 386420 42424
rect 226300 42384 386420 42412
rect 226300 42372 226306 42384
rect 386414 42372 386420 42384
rect 386472 42372 386478 42424
rect 345014 42304 345020 42356
rect 345072 42344 345078 42356
rect 506474 42344 506480 42356
rect 345072 42316 506480 42344
rect 345072 42304 345078 42316
rect 506474 42304 506480 42316
rect 506532 42304 506538 42356
rect 331858 42236 331864 42288
rect 331916 42276 331922 42288
rect 495434 42276 495440 42288
rect 331916 42248 495440 42276
rect 331916 42236 331922 42248
rect 495434 42236 495440 42248
rect 495492 42236 495498 42288
rect 197262 42168 197268 42220
rect 197320 42208 197326 42220
rect 485774 42208 485780 42220
rect 197320 42180 485780 42208
rect 197320 42168 197326 42180
rect 485774 42168 485780 42180
rect 485832 42168 485838 42220
rect 129734 42100 129740 42152
rect 129792 42140 129798 42152
rect 437474 42140 437480 42152
rect 129792 42112 437480 42140
rect 129792 42100 129798 42112
rect 437474 42100 437480 42112
rect 437532 42100 437538 42152
rect 80054 42032 80060 42084
rect 80112 42072 80118 42084
rect 109862 42072 109868 42084
rect 80112 42044 109868 42072
rect 80112 42032 80118 42044
rect 109862 42032 109868 42044
rect 109920 42032 109926 42084
rect 189074 42032 189080 42084
rect 189132 42072 189138 42084
rect 552290 42072 552296 42084
rect 189132 42044 552296 42072
rect 189132 42032 189138 42044
rect 552290 42032 552296 42044
rect 552348 42032 552354 42084
rect 241330 40944 241336 40996
rect 241388 40984 241394 40996
rect 336734 40984 336740 40996
rect 241388 40956 336740 40984
rect 241388 40944 241394 40956
rect 336734 40944 336740 40956
rect 336792 40944 336798 40996
rect 337378 40944 337384 40996
rect 337436 40984 337442 40996
rect 477494 40984 477500 40996
rect 337436 40956 477500 40984
rect 337436 40944 337442 40956
rect 477494 40944 477500 40956
rect 477552 40944 477558 40996
rect 333974 40876 333980 40928
rect 334032 40916 334038 40928
rect 510890 40916 510896 40928
rect 334032 40888 510896 40916
rect 334032 40876 334038 40888
rect 510890 40876 510896 40888
rect 510948 40876 510954 40928
rect 131114 40808 131120 40860
rect 131172 40848 131178 40860
rect 300118 40848 300124 40860
rect 131172 40820 300124 40848
rect 131172 40808 131178 40820
rect 300118 40808 300124 40820
rect 300176 40808 300182 40860
rect 329282 40808 329288 40860
rect 329340 40848 329346 40860
rect 506474 40848 506480 40860
rect 329340 40820 506480 40848
rect 329340 40808 329346 40820
rect 506474 40808 506480 40820
rect 506532 40808 506538 40860
rect 215294 40740 215300 40792
rect 215352 40780 215358 40792
rect 412634 40780 412640 40792
rect 215352 40752 412640 40780
rect 215352 40740 215358 40752
rect 412634 40740 412640 40752
rect 412692 40740 412698 40792
rect 27614 40672 27620 40724
rect 27672 40712 27678 40724
rect 125042 40712 125048 40724
rect 27672 40684 125048 40712
rect 27672 40672 27678 40684
rect 125042 40672 125048 40684
rect 125100 40672 125106 40724
rect 182174 40672 182180 40724
rect 182232 40712 182238 40724
rect 554774 40712 554780 40724
rect 182232 40684 554780 40712
rect 182232 40672 182238 40684
rect 554774 40672 554780 40684
rect 554832 40672 554838 40724
rect 251266 39652 251272 39704
rect 251324 39692 251330 39704
rect 402974 39692 402980 39704
rect 251324 39664 402980 39692
rect 251324 39652 251330 39664
rect 402974 39652 402980 39664
rect 403032 39652 403038 39704
rect 224678 39584 224684 39636
rect 224736 39624 224742 39636
rect 393314 39624 393320 39636
rect 224736 39596 393320 39624
rect 224736 39584 224742 39596
rect 393314 39584 393320 39596
rect 393372 39584 393378 39636
rect 327718 39516 327724 39568
rect 327776 39556 327782 39568
rect 509234 39556 509240 39568
rect 327776 39528 509240 39556
rect 327776 39516 327782 39528
rect 509234 39516 509240 39528
rect 509292 39516 509298 39568
rect 327074 39448 327080 39500
rect 327132 39488 327138 39500
rect 511994 39488 512000 39500
rect 327132 39460 512000 39488
rect 327132 39448 327138 39460
rect 511994 39448 512000 39460
rect 512052 39448 512058 39500
rect 151906 39380 151912 39432
rect 151964 39420 151970 39432
rect 431954 39420 431960 39432
rect 151964 39392 431960 39420
rect 151964 39380 151970 39392
rect 431954 39380 431960 39392
rect 432012 39380 432018 39432
rect 52546 39312 52552 39364
rect 52604 39352 52610 39364
rect 84838 39352 84844 39364
rect 52604 39324 84844 39352
rect 52604 39312 52610 39324
rect 84838 39312 84844 39324
rect 84896 39312 84902 39364
rect 178034 39312 178040 39364
rect 178092 39352 178098 39364
rect 556338 39352 556344 39364
rect 178092 39324 556344 39352
rect 178092 39312 178098 39324
rect 556338 39312 556344 39324
rect 556396 39312 556402 39364
rect 253934 38224 253940 38276
rect 253992 38264 253998 38276
rect 401594 38264 401600 38276
rect 253992 38236 401600 38264
rect 253992 38224 253998 38236
rect 401594 38224 401600 38236
rect 401652 38224 401658 38276
rect 220630 38156 220636 38208
rect 220688 38196 220694 38208
rect 407114 38196 407120 38208
rect 220688 38168 407120 38196
rect 220688 38156 220694 38168
rect 407114 38156 407120 38168
rect 407172 38156 407178 38208
rect 324314 38088 324320 38140
rect 324372 38128 324378 38140
rect 513466 38128 513472 38140
rect 324372 38100 513472 38128
rect 324372 38088 324378 38100
rect 513466 38088 513472 38100
rect 513524 38088 513530 38140
rect 322198 38020 322204 38072
rect 322256 38060 322262 38072
rect 527174 38060 527180 38072
rect 322256 38032 527180 38060
rect 322256 38020 322262 38032
rect 527174 38020 527180 38032
rect 527232 38020 527238 38072
rect 158714 37952 158720 38004
rect 158772 37992 158778 38004
rect 429194 37992 429200 38004
rect 158772 37964 429200 37992
rect 158772 37952 158778 37964
rect 429194 37952 429200 37964
rect 429252 37952 429258 38004
rect 448514 37952 448520 38004
rect 448572 37992 448578 38004
rect 477770 37992 477776 38004
rect 448572 37964 477776 37992
rect 448572 37952 448578 37964
rect 477770 37952 477776 37964
rect 477828 37952 477834 38004
rect 20714 37884 20720 37936
rect 20772 37924 20778 37936
rect 159358 37924 159364 37936
rect 20772 37896 159364 37924
rect 20772 37884 20778 37896
rect 159358 37884 159364 37896
rect 159416 37884 159422 37936
rect 175274 37884 175280 37936
rect 175332 37924 175338 37936
rect 556522 37924 556528 37936
rect 175332 37896 556528 37924
rect 175332 37884 175338 37896
rect 556522 37884 556528 37896
rect 556580 37884 556586 37936
rect 230382 36796 230388 36848
rect 230440 36836 230446 36848
rect 372614 36836 372620 36848
rect 230440 36808 372620 36836
rect 230440 36796 230446 36808
rect 372614 36796 372620 36808
rect 372672 36796 372678 36848
rect 292666 36728 292672 36780
rect 292724 36768 292730 36780
rect 523218 36768 523224 36780
rect 292724 36740 523224 36768
rect 292724 36728 292730 36740
rect 523218 36728 523224 36740
rect 523276 36728 523282 36780
rect 249610 36660 249616 36712
rect 249668 36700 249674 36712
rect 304994 36700 305000 36712
rect 249668 36672 305000 36700
rect 249668 36660 249674 36672
rect 304994 36660 305000 36672
rect 305052 36660 305058 36712
rect 310422 36660 310428 36712
rect 310480 36700 310486 36712
rect 552014 36700 552020 36712
rect 310480 36672 552020 36700
rect 310480 36660 310486 36672
rect 552014 36660 552020 36672
rect 552072 36660 552078 36712
rect 136634 36592 136640 36644
rect 136692 36632 136698 36644
rect 436370 36632 436376 36644
rect 136692 36604 436376 36632
rect 136692 36592 136698 36604
rect 436370 36592 436376 36604
rect 436428 36592 436434 36644
rect 444374 36592 444380 36644
rect 444432 36632 444438 36644
rect 477586 36632 477592 36644
rect 444432 36604 477592 36632
rect 444432 36592 444438 36604
rect 477586 36592 477592 36604
rect 477644 36592 477650 36644
rect 171134 36524 171140 36576
rect 171192 36564 171198 36576
rect 557626 36564 557632 36576
rect 171192 36536 557632 36564
rect 171192 36524 171198 36536
rect 557626 36524 557632 36536
rect 557684 36524 557690 36576
rect 364978 35572 364984 35624
rect 365036 35612 365042 35624
rect 382550 35612 382556 35624
rect 365036 35584 382556 35612
rect 365036 35572 365042 35584
rect 382550 35572 382556 35584
rect 382608 35572 382614 35624
rect 332594 35504 332600 35556
rect 332652 35544 332658 35556
rect 378226 35544 378232 35556
rect 332652 35516 378232 35544
rect 332652 35504 332658 35516
rect 378226 35504 378232 35516
rect 378284 35504 378290 35556
rect 352558 35436 352564 35488
rect 352616 35476 352622 35488
rect 423950 35476 423956 35488
rect 352616 35448 423956 35476
rect 352616 35436 352622 35448
rect 423950 35436 423956 35448
rect 424008 35436 424014 35488
rect 231762 35368 231768 35420
rect 231820 35408 231826 35420
rect 368474 35408 368480 35420
rect 231820 35380 368480 35408
rect 231820 35368 231826 35380
rect 368474 35368 368480 35380
rect 368532 35368 368538 35420
rect 423766 35368 423772 35420
rect 423824 35408 423830 35420
rect 484486 35408 484492 35420
rect 423824 35380 484492 35408
rect 423824 35368 423830 35380
rect 484486 35368 484492 35380
rect 484544 35368 484550 35420
rect 179414 35300 179420 35352
rect 179472 35340 179478 35352
rect 423674 35340 423680 35352
rect 179472 35312 423680 35340
rect 179472 35300 179478 35312
rect 423674 35300 423680 35312
rect 423732 35300 423738 35352
rect 446398 35300 446404 35352
rect 446456 35340 446462 35352
rect 554774 35340 554780 35352
rect 446456 35312 554780 35340
rect 446456 35300 446462 35312
rect 554774 35300 554780 35312
rect 554832 35300 554838 35352
rect 256694 35232 256700 35284
rect 256752 35272 256758 35284
rect 532694 35272 532700 35284
rect 256752 35244 532700 35272
rect 256752 35232 256758 35244
rect 532694 35232 532700 35244
rect 532752 35232 532758 35284
rect 153194 35164 153200 35216
rect 153252 35204 153258 35216
rect 563054 35204 563060 35216
rect 153252 35176 563060 35204
rect 153252 35164 153258 35176
rect 563054 35164 563060 35176
rect 563112 35164 563118 35216
rect 358262 34076 358268 34128
rect 358320 34116 358326 34128
rect 402974 34116 402980 34128
rect 358320 34088 402980 34116
rect 358320 34076 358326 34088
rect 402974 34076 402980 34088
rect 403032 34076 403038 34128
rect 317414 34008 317420 34060
rect 317472 34048 317478 34060
rect 382274 34048 382280 34060
rect 317472 34020 382280 34048
rect 317472 34008 317478 34020
rect 382274 34008 382280 34020
rect 382332 34008 382338 34060
rect 190454 33940 190460 33992
rect 190512 33980 190518 33992
rect 419810 33980 419816 33992
rect 190512 33952 419816 33980
rect 190512 33940 190518 33952
rect 419810 33940 419816 33952
rect 419868 33940 419874 33992
rect 447778 33940 447784 33992
rect 447836 33980 447842 33992
rect 550634 33980 550640 33992
rect 447836 33952 550640 33980
rect 447836 33940 447842 33952
rect 550634 33940 550640 33952
rect 550692 33940 550698 33992
rect 252554 33872 252560 33924
rect 252612 33912 252618 33924
rect 534074 33912 534080 33924
rect 252612 33884 534080 33912
rect 252612 33872 252618 33884
rect 534074 33872 534080 33884
rect 534132 33872 534138 33924
rect 51074 33804 51080 33856
rect 51132 33844 51138 33856
rect 151078 33844 151084 33856
rect 51132 33816 151084 33844
rect 51132 33804 51138 33816
rect 151078 33804 151084 33816
rect 151136 33804 151142 33856
rect 180702 33804 180708 33856
rect 180760 33844 180766 33856
rect 542354 33844 542360 33856
rect 180760 33816 542360 33844
rect 180760 33804 180766 33816
rect 542354 33804 542360 33816
rect 542412 33804 542418 33856
rect 150434 33736 150440 33788
rect 150492 33776 150498 33788
rect 564618 33776 564624 33788
rect 150492 33748 564624 33776
rect 150492 33736 150498 33748
rect 564618 33736 564624 33748
rect 564676 33736 564682 33788
rect 289814 32716 289820 32768
rect 289872 32756 289878 32768
rect 390830 32756 390836 32768
rect 289872 32728 390836 32756
rect 289872 32716 289878 32728
rect 390830 32716 390836 32728
rect 390888 32716 390894 32768
rect 356698 32648 356704 32700
rect 356756 32688 356762 32700
rect 409874 32688 409880 32700
rect 356756 32660 409880 32688
rect 356756 32648 356762 32660
rect 409874 32648 409880 32660
rect 409932 32648 409938 32700
rect 224862 32580 224868 32632
rect 224920 32620 224926 32632
rect 390554 32620 390560 32632
rect 224920 32592 390560 32620
rect 224920 32580 224926 32592
rect 390554 32580 390560 32592
rect 390612 32580 390618 32632
rect 437474 32580 437480 32632
rect 437532 32620 437538 32632
rect 480254 32620 480260 32632
rect 437532 32592 480260 32620
rect 437532 32580 437538 32592
rect 480254 32580 480260 32592
rect 480312 32580 480318 32632
rect 212534 32512 212540 32564
rect 212592 32552 212598 32564
rect 276658 32552 276664 32564
rect 212592 32524 276664 32552
rect 212592 32512 212598 32524
rect 276658 32512 276664 32524
rect 276716 32512 276722 32564
rect 277394 32512 277400 32564
rect 277452 32552 277458 32564
rect 527358 32552 527364 32564
rect 277452 32524 527364 32552
rect 277452 32512 277458 32524
rect 527358 32512 527364 32524
rect 527416 32512 527422 32564
rect 184934 32444 184940 32496
rect 184992 32484 184998 32496
rect 284938 32484 284944 32496
rect 184992 32456 284944 32484
rect 184992 32444 184998 32456
rect 284938 32444 284944 32456
rect 284996 32444 285002 32496
rect 307570 32444 307576 32496
rect 307628 32484 307634 32496
rect 563054 32484 563060 32496
rect 307628 32456 563060 32484
rect 307628 32444 307634 32456
rect 563054 32444 563060 32456
rect 563112 32444 563118 32496
rect 26234 32376 26240 32428
rect 26292 32416 26298 32428
rect 158162 32416 158168 32428
rect 26292 32388 158168 32416
rect 26292 32376 26298 32388
rect 158162 32376 158168 32388
rect 158220 32376 158226 32428
rect 164234 32376 164240 32428
rect 164292 32416 164298 32428
rect 560386 32416 560392 32428
rect 164292 32388 560392 32416
rect 164292 32376 164298 32388
rect 560386 32376 560392 32388
rect 560444 32376 560450 32428
rect 296714 31288 296720 31340
rect 296772 31328 296778 31340
rect 389266 31328 389272 31340
rect 296772 31300 389272 31328
rect 296772 31288 296778 31300
rect 389266 31288 389272 31300
rect 389324 31288 389330 31340
rect 398834 31288 398840 31340
rect 398892 31328 398898 31340
rect 491294 31328 491300 31340
rect 398892 31300 491300 31328
rect 398892 31288 398898 31300
rect 491294 31288 491300 31300
rect 491352 31288 491358 31340
rect 149054 31220 149060 31272
rect 149112 31260 149118 31272
rect 294598 31260 294604 31272
rect 149112 31232 294604 31260
rect 149112 31220 149118 31232
rect 294598 31220 294604 31232
rect 294656 31220 294662 31272
rect 303338 31220 303344 31272
rect 303396 31260 303402 31272
rect 576118 31260 576124 31272
rect 303396 31232 576124 31260
rect 303396 31220 303402 31232
rect 576118 31220 576124 31232
rect 576176 31220 576182 31272
rect 242894 31152 242900 31204
rect 242952 31192 242958 31204
rect 536926 31192 536932 31204
rect 242952 31164 536932 31192
rect 242952 31152 242958 31164
rect 536926 31152 536932 31164
rect 536984 31152 536990 31204
rect 126974 31084 126980 31136
rect 127032 31124 127038 31136
rect 438854 31124 438860 31136
rect 127032 31096 438860 31124
rect 127032 31084 127038 31096
rect 438854 31084 438860 31096
rect 438912 31084 438918 31136
rect 449342 31084 449348 31136
rect 449400 31124 449406 31136
rect 547874 31124 547880 31136
rect 449400 31096 547880 31124
rect 449400 31084 449406 31096
rect 547874 31084 547880 31096
rect 547932 31084 547938 31136
rect 41414 31016 41420 31068
rect 41472 31056 41478 31068
rect 120902 31056 120908 31068
rect 41472 31028 120908 31056
rect 41472 31016 41478 31028
rect 120902 31016 120908 31028
rect 120960 31016 120966 31068
rect 179046 31016 179052 31068
rect 179104 31056 179110 31068
rect 547138 31056 547144 31068
rect 179104 31028 547144 31056
rect 179104 31016 179110 31028
rect 547138 31016 547144 31028
rect 547196 31016 547202 31068
rect 394694 29928 394700 29980
rect 394752 29968 394758 29980
rect 492674 29968 492680 29980
rect 394752 29940 492680 29968
rect 394752 29928 394758 29940
rect 492674 29928 492680 29940
rect 492732 29928 492738 29980
rect 260834 29860 260840 29912
rect 260892 29900 260898 29912
rect 399110 29900 399116 29912
rect 260892 29872 399116 29900
rect 260892 29860 260898 29872
rect 399110 29860 399116 29872
rect 399168 29860 399174 29912
rect 330478 29792 330484 29844
rect 330536 29832 330542 29844
rect 498194 29832 498200 29844
rect 330536 29804 498200 29832
rect 330536 29792 330542 29804
rect 498194 29792 498200 29804
rect 498252 29792 498258 29844
rect 165614 29724 165620 29776
rect 165672 29764 165678 29776
rect 427998 29764 428004 29776
rect 165672 29736 428004 29764
rect 165672 29724 165678 29736
rect 427998 29724 428004 29736
rect 428056 29724 428062 29776
rect 449158 29724 449164 29776
rect 449216 29764 449222 29776
rect 543734 29764 543740 29776
rect 449216 29736 543740 29764
rect 449216 29724 449222 29736
rect 543734 29724 543740 29736
rect 543792 29724 543798 29776
rect 224954 29656 224960 29708
rect 225012 29696 225018 29708
rect 542446 29696 542452 29708
rect 225012 29668 542452 29696
rect 225012 29656 225018 29668
rect 542446 29656 542452 29668
rect 542504 29656 542510 29708
rect 34514 29588 34520 29640
rect 34572 29628 34578 29640
rect 122098 29628 122104 29640
rect 34572 29600 122104 29628
rect 34572 29588 34578 29600
rect 122098 29588 122104 29600
rect 122156 29588 122162 29640
rect 183186 29588 183192 29640
rect 183244 29628 183250 29640
rect 535454 29628 535460 29640
rect 183244 29600 535460 29628
rect 183244 29588 183250 29600
rect 535454 29588 535460 29600
rect 535512 29588 535518 29640
rect 387794 28568 387800 28620
rect 387852 28608 387858 28620
rect 494054 28608 494060 28620
rect 387852 28580 494060 28608
rect 387852 28568 387858 28580
rect 494054 28568 494060 28580
rect 494112 28568 494118 28620
rect 271874 28500 271880 28552
rect 271932 28540 271938 28552
rect 396074 28540 396080 28552
rect 271932 28512 396080 28540
rect 271932 28500 271938 28512
rect 396074 28500 396080 28512
rect 396132 28500 396138 28552
rect 329098 28432 329104 28484
rect 329156 28472 329162 28484
rect 502334 28472 502340 28484
rect 329156 28444 502340 28472
rect 329156 28432 329162 28444
rect 502334 28432 502340 28444
rect 502392 28432 502398 28484
rect 172514 28364 172520 28416
rect 172572 28404 172578 28416
rect 425146 28404 425152 28416
rect 172572 28376 425152 28404
rect 172572 28364 172578 28376
rect 425146 28364 425152 28376
rect 425204 28364 425210 28416
rect 450538 28364 450544 28416
rect 450596 28404 450602 28416
rect 539870 28404 539876 28416
rect 450596 28376 539876 28404
rect 450596 28364 450602 28376
rect 539870 28364 539876 28376
rect 539928 28364 539934 28416
rect 220814 28296 220820 28348
rect 220872 28336 220878 28348
rect 544010 28336 544016 28348
rect 220872 28308 544016 28336
rect 220872 28296 220878 28308
rect 544010 28296 544016 28308
rect 544068 28296 544074 28348
rect 16574 28228 16580 28280
rect 16632 28268 16638 28280
rect 160738 28268 160744 28280
rect 16632 28240 160744 28268
rect 16632 28228 16638 28240
rect 160738 28228 160744 28240
rect 160796 28228 160802 28280
rect 182082 28228 182088 28280
rect 182140 28268 182146 28280
rect 538858 28268 538864 28280
rect 182140 28240 538864 28268
rect 182140 28228 182146 28240
rect 538858 28228 538864 28240
rect 538916 28228 538922 28280
rect 187694 27208 187700 27260
rect 187752 27248 187758 27260
rect 283558 27248 283564 27260
rect 187752 27220 283564 27248
rect 187752 27208 187758 27220
rect 283558 27208 283564 27220
rect 283616 27208 283622 27260
rect 353938 27208 353944 27260
rect 353996 27248 354002 27260
rect 416774 27248 416780 27260
rect 353996 27220 416780 27248
rect 353996 27208 354002 27220
rect 416774 27208 416780 27220
rect 416832 27208 416838 27260
rect 282914 27140 282920 27192
rect 282972 27180 282978 27192
rect 393406 27180 393412 27192
rect 282972 27152 393412 27180
rect 282972 27140 282978 27152
rect 393406 27140 393412 27152
rect 393464 27140 393470 27192
rect 217962 27072 217968 27124
rect 218020 27112 218026 27124
rect 415394 27112 415400 27124
rect 218020 27084 415400 27112
rect 218020 27072 218026 27084
rect 415394 27072 415400 27084
rect 415452 27072 415458 27124
rect 433334 27072 433340 27124
rect 433392 27112 433398 27124
rect 481818 27112 481824 27124
rect 433392 27084 481824 27112
rect 433392 27072 433398 27084
rect 481818 27072 481824 27084
rect 481876 27072 481882 27124
rect 270494 27004 270500 27056
rect 270552 27044 270558 27056
rect 528554 27044 528560 27056
rect 270552 27016 528560 27044
rect 270552 27004 270558 27016
rect 528554 27004 528560 27016
rect 528612 27004 528618 27056
rect 135346 26936 135352 26988
rect 135404 26976 135410 26988
rect 298738 26976 298744 26988
rect 135404 26948 298744 26976
rect 135404 26936 135410 26948
rect 298738 26936 298744 26948
rect 298796 26936 298802 26988
rect 306282 26936 306288 26988
rect 306340 26976 306346 26988
rect 565814 26976 565820 26988
rect 306340 26948 565820 26976
rect 306340 26936 306346 26948
rect 565814 26936 565820 26948
rect 565872 26936 565878 26988
rect 17954 26868 17960 26920
rect 18012 26908 18018 26920
rect 126238 26908 126244 26920
rect 18012 26880 126244 26908
rect 18012 26868 18018 26880
rect 126238 26868 126244 26880
rect 126296 26868 126302 26920
rect 160094 26868 160100 26920
rect 160152 26908 160158 26920
rect 560570 26908 560576 26920
rect 160152 26880 560576 26908
rect 160152 26868 160158 26880
rect 560570 26868 560576 26880
rect 560628 26868 560634 26920
rect 307754 25848 307760 25900
rect 307812 25888 307818 25900
rect 386598 25888 386604 25900
rect 307812 25860 386604 25888
rect 307812 25848 307818 25860
rect 386598 25848 386604 25860
rect 386656 25848 386662 25900
rect 383654 25780 383660 25832
rect 383712 25820 383718 25832
rect 495526 25820 495532 25832
rect 383712 25792 495532 25820
rect 383712 25780 383718 25792
rect 495526 25780 495532 25792
rect 495584 25780 495590 25832
rect 235994 25712 236000 25764
rect 236052 25752 236058 25764
rect 407298 25752 407304 25764
rect 236052 25724 407304 25752
rect 236052 25712 236058 25724
rect 407298 25712 407304 25724
rect 407356 25712 407362 25764
rect 461762 25712 461768 25764
rect 461820 25752 461826 25764
rect 500954 25752 500960 25764
rect 461820 25724 500960 25752
rect 461820 25712 461826 25724
rect 500954 25712 500960 25724
rect 501012 25712 501018 25764
rect 202874 25644 202880 25696
rect 202932 25684 202938 25696
rect 548058 25684 548064 25696
rect 202932 25656 548064 25684
rect 202932 25644 202938 25656
rect 548058 25644 548064 25656
rect 548116 25644 548122 25696
rect 28994 25576 29000 25628
rect 29052 25616 29058 25628
rect 157978 25616 157984 25628
rect 29052 25588 157984 25616
rect 29052 25576 29058 25588
rect 157978 25576 157984 25588
rect 158036 25576 158042 25628
rect 177942 25576 177948 25628
rect 178000 25616 178006 25628
rect 553486 25616 553492 25628
rect 178000 25588 553492 25616
rect 178000 25576 178006 25588
rect 553486 25576 553492 25588
rect 553544 25576 553550 25628
rect 157334 25508 157340 25560
rect 157392 25548 157398 25560
rect 561766 25548 561772 25560
rect 157392 25520 561772 25548
rect 157392 25508 157398 25520
rect 561766 25508 561772 25520
rect 561824 25508 561830 25560
rect 278774 24420 278780 24472
rect 278832 24460 278838 24472
rect 394878 24460 394884 24472
rect 278832 24432 394884 24460
rect 278832 24420 278838 24432
rect 394878 24420 394884 24432
rect 394936 24420 394942 24472
rect 376754 24352 376760 24404
rect 376812 24392 376818 24404
rect 498378 24392 498384 24404
rect 376812 24364 498384 24392
rect 376812 24352 376818 24364
rect 498378 24352 498384 24364
rect 498436 24352 498442 24404
rect 333238 24284 333244 24336
rect 333296 24324 333302 24336
rect 491294 24324 491300 24336
rect 333296 24296 491300 24324
rect 333296 24284 333302 24296
rect 491294 24284 491300 24296
rect 491352 24284 491358 24336
rect 176654 24216 176660 24268
rect 176712 24256 176718 24268
rect 423858 24256 423864 24268
rect 176712 24228 423864 24256
rect 176712 24216 176718 24228
rect 423858 24216 423864 24228
rect 423916 24216 423922 24268
rect 464338 24216 464344 24268
rect 464396 24256 464402 24268
rect 494054 24256 494060 24268
rect 464396 24228 494060 24256
rect 464396 24216 464402 24228
rect 494054 24216 494060 24228
rect 494112 24216 494118 24268
rect 184842 24148 184848 24200
rect 184900 24188 184906 24200
rect 528554 24188 528560 24200
rect 184900 24160 528560 24188
rect 184900 24148 184906 24160
rect 528554 24148 528560 24160
rect 528612 24148 528618 24200
rect 74442 24080 74448 24132
rect 74500 24120 74506 24132
rect 88334 24120 88340 24132
rect 74500 24092 88340 24120
rect 74500 24080 74506 24092
rect 88334 24080 88340 24092
rect 88392 24080 88398 24132
rect 185026 24080 185032 24132
rect 185084 24120 185090 24132
rect 553394 24120 553400 24132
rect 185084 24092 553400 24120
rect 185084 24080 185090 24092
rect 553394 24080 553400 24092
rect 553452 24080 553458 24132
rect 97994 23808 98000 23860
rect 98052 23848 98058 23860
rect 104158 23848 104164 23860
rect 98052 23820 104164 23848
rect 98052 23808 98058 23820
rect 104158 23808 104164 23820
rect 104216 23808 104222 23860
rect 194594 23060 194600 23112
rect 194652 23100 194658 23112
rect 282362 23100 282368 23112
rect 194652 23072 282368 23100
rect 194652 23060 194658 23072
rect 282362 23060 282368 23072
rect 282420 23060 282426 23112
rect 357434 23060 357440 23112
rect 357492 23100 357498 23112
rect 371234 23100 371240 23112
rect 357492 23072 371240 23100
rect 357492 23060 357498 23072
rect 371234 23060 371240 23072
rect 371292 23060 371298 23112
rect 264974 22992 264980 23044
rect 265032 23032 265038 23044
rect 398926 23032 398932 23044
rect 265032 23004 398932 23032
rect 265032 22992 265038 23004
rect 398926 22992 398932 23004
rect 398984 22992 398990 23044
rect 223482 22924 223488 22976
rect 223540 22964 223546 22976
rect 397454 22964 397460 22976
rect 223540 22936 397460 22964
rect 223540 22924 223546 22936
rect 397454 22924 397460 22936
rect 397512 22924 397518 22976
rect 426434 22924 426440 22976
rect 426492 22964 426498 22976
rect 483014 22964 483020 22976
rect 426492 22936 483020 22964
rect 426492 22924 426498 22936
rect 483014 22924 483020 22936
rect 483072 22924 483078 22976
rect 267826 22856 267832 22908
rect 267884 22896 267890 22908
rect 529934 22896 529940 22908
rect 267884 22868 529940 22896
rect 267884 22856 267890 22868
rect 529934 22856 529940 22868
rect 529992 22856 529998 22908
rect 144914 22788 144920 22840
rect 144972 22828 144978 22840
rect 295978 22828 295984 22840
rect 144972 22800 295984 22828
rect 144972 22788 144978 22800
rect 295978 22788 295984 22800
rect 296036 22788 296042 22840
rect 304902 22788 304908 22840
rect 304960 22828 304966 22840
rect 569954 22828 569960 22840
rect 304960 22800 569960 22828
rect 304960 22788 304966 22800
rect 569954 22788 569960 22800
rect 570012 22788 570018 22840
rect 77294 22720 77300 22772
rect 77352 22760 77358 22772
rect 109678 22760 109684 22772
rect 77352 22732 109684 22760
rect 77352 22720 77358 22732
rect 109678 22720 109684 22732
rect 109736 22720 109742 22772
rect 125594 22720 125600 22772
rect 125652 22760 125658 22772
rect 571334 22760 571340 22772
rect 125652 22732 571340 22760
rect 125652 22720 125658 22732
rect 571334 22720 571340 22732
rect 571392 22720 571398 22772
rect 349246 21700 349252 21752
rect 349304 21740 349310 21752
rect 374086 21740 374092 21752
rect 349304 21712 374092 21740
rect 349304 21700 349310 21712
rect 374086 21700 374092 21712
rect 374144 21700 374150 21752
rect 220446 21632 220452 21684
rect 220504 21672 220510 21684
rect 404354 21672 404360 21684
rect 220504 21644 404360 21672
rect 220504 21632 220510 21644
rect 404354 21632 404360 21644
rect 404412 21632 404418 21684
rect 408494 21632 408500 21684
rect 408552 21672 408558 21684
rect 488626 21672 488632 21684
rect 408552 21644 488632 21672
rect 408552 21632 408558 21644
rect 488626 21632 488632 21644
rect 488684 21632 488690 21684
rect 216306 21564 216312 21616
rect 216364 21604 216370 21616
rect 422294 21604 422300 21616
rect 216364 21576 422300 21604
rect 216364 21564 216370 21576
rect 422294 21564 422300 21576
rect 422352 21564 422358 21616
rect 213822 21496 213828 21548
rect 213880 21536 213886 21548
rect 429194 21536 429200 21548
rect 213880 21508 429200 21536
rect 213880 21496 213886 21508
rect 429194 21496 429200 21508
rect 429252 21496 429258 21548
rect 462314 21496 462320 21548
rect 462372 21536 462378 21548
rect 473538 21536 473544 21548
rect 462372 21508 473544 21536
rect 462372 21496 462378 21508
rect 473538 21496 473544 21508
rect 473596 21496 473602 21548
rect 212350 21428 212356 21480
rect 212408 21468 212414 21480
rect 431954 21468 431960 21480
rect 212408 21440 431960 21468
rect 212408 21428 212414 21440
rect 431954 21428 431960 21440
rect 432012 21428 432018 21480
rect 465902 21428 465908 21480
rect 465960 21468 465966 21480
rect 490190 21468 490196 21480
rect 465960 21440 490196 21468
rect 465960 21428 465966 21440
rect 490190 21428 490196 21440
rect 490248 21428 490254 21480
rect 35894 21360 35900 21412
rect 35952 21400 35958 21412
rect 155218 21400 155224 21412
rect 35952 21372 155224 21400
rect 35952 21360 35958 21372
rect 155218 21360 155224 21372
rect 155276 21360 155282 21412
rect 212166 21360 212172 21412
rect 212224 21400 212230 21412
rect 436094 21400 436100 21412
rect 212224 21372 436100 21400
rect 212224 21360 212230 21372
rect 436094 21360 436100 21372
rect 436152 21360 436158 21412
rect 443638 21360 443644 21412
rect 443696 21400 443702 21412
rect 564434 21400 564440 21412
rect 443696 21372 564440 21400
rect 443696 21360 443702 21372
rect 564434 21360 564440 21372
rect 564492 21360 564498 21412
rect 228726 20408 228732 20460
rect 228784 20448 228790 20460
rect 375374 20448 375380 20460
rect 228784 20420 375380 20448
rect 228784 20408 228790 20420
rect 375374 20408 375380 20420
rect 375432 20408 375438 20460
rect 227622 20340 227628 20392
rect 227680 20380 227686 20392
rect 382366 20380 382372 20392
rect 227680 20352 382372 20380
rect 227680 20340 227686 20352
rect 382366 20340 382372 20352
rect 382424 20340 382430 20392
rect 176562 20272 176568 20324
rect 176620 20312 176626 20324
rect 556246 20312 556252 20324
rect 176620 20284 556252 20312
rect 176620 20272 176626 20284
rect 556246 20272 556252 20284
rect 556304 20272 556310 20324
rect 175090 20204 175096 20256
rect 175148 20244 175154 20256
rect 560294 20244 560300 20256
rect 175148 20216 560300 20244
rect 175148 20204 175154 20216
rect 560294 20204 560300 20216
rect 560352 20204 560358 20256
rect 174906 20136 174912 20188
rect 174964 20176 174970 20188
rect 564526 20176 564532 20188
rect 174964 20148 564532 20176
rect 174964 20136 174970 20148
rect 564526 20136 564532 20148
rect 564584 20136 564590 20188
rect 172422 20068 172428 20120
rect 172480 20108 172486 20120
rect 571334 20108 571340 20120
rect 172480 20080 571340 20108
rect 172480 20068 172486 20080
rect 571334 20068 571340 20080
rect 571392 20068 571398 20120
rect 170766 20000 170772 20052
rect 170824 20040 170830 20052
rect 574094 20040 574100 20052
rect 170824 20012 574100 20040
rect 170824 20000 170830 20012
rect 574094 20000 574100 20012
rect 574152 20000 574158 20052
rect 33134 19932 33140 19984
rect 33192 19972 33198 19984
rect 156598 19972 156604 19984
rect 33192 19944 156604 19972
rect 33192 19932 33198 19944
rect 156598 19932 156604 19944
rect 156656 19932 156662 19984
rect 170950 19932 170956 19984
rect 171008 19972 171014 19984
rect 578234 19972 578240 19984
rect 171008 19944 578240 19972
rect 171008 19932 171014 19944
rect 578234 19932 578240 19944
rect 578292 19932 578298 19984
rect 195790 19116 195796 19168
rect 195848 19156 195854 19168
rect 490006 19156 490012 19168
rect 195848 19128 490012 19156
rect 195848 19116 195854 19128
rect 490006 19116 490012 19128
rect 490064 19116 490070 19168
rect 195606 19048 195612 19100
rect 195664 19088 195670 19100
rect 492674 19088 492680 19100
rect 195664 19060 492680 19088
rect 195664 19048 195670 19060
rect 492674 19048 492680 19060
rect 492732 19048 492738 19100
rect 194502 18980 194508 19032
rect 194560 19020 194566 19032
rect 496906 19020 496912 19032
rect 194560 18992 496912 19020
rect 194560 18980 194566 18992
rect 496906 18980 496912 18992
rect 496964 18980 496970 19032
rect 193122 18912 193128 18964
rect 193180 18952 193186 18964
rect 499574 18952 499580 18964
rect 193180 18924 499580 18952
rect 193180 18912 193186 18924
rect 499574 18912 499580 18924
rect 499632 18912 499638 18964
rect 191650 18844 191656 18896
rect 191708 18884 191714 18896
rect 503714 18884 503720 18896
rect 191708 18856 503720 18884
rect 191708 18844 191714 18856
rect 503714 18844 503720 18856
rect 503772 18844 503778 18896
rect 191466 18776 191472 18828
rect 191524 18816 191530 18828
rect 506566 18816 506572 18828
rect 191524 18788 506572 18816
rect 191524 18776 191530 18788
rect 506566 18776 506572 18788
rect 506624 18776 506630 18828
rect 190362 18708 190368 18760
rect 190420 18748 190426 18760
rect 510614 18748 510620 18760
rect 190420 18720 510620 18748
rect 190420 18708 190426 18720
rect 510614 18708 510620 18720
rect 510672 18708 510678 18760
rect 187510 18640 187516 18692
rect 187568 18680 187574 18692
rect 517514 18680 517520 18692
rect 187568 18652 517520 18680
rect 187568 18640 187574 18652
rect 517514 18640 517520 18652
rect 517572 18640 517578 18692
rect 67634 18572 67640 18624
rect 67692 18612 67698 18624
rect 80882 18612 80888 18624
rect 67692 18584 80888 18612
rect 67692 18572 67698 18584
rect 80882 18572 80888 18584
rect 80940 18572 80946 18624
rect 86954 18572 86960 18624
rect 87012 18612 87018 18624
rect 106918 18612 106924 18624
rect 87012 18584 106924 18612
rect 87012 18572 87018 18584
rect 106918 18572 106924 18584
rect 106976 18572 106982 18624
rect 107654 18572 107660 18624
rect 107712 18612 107718 18624
rect 134518 18612 134524 18624
rect 107712 18584 134524 18612
rect 107712 18572 107718 18584
rect 134518 18572 134524 18584
rect 134576 18572 134582 18624
rect 187326 18572 187332 18624
rect 187384 18612 187390 18624
rect 521654 18612 521660 18624
rect 187384 18584 521660 18612
rect 187384 18572 187390 18584
rect 521654 18572 521660 18584
rect 521712 18572 521718 18624
rect 351178 17824 351184 17876
rect 351236 17864 351242 17876
rect 427814 17864 427820 17876
rect 351236 17836 427820 17864
rect 351236 17824 351242 17836
rect 427814 17824 427820 17836
rect 427872 17824 427878 17876
rect 349798 17756 349804 17808
rect 349856 17796 349862 17808
rect 432046 17796 432052 17808
rect 349856 17768 432052 17796
rect 349856 17756 349862 17768
rect 432046 17756 432052 17768
rect 432104 17756 432110 17808
rect 349982 17688 349988 17740
rect 350040 17728 350046 17740
rect 434714 17728 434720 17740
rect 350040 17700 434720 17728
rect 350040 17688 350046 17700
rect 434714 17688 434720 17700
rect 434772 17688 434778 17740
rect 348418 17620 348424 17672
rect 348476 17660 348482 17672
rect 438854 17660 438860 17672
rect 348476 17632 438860 17660
rect 348476 17620 348482 17632
rect 438854 17620 438860 17632
rect 438912 17620 438918 17672
rect 440326 17620 440332 17672
rect 440384 17660 440390 17672
rect 478874 17660 478880 17672
rect 440384 17632 478880 17660
rect 440384 17620 440390 17632
rect 478874 17620 478880 17632
rect 478932 17620 478938 17672
rect 347038 17552 347044 17604
rect 347096 17592 347102 17604
rect 441614 17592 441620 17604
rect 347096 17564 441620 17592
rect 347096 17552 347102 17564
rect 441614 17552 441620 17564
rect 441672 17552 441678 17604
rect 251082 17484 251088 17536
rect 251140 17524 251146 17536
rect 300854 17524 300860 17536
rect 251140 17496 300860 17524
rect 251140 17484 251146 17496
rect 300854 17484 300860 17496
rect 300912 17484 300918 17536
rect 345658 17484 345664 17536
rect 345716 17524 345722 17536
rect 445754 17524 445760 17536
rect 345716 17496 445760 17524
rect 345716 17484 345722 17496
rect 445754 17484 445760 17496
rect 445812 17484 445818 17536
rect 209866 17416 209872 17468
rect 209924 17456 209930 17468
rect 278222 17456 278228 17468
rect 209924 17428 278228 17456
rect 209924 17416 209930 17428
rect 278222 17416 278228 17428
rect 278280 17416 278286 17468
rect 345842 17416 345848 17468
rect 345900 17456 345906 17468
rect 448606 17456 448612 17468
rect 345900 17428 448612 17456
rect 345900 17416 345906 17428
rect 448606 17416 448612 17428
rect 448664 17416 448670 17468
rect 451274 17416 451280 17468
rect 451332 17456 451338 17468
rect 476206 17456 476212 17468
rect 451332 17428 476212 17456
rect 451332 17416 451338 17428
rect 476206 17416 476212 17428
rect 476264 17416 476270 17468
rect 241146 17348 241152 17400
rect 241204 17388 241210 17400
rect 332686 17388 332692 17400
rect 241204 17360 332692 17388
rect 241204 17348 241210 17360
rect 332686 17348 332692 17360
rect 332744 17348 332750 17400
rect 344278 17348 344284 17400
rect 344336 17388 344342 17400
rect 452654 17388 452660 17400
rect 344336 17360 452660 17388
rect 344336 17348 344342 17360
rect 452654 17348 452660 17360
rect 452712 17348 452718 17400
rect 63494 17280 63500 17332
rect 63552 17320 63558 17332
rect 80698 17320 80704 17332
rect 63552 17292 80704 17320
rect 63552 17280 63558 17292
rect 80698 17280 80704 17292
rect 80756 17280 80762 17332
rect 169754 17280 169760 17332
rect 169812 17320 169818 17332
rect 289078 17320 289084 17332
rect 169812 17292 289084 17320
rect 169812 17280 169818 17292
rect 289078 17280 289084 17292
rect 289136 17280 289142 17332
rect 342898 17280 342904 17332
rect 342956 17320 342962 17332
rect 456886 17320 456892 17332
rect 342956 17292 456892 17320
rect 342956 17280 342962 17292
rect 456886 17280 456892 17292
rect 456944 17280 456950 17332
rect 465718 17280 465724 17332
rect 465776 17320 465782 17332
rect 487154 17320 487160 17332
rect 465776 17292 487160 17320
rect 465776 17280 465782 17292
rect 487154 17280 487160 17292
rect 487212 17280 487218 17332
rect 72878 17212 72884 17264
rect 72936 17252 72942 17264
rect 95234 17252 95240 17264
rect 72936 17224 95240 17252
rect 72936 17212 72942 17224
rect 95234 17212 95240 17224
rect 95292 17212 95298 17264
rect 100754 17212 100760 17264
rect 100812 17252 100818 17264
rect 137462 17252 137468 17264
rect 100812 17224 137468 17252
rect 100812 17212 100818 17224
rect 137462 17212 137468 17224
rect 137520 17212 137526 17264
rect 154574 17212 154580 17264
rect 154632 17252 154638 17264
rect 430666 17252 430672 17264
rect 154632 17224 430672 17252
rect 154632 17212 154638 17224
rect 430666 17212 430672 17224
rect 430724 17212 430730 17264
rect 456058 17212 456064 17264
rect 456116 17252 456122 17264
rect 523126 17252 523132 17264
rect 456116 17224 523132 17252
rect 456116 17212 456122 17224
rect 523126 17212 523132 17224
rect 523184 17212 523190 17264
rect 238662 16192 238668 16244
rect 238720 16232 238726 16244
rect 344554 16232 344560 16244
rect 238720 16204 344560 16232
rect 238720 16192 238726 16204
rect 344554 16192 344560 16204
rect 344612 16192 344618 16244
rect 366542 16192 366548 16244
rect 366600 16232 366606 16244
rect 374086 16232 374092 16244
rect 366600 16204 374092 16232
rect 366600 16192 366606 16204
rect 374086 16192 374092 16204
rect 374144 16192 374150 16244
rect 237190 16124 237196 16176
rect 237248 16164 237254 16176
rect 348050 16164 348056 16176
rect 237248 16136 348056 16164
rect 237248 16124 237254 16136
rect 348050 16124 348056 16136
rect 348108 16124 348114 16176
rect 363598 16124 363604 16176
rect 363656 16164 363662 16176
rect 385954 16164 385960 16176
rect 363656 16136 385960 16164
rect 363656 16124 363662 16136
rect 385954 16124 385960 16136
rect 386012 16124 386018 16176
rect 237006 16056 237012 16108
rect 237064 16096 237070 16108
rect 351178 16096 351184 16108
rect 237064 16068 351184 16096
rect 237064 16056 237070 16068
rect 351178 16056 351184 16068
rect 351236 16056 351242 16108
rect 360838 16056 360844 16108
rect 360896 16096 360902 16108
rect 396074 16096 396080 16108
rect 360896 16068 396080 16096
rect 360896 16056 360902 16068
rect 396074 16056 396080 16068
rect 396132 16056 396138 16108
rect 467098 16056 467104 16108
rect 467156 16096 467162 16108
rect 484026 16096 484032 16108
rect 467156 16068 484032 16096
rect 467156 16056 467162 16068
rect 484026 16056 484032 16068
rect 484084 16056 484090 16108
rect 234522 15988 234528 16040
rect 234580 16028 234586 16040
rect 357526 16028 357532 16040
rect 234580 16000 357532 16028
rect 234580 15988 234586 16000
rect 357526 15988 357532 16000
rect 357584 15988 357590 16040
rect 358078 15988 358084 16040
rect 358136 16028 358142 16040
rect 407206 16028 407212 16040
rect 358136 16000 407212 16028
rect 358136 15988 358142 16000
rect 407206 15988 407212 16000
rect 407264 15988 407270 16040
rect 420178 15988 420184 16040
rect 420236 16028 420242 16040
rect 485958 16028 485964 16040
rect 420236 16000 485964 16028
rect 420236 15988 420242 16000
rect 485958 15988 485964 16000
rect 486016 15988 486022 16040
rect 232866 15920 232872 15972
rect 232924 15960 232930 15972
rect 365714 15960 365720 15972
rect 232924 15932 365720 15960
rect 232924 15920 232930 15932
rect 365714 15920 365720 15932
rect 365772 15920 365778 15972
rect 366358 15920 366364 15972
rect 366416 15960 366422 15972
rect 378318 15960 378324 15972
rect 366416 15932 378324 15960
rect 366416 15920 366422 15932
rect 378318 15920 378324 15932
rect 378376 15920 378382 15972
rect 381170 15920 381176 15972
rect 381228 15960 381234 15972
rect 496814 15960 496820 15972
rect 381228 15932 496820 15960
rect 381228 15920 381234 15932
rect 496814 15920 496820 15932
rect 496872 15920 496878 15972
rect 73338 15852 73344 15904
rect 73396 15892 73402 15904
rect 111058 15892 111064 15904
rect 73396 15864 111064 15892
rect 73396 15852 73402 15864
rect 111058 15852 111064 15864
rect 111116 15852 111122 15904
rect 114738 15852 114744 15904
rect 114796 15892 114802 15904
rect 133138 15892 133144 15904
rect 114796 15864 133144 15892
rect 114796 15852 114802 15864
rect 133138 15852 133144 15864
rect 133196 15852 133202 15904
rect 147858 15852 147864 15904
rect 147916 15892 147922 15904
rect 432138 15892 432144 15904
rect 147916 15864 432144 15892
rect 147916 15852 147922 15864
rect 432138 15852 432144 15864
rect 432196 15852 432202 15904
rect 461578 15852 461584 15904
rect 461636 15892 461642 15904
rect 505370 15892 505376 15904
rect 461636 15864 505376 15892
rect 461636 15852 461642 15864
rect 505370 15852 505376 15864
rect 505428 15852 505434 15904
rect 367738 15308 367744 15360
rect 367796 15348 367802 15360
rect 371234 15348 371240 15360
rect 367796 15320 371240 15348
rect 367796 15308 367802 15320
rect 371234 15308 371240 15320
rect 371292 15308 371298 15360
rect 260742 14696 260748 14748
rect 260800 14736 260806 14748
rect 270034 14736 270040 14748
rect 260800 14708 270040 14736
rect 260800 14696 260806 14708
rect 270034 14696 270040 14708
rect 270092 14696 270098 14748
rect 320818 14696 320824 14748
rect 320876 14736 320882 14748
rect 534442 14736 534448 14748
rect 320876 14708 534448 14736
rect 320876 14696 320882 14708
rect 534442 14696 534448 14708
rect 534500 14696 534506 14748
rect 249426 14628 249432 14680
rect 249484 14668 249490 14680
rect 307846 14668 307852 14680
rect 249484 14640 307852 14668
rect 249484 14628 249490 14640
rect 307846 14628 307852 14640
rect 307904 14628 307910 14680
rect 319438 14628 319444 14680
rect 319496 14668 319502 14680
rect 538214 14668 538220 14680
rect 319496 14640 538220 14668
rect 319496 14628 319502 14640
rect 538214 14628 538220 14640
rect 538272 14628 538278 14680
rect 198734 14560 198740 14612
rect 198792 14600 198798 14612
rect 280798 14600 280804 14612
rect 198792 14572 280804 14600
rect 198792 14560 198798 14572
rect 280798 14560 280804 14572
rect 280856 14560 280862 14612
rect 318058 14560 318064 14612
rect 318116 14600 318122 14612
rect 541986 14600 541992 14612
rect 318116 14572 541992 14600
rect 318116 14560 318122 14572
rect 541986 14560 541992 14572
rect 542044 14560 542050 14612
rect 101950 14492 101956 14544
rect 102008 14532 102014 14544
rect 105630 14532 105636 14544
rect 102008 14504 105636 14532
rect 102008 14492 102014 14504
rect 105630 14492 105636 14504
rect 105688 14492 105694 14544
rect 167178 14492 167184 14544
rect 167236 14532 167242 14544
rect 290458 14532 290464 14544
rect 167236 14504 290464 14532
rect 167236 14492 167242 14504
rect 290458 14492 290464 14504
rect 290516 14492 290522 14544
rect 311802 14492 311808 14544
rect 311860 14532 311866 14544
rect 548610 14532 548616 14544
rect 311860 14504 548616 14532
rect 311860 14492 311866 14504
rect 548610 14492 548616 14504
rect 548668 14492 548674 14544
rect 66714 14424 66720 14476
rect 66772 14464 66778 14476
rect 113818 14464 113824 14476
rect 66772 14436 113824 14464
rect 66772 14424 66778 14436
rect 113818 14424 113824 14436
rect 113876 14424 113882 14476
rect 128170 14424 128176 14476
rect 128228 14464 128234 14476
rect 301498 14464 301504 14476
rect 128228 14436 301504 14464
rect 128228 14424 128234 14436
rect 301498 14424 301504 14436
rect 301556 14424 301562 14476
rect 307386 14424 307392 14476
rect 307444 14464 307450 14476
rect 559282 14464 559288 14476
rect 307444 14436 559288 14464
rect 307444 14424 307450 14436
rect 559282 14424 559288 14436
rect 559340 14424 559346 14476
rect 469858 13744 469864 13796
rect 469916 13784 469922 13796
rect 470686 13784 470692 13796
rect 469916 13756 470692 13784
rect 469916 13744 469922 13756
rect 470686 13744 470692 13756
rect 470744 13744 470750 13796
rect 248322 13472 248328 13524
rect 248380 13512 248386 13524
rect 312170 13512 312176 13524
rect 248380 13484 312176 13512
rect 248380 13472 248386 13484
rect 312170 13472 312176 13484
rect 312228 13472 312234 13524
rect 353570 13472 353576 13524
rect 353628 13512 353634 13524
rect 372706 13512 372712 13524
rect 353628 13484 372712 13512
rect 353628 13472 353634 13484
rect 372706 13472 372712 13484
rect 372764 13472 372770 13524
rect 246942 13404 246948 13456
rect 247000 13444 247006 13456
rect 316218 13444 316224 13456
rect 247000 13416 316224 13444
rect 247000 13404 247006 13416
rect 316218 13404 316224 13416
rect 316276 13404 316282 13456
rect 359458 13404 359464 13456
rect 359516 13444 359522 13456
rect 398926 13444 398932 13456
rect 359516 13416 398932 13444
rect 359516 13404 359522 13416
rect 398926 13404 398932 13416
rect 398984 13404 398990 13456
rect 245286 13336 245292 13388
rect 245344 13376 245350 13388
rect 319714 13376 319720 13388
rect 245344 13348 319720 13376
rect 245344 13336 245350 13348
rect 319714 13336 319720 13348
rect 319772 13336 319778 13388
rect 322106 13336 322112 13388
rect 322164 13376 322170 13388
rect 382458 13376 382464 13388
rect 322164 13348 382464 13376
rect 322164 13336 322170 13348
rect 382458 13336 382464 13348
rect 382516 13336 382522 13388
rect 311434 13268 311440 13320
rect 311492 13308 311498 13320
rect 385034 13308 385040 13320
rect 311492 13280 385040 13308
rect 311492 13268 311498 13280
rect 385034 13268 385040 13280
rect 385092 13268 385098 13320
rect 468478 13268 468484 13320
rect 468536 13308 468542 13320
rect 480530 13308 480536 13320
rect 468536 13280 480536 13308
rect 468536 13268 468542 13280
rect 480530 13268 480536 13280
rect 480588 13268 480594 13320
rect 245470 13200 245476 13252
rect 245528 13240 245534 13252
rect 322934 13240 322940 13252
rect 245528 13212 322940 13240
rect 245528 13200 245534 13212
rect 322934 13200 322940 13212
rect 322992 13200 322998 13252
rect 336274 13200 336280 13252
rect 336332 13240 336338 13252
rect 378410 13240 378416 13252
rect 336332 13212 378416 13240
rect 336332 13200 336338 13212
rect 378410 13200 378416 13212
rect 378468 13200 378474 13252
rect 402514 13200 402520 13252
rect 402572 13240 402578 13252
rect 489914 13240 489920 13252
rect 402572 13212 489920 13240
rect 402572 13200 402578 13212
rect 489914 13200 489920 13212
rect 489972 13200 489978 13252
rect 73062 13132 73068 13184
rect 73120 13172 73126 13184
rect 92474 13172 92480 13184
rect 73120 13144 92480 13172
rect 73120 13132 73126 13144
rect 92474 13132 92480 13144
rect 92532 13132 92538 13184
rect 94406 13132 94412 13184
rect 94464 13172 94470 13184
rect 105722 13172 105728 13184
rect 94464 13144 105728 13172
rect 94464 13132 94470 13144
rect 105722 13132 105728 13144
rect 105780 13132 105786 13184
rect 242802 13132 242808 13184
rect 242860 13172 242866 13184
rect 330386 13172 330392 13184
rect 242860 13144 330392 13172
rect 242860 13132 242866 13144
rect 330386 13132 330392 13144
rect 330444 13132 330450 13184
rect 341518 13132 341524 13184
rect 341576 13172 341582 13184
rect 459922 13172 459928 13184
rect 341576 13144 459928 13172
rect 341576 13132 341582 13144
rect 459922 13132 459928 13144
rect 459980 13132 459986 13184
rect 462958 13132 462964 13184
rect 463016 13172 463022 13184
rect 498286 13172 498292 13184
rect 463016 13144 498292 13172
rect 463016 13132 463022 13144
rect 498286 13132 498292 13144
rect 498344 13132 498350 13184
rect 60826 13064 60832 13116
rect 60884 13104 60890 13116
rect 82078 13104 82084 13116
rect 60884 13076 82084 13104
rect 60884 13064 60890 13076
rect 82078 13064 82084 13076
rect 82136 13064 82142 13116
rect 97442 13064 97448 13116
rect 97500 13104 97506 13116
rect 137278 13104 137284 13116
rect 97500 13076 137284 13104
rect 97500 13064 97506 13076
rect 137278 13064 137284 13076
rect 137336 13064 137342 13116
rect 156138 13064 156144 13116
rect 156196 13104 156202 13116
rect 293218 13104 293224 13116
rect 156196 13076 293224 13104
rect 156196 13064 156202 13076
rect 293218 13064 293224 13076
rect 293276 13064 293282 13116
rect 320450 13064 320456 13116
rect 320508 13104 320514 13116
rect 514846 13104 514852 13116
rect 320508 13076 514852 13104
rect 320508 13064 320514 13076
rect 514846 13064 514852 13076
rect 514904 13064 514910 13116
rect 465810 12928 465816 12980
rect 465868 12968 465874 12980
rect 471974 12968 471980 12980
rect 465868 12940 471980 12968
rect 465868 12928 465874 12940
rect 471974 12928 471980 12940
rect 472032 12928 472038 12980
rect 259362 12248 259368 12300
rect 259420 12288 259426 12300
rect 273254 12288 273260 12300
rect 259420 12260 273260 12288
rect 259420 12248 259426 12260
rect 273254 12248 273260 12260
rect 273312 12248 273318 12300
rect 257890 12180 257896 12232
rect 257948 12220 257954 12232
rect 276658 12220 276664 12232
rect 257948 12192 276664 12220
rect 257948 12180 257954 12192
rect 276658 12180 276664 12192
rect 276716 12180 276722 12232
rect 257706 12112 257712 12164
rect 257764 12152 257770 12164
rect 280706 12152 280712 12164
rect 257764 12124 280712 12152
rect 257764 12112 257770 12124
rect 280706 12112 280712 12124
rect 280764 12112 280770 12164
rect 255222 12044 255228 12096
rect 255280 12084 255286 12096
rect 287330 12084 287336 12096
rect 255280 12056 287336 12084
rect 255280 12044 255286 12056
rect 287330 12044 287336 12056
rect 287388 12044 287394 12096
rect 346946 12044 346952 12096
rect 347004 12084 347010 12096
rect 374270 12084 374276 12096
rect 347004 12056 374276 12084
rect 347004 12044 347010 12056
rect 374270 12044 374276 12056
rect 374328 12044 374334 12096
rect 253750 11976 253756 12028
rect 253808 12016 253814 12028
rect 291378 12016 291384 12028
rect 253808 11988 291384 12016
rect 253808 11976 253814 11988
rect 291378 11976 291384 11988
rect 291436 11976 291442 12028
rect 339494 11976 339500 12028
rect 339552 12016 339558 12028
rect 376846 12016 376852 12028
rect 339552 11988 376852 12016
rect 339552 11976 339558 11988
rect 376846 11976 376852 11988
rect 376904 11976 376910 12028
rect 253566 11908 253572 11960
rect 253624 11948 253630 11960
rect 294874 11948 294880 11960
rect 253624 11920 294880 11948
rect 253624 11908 253630 11920
rect 294874 11908 294880 11920
rect 294932 11908 294938 11960
rect 324406 11908 324412 11960
rect 324464 11948 324470 11960
rect 380986 11948 380992 11960
rect 324464 11920 380992 11948
rect 324464 11908 324470 11920
rect 380986 11908 380992 11920
rect 381044 11908 381050 11960
rect 455690 11908 455696 11960
rect 455748 11948 455754 11960
rect 474734 11948 474740 11960
rect 455748 11920 474740 11948
rect 455748 11908 455754 11920
rect 474734 11908 474740 11920
rect 474792 11908 474798 11960
rect 252462 11840 252468 11892
rect 252520 11880 252526 11892
rect 298094 11880 298100 11892
rect 252520 11852 298100 11880
rect 252520 11840 252526 11852
rect 298094 11840 298100 11852
rect 298152 11840 298158 11892
rect 314654 11840 314660 11892
rect 314712 11880 314718 11892
rect 383746 11880 383752 11892
rect 314712 11852 383752 11880
rect 314712 11840 314718 11852
rect 383746 11840 383752 11852
rect 383804 11840 383810 11892
rect 412634 11840 412640 11892
rect 412692 11880 412698 11892
rect 487246 11880 487252 11892
rect 412692 11852 487252 11880
rect 412692 11840 412698 11852
rect 487246 11840 487252 11852
rect 487304 11840 487310 11892
rect 71682 11772 71688 11824
rect 71740 11812 71746 11824
rect 99834 11812 99840 11824
rect 71740 11784 99840 11812
rect 71740 11772 71746 11784
rect 99834 11772 99840 11784
rect 99892 11772 99898 11824
rect 102042 11772 102048 11824
rect 102100 11812 102106 11824
rect 109034 11812 109040 11824
rect 102100 11784 109040 11812
rect 102100 11772 102106 11784
rect 109034 11772 109040 11784
rect 109092 11772 109098 11824
rect 256602 11772 256608 11824
rect 256660 11812 256666 11824
rect 284294 11812 284300 11824
rect 256660 11784 284300 11812
rect 256660 11772 256666 11784
rect 284294 11772 284300 11784
rect 284352 11772 284358 11824
rect 286594 11772 286600 11824
rect 286652 11812 286658 11824
rect 392026 11812 392032 11824
rect 286652 11784 392032 11812
rect 286652 11772 286658 11784
rect 392026 11772 392032 11784
rect 392084 11772 392090 11824
rect 405734 11772 405740 11824
rect 405792 11812 405798 11824
rect 490098 11812 490104 11824
rect 405792 11784 490104 11812
rect 405792 11772 405798 11784
rect 490098 11772 490104 11784
rect 490156 11772 490162 11824
rect 56778 11704 56784 11756
rect 56836 11744 56842 11756
rect 83458 11744 83464 11756
rect 56836 11716 83464 11744
rect 56836 11704 56842 11716
rect 83458 11704 83464 11716
rect 83516 11704 83522 11756
rect 89898 11704 89904 11756
rect 89956 11744 89962 11756
rect 140038 11744 140044 11756
rect 89956 11716 140044 11744
rect 89956 11704 89962 11716
rect 140038 11704 140044 11716
rect 140096 11704 140102 11756
rect 143534 11704 143540 11756
rect 143592 11744 143598 11756
rect 144730 11744 144736 11756
rect 143592 11716 144736 11744
rect 143592 11704 143598 11716
rect 144730 11704 144736 11716
rect 144788 11704 144794 11756
rect 297358 11744 297364 11756
rect 151786 11716 297364 11744
rect 142154 11636 142160 11688
rect 142212 11676 142218 11688
rect 151786 11676 151814 11716
rect 297358 11704 297364 11716
rect 297416 11704 297422 11756
rect 299474 11704 299480 11756
rect 299532 11744 299538 11756
rect 387886 11744 387892 11756
rect 299532 11716 387892 11744
rect 299532 11704 299538 11716
rect 387886 11704 387892 11716
rect 387944 11704 387950 11756
rect 390646 11704 390652 11756
rect 390704 11744 390710 11756
rect 494238 11744 494244 11756
rect 390704 11716 494244 11744
rect 390704 11704 390710 11716
rect 494238 11704 494244 11716
rect 494296 11704 494302 11756
rect 142212 11648 151814 11676
rect 142212 11636 142218 11648
rect 259454 11636 259460 11688
rect 259512 11676 259518 11688
rect 260650 11676 260656 11688
rect 259512 11648 260656 11676
rect 259512 11636 259518 11648
rect 260650 11636 260656 11648
rect 260708 11636 260714 11688
rect 259454 10956 259460 11008
rect 259512 10996 259518 11008
rect 262858 10996 262864 11008
rect 259512 10968 262864 10996
rect 259512 10956 259518 10968
rect 262858 10956 262864 10968
rect 262916 10956 262922 11008
rect 361114 10820 361120 10872
rect 361172 10860 361178 10872
rect 370130 10860 370136 10872
rect 361172 10832 370136 10860
rect 361172 10820 361178 10832
rect 370130 10820 370136 10832
rect 370188 10820 370194 10872
rect 245194 10684 245200 10736
rect 245252 10724 245258 10736
rect 266998 10724 267004 10736
rect 245252 10696 267004 10724
rect 245252 10684 245258 10696
rect 266998 10684 267004 10696
rect 267056 10684 267062 10736
rect 370130 10684 370136 10736
rect 370188 10724 370194 10736
rect 499666 10724 499672 10736
rect 370188 10696 499672 10724
rect 370188 10684 370194 10696
rect 499666 10684 499672 10696
rect 499724 10684 499730 10736
rect 237650 10616 237656 10668
rect 237708 10656 237714 10668
rect 269942 10656 269948 10668
rect 237708 10628 269948 10656
rect 237708 10616 237714 10628
rect 269942 10616 269948 10628
rect 270000 10616 270006 10668
rect 365806 10616 365812 10668
rect 365864 10656 365870 10668
rect 501046 10656 501052 10668
rect 365864 10628 501052 10656
rect 365864 10616 365870 10628
rect 501046 10616 501052 10628
rect 501104 10616 501110 10668
rect 234614 10548 234620 10600
rect 234672 10588 234678 10600
rect 269758 10588 269764 10600
rect 234672 10560 269764 10588
rect 234672 10548 234678 10560
rect 269758 10548 269764 10560
rect 269816 10548 269822 10600
rect 363506 10548 363512 10600
rect 363564 10588 363570 10600
rect 502518 10588 502524 10600
rect 363564 10560 502524 10588
rect 363564 10548 363570 10560
rect 502518 10548 502524 10560
rect 502576 10548 502582 10600
rect 226334 10480 226340 10532
rect 226392 10520 226398 10532
rect 272518 10520 272524 10532
rect 226392 10492 272524 10520
rect 226392 10480 226398 10492
rect 272518 10480 272524 10492
rect 272576 10480 272582 10532
rect 359458 10480 359464 10532
rect 359516 10520 359522 10532
rect 502702 10520 502708 10532
rect 359516 10492 502708 10520
rect 359516 10480 359522 10492
rect 502702 10480 502708 10492
rect 502760 10480 502766 10532
rect 235902 10412 235908 10464
rect 235960 10452 235966 10464
rect 355226 10452 355232 10464
rect 235960 10424 355232 10452
rect 235960 10412 235966 10424
rect 355226 10412 355232 10424
rect 355284 10412 355290 10464
rect 356330 10412 356336 10464
rect 356388 10452 356394 10464
rect 503806 10452 503812 10464
rect 356388 10424 503812 10452
rect 356388 10412 356394 10424
rect 503806 10412 503812 10424
rect 503864 10412 503870 10464
rect 91554 10344 91560 10396
rect 91612 10384 91618 10396
rect 105538 10384 105544 10396
rect 91612 10356 105544 10384
rect 91612 10344 91618 10356
rect 105538 10344 105544 10356
rect 105596 10344 105602 10396
rect 223574 10344 223580 10396
rect 223632 10384 223638 10396
rect 274082 10384 274088 10396
rect 223632 10356 274088 10384
rect 223632 10344 223638 10356
rect 274082 10344 274088 10356
rect 274140 10344 274146 10396
rect 352834 10344 352840 10396
rect 352892 10384 352898 10396
rect 505186 10384 505192 10396
rect 352892 10356 505192 10384
rect 352892 10344 352898 10356
rect 505186 10344 505192 10356
rect 505244 10344 505250 10396
rect 65058 10276 65064 10328
rect 65116 10316 65122 10328
rect 146938 10316 146944 10328
rect 65116 10288 146944 10316
rect 65116 10276 65122 10288
rect 146938 10276 146944 10288
rect 146996 10276 147002 10328
rect 219986 10276 219992 10328
rect 220044 10316 220050 10328
rect 273898 10316 273904 10328
rect 220044 10288 273904 10316
rect 220044 10276 220050 10288
rect 273898 10276 273904 10288
rect 273956 10276 273962 10328
rect 340966 10276 340972 10328
rect 341024 10316 341030 10328
rect 507854 10316 507860 10328
rect 341024 10288 507860 10316
rect 341024 10276 341030 10288
rect 507854 10276 507860 10288
rect 507912 10276 507918 10328
rect 77018 9596 77024 9648
rect 77076 9636 77082 9648
rect 78582 9636 78588 9648
rect 77076 9608 78588 9636
rect 77076 9596 77082 9608
rect 78582 9596 78588 9608
rect 78640 9596 78646 9648
rect 151722 9596 151728 9648
rect 151780 9636 151786 9648
rect 153010 9636 153016 9648
rect 151780 9608 153016 9636
rect 151780 9596 151786 9608
rect 153010 9596 153016 9608
rect 153068 9596 153074 9648
rect 255866 9460 255872 9512
rect 255924 9500 255930 9512
rect 264238 9500 264244 9512
rect 255924 9472 264244 9500
rect 255924 9460 255930 9472
rect 264238 9460 264244 9472
rect 264296 9460 264302 9512
rect 241698 9392 241704 9444
rect 241756 9432 241762 9444
rect 268378 9432 268384 9444
rect 241756 9404 268384 9432
rect 241756 9392 241762 9404
rect 268378 9392 268384 9404
rect 268436 9392 268442 9444
rect 231026 9324 231032 9376
rect 231084 9364 231090 9376
rect 271138 9364 271144 9376
rect 231084 9336 271144 9364
rect 231084 9324 231090 9336
rect 271138 9324 271144 9336
rect 271196 9324 271202 9376
rect 310238 9324 310244 9376
rect 310296 9364 310302 9376
rect 517606 9364 517612 9376
rect 310296 9336 517612 9364
rect 310296 9324 310302 9336
rect 517606 9324 517612 9336
rect 517664 9324 517670 9376
rect 216858 9256 216864 9308
rect 216916 9296 216922 9308
rect 275278 9296 275284 9308
rect 216916 9268 275284 9296
rect 216916 9256 216922 9268
rect 275278 9256 275284 9268
rect 275336 9256 275342 9308
rect 306742 9256 306748 9308
rect 306800 9296 306806 9308
rect 518986 9296 518992 9308
rect 306800 9268 518992 9296
rect 306800 9256 306806 9268
rect 518986 9256 518992 9268
rect 519044 9256 519050 9308
rect 181438 9188 181444 9240
rect 181496 9228 181502 9240
rect 286502 9228 286508 9240
rect 181496 9200 286508 9228
rect 181496 9188 181502 9200
rect 286502 9188 286508 9200
rect 286560 9188 286566 9240
rect 303154 9188 303160 9240
rect 303212 9228 303218 9240
rect 519170 9228 519176 9240
rect 303212 9200 519176 9228
rect 303212 9188 303218 9200
rect 519170 9188 519176 9200
rect 519228 9188 519234 9240
rect 177850 9120 177856 9172
rect 177908 9160 177914 9172
rect 286318 9160 286324 9172
rect 177908 9132 286324 9160
rect 177908 9120 177914 9132
rect 286318 9120 286324 9132
rect 286376 9120 286382 9172
rect 299658 9120 299664 9172
rect 299716 9160 299722 9172
rect 520366 9160 520372 9172
rect 299716 9132 520372 9160
rect 299716 9120 299722 9132
rect 520366 9120 520372 9132
rect 520424 9120 520430 9172
rect 174262 9052 174268 9104
rect 174320 9092 174326 9104
rect 287698 9092 287704 9104
rect 174320 9064 287704 9092
rect 174320 9052 174326 9064
rect 287698 9052 287704 9064
rect 287756 9052 287762 9104
rect 296070 9052 296076 9104
rect 296128 9092 296134 9104
rect 521746 9092 521752 9104
rect 296128 9064 521752 9092
rect 296128 9052 296134 9064
rect 521746 9052 521752 9064
rect 521804 9052 521810 9104
rect 84470 8984 84476 9036
rect 84528 9024 84534 9036
rect 108298 9024 108304 9036
rect 84528 8996 108304 9024
rect 84528 8984 84534 8996
rect 108298 8984 108304 8996
rect 108356 8984 108362 9036
rect 192018 8984 192024 9036
rect 192076 9024 192082 9036
rect 282178 9024 282184 9036
rect 192076 8996 282184 9024
rect 192076 8984 192082 8996
rect 282178 8984 282184 8996
rect 282236 8984 282242 9036
rect 285398 8984 285404 9036
rect 285456 9024 285462 9036
rect 524506 9024 524512 9036
rect 285456 8996 524512 9024
rect 285456 8984 285462 8996
rect 524506 8984 524512 8996
rect 524564 8984 524570 9036
rect 62022 8916 62028 8968
rect 62080 8956 62086 8968
rect 148318 8956 148324 8968
rect 62080 8928 148324 8956
rect 62080 8916 62086 8928
rect 148318 8916 148324 8928
rect 148376 8916 148382 8968
rect 206186 8916 206192 8968
rect 206244 8956 206250 8968
rect 278038 8956 278044 8968
rect 206244 8928 278044 8956
rect 206244 8916 206250 8928
rect 278038 8916 278044 8928
rect 278096 8916 278102 8968
rect 281902 8916 281908 8968
rect 281960 8956 281966 8968
rect 525794 8956 525800 8968
rect 281960 8928 525800 8956
rect 281960 8916 281966 8928
rect 525794 8916 525800 8928
rect 525852 8916 525858 8968
rect 249978 7964 249984 8016
rect 250036 8004 250042 8016
rect 535638 8004 535644 8016
rect 250036 7976 535644 8004
rect 250036 7964 250042 7976
rect 535638 7964 535644 7976
rect 535696 7964 535702 8016
rect 246390 7896 246396 7948
rect 246448 7936 246454 7948
rect 535822 7936 535828 7948
rect 246448 7908 535828 7936
rect 246448 7896 246454 7908
rect 535822 7896 535828 7908
rect 535880 7896 535886 7948
rect 45462 7828 45468 7880
rect 45520 7868 45526 7880
rect 119338 7868 119344 7880
rect 45520 7840 119344 7868
rect 45520 7828 45526 7840
rect 119338 7828 119344 7840
rect 119396 7828 119402 7880
rect 239306 7828 239312 7880
rect 239364 7868 239370 7880
rect 538306 7868 538312 7880
rect 239364 7840 538312 7868
rect 239364 7828 239370 7840
rect 538306 7828 538312 7840
rect 538364 7828 538370 7880
rect 38378 7760 38384 7812
rect 38436 7800 38442 7812
rect 120718 7800 120724 7812
rect 38436 7772 120724 7800
rect 38436 7760 38442 7772
rect 120718 7760 120724 7772
rect 120776 7760 120782 7812
rect 235810 7760 235816 7812
rect 235868 7800 235874 7812
rect 539778 7800 539784 7812
rect 235868 7772 539784 7800
rect 235868 7760 235874 7772
rect 539778 7760 539784 7772
rect 539836 7760 539842 7812
rect 31294 7692 31300 7744
rect 31352 7732 31358 7744
rect 123478 7732 123484 7744
rect 31352 7704 123484 7732
rect 31352 7692 31358 7704
rect 123478 7692 123484 7704
rect 123536 7692 123542 7744
rect 232222 7692 232228 7744
rect 232280 7732 232286 7744
rect 539594 7732 539600 7744
rect 232280 7704 539600 7732
rect 232280 7692 232286 7704
rect 539594 7692 539600 7704
rect 539652 7692 539658 7744
rect 23014 7624 23020 7676
rect 23072 7664 23078 7676
rect 124858 7664 124864 7676
rect 23072 7636 124864 7664
rect 23072 7624 23078 7636
rect 124858 7624 124864 7636
rect 124916 7624 124922 7676
rect 228726 7624 228732 7676
rect 228784 7664 228790 7676
rect 541066 7664 541072 7676
rect 228784 7636 541072 7664
rect 228784 7624 228790 7636
rect 541066 7624 541072 7636
rect 541124 7624 541130 7676
rect 13538 7556 13544 7608
rect 13596 7596 13602 7608
rect 127618 7596 127624 7608
rect 13596 7568 127624 7596
rect 13596 7556 13602 7568
rect 127618 7556 127624 7568
rect 127676 7556 127682 7608
rect 132954 7556 132960 7608
rect 133012 7596 133018 7608
rect 568850 7596 568856 7608
rect 133012 7568 568856 7596
rect 133012 7556 133018 7568
rect 568850 7556 568856 7568
rect 568908 7556 568914 7608
rect 523034 7488 523040 7540
rect 523092 7528 523098 7540
rect 523862 7528 523868 7540
rect 523092 7500 523868 7528
rect 523092 7488 523098 7500
rect 523862 7488 523868 7500
rect 523920 7488 523926 7540
rect 247586 6536 247592 6588
rect 247644 6576 247650 6588
rect 403158 6576 403164 6588
rect 247644 6548 403164 6576
rect 247644 6536 247650 6548
rect 403158 6536 403164 6548
rect 403216 6536 403222 6588
rect 75822 6468 75828 6520
rect 75880 6508 75886 6520
rect 85666 6508 85672 6520
rect 75880 6480 85672 6508
rect 75880 6468 75886 6480
rect 85666 6468 85672 6480
rect 85724 6468 85730 6520
rect 244090 6468 244096 6520
rect 244148 6508 244154 6520
rect 404446 6508 404452 6520
rect 244148 6480 404452 6508
rect 244148 6468 244154 6480
rect 404446 6468 404452 6480
rect 404504 6468 404510 6520
rect 70302 6400 70308 6452
rect 70360 6440 70366 6452
rect 112438 6440 112444 6452
rect 70360 6412 112444 6440
rect 70360 6400 70366 6412
rect 112438 6400 112444 6412
rect 112496 6400 112502 6452
rect 240502 6400 240508 6452
rect 240560 6440 240566 6452
rect 405826 6440 405832 6452
rect 240560 6412 405832 6440
rect 240560 6400 240566 6412
rect 405826 6400 405832 6412
rect 405884 6400 405890 6452
rect 59630 6332 59636 6384
rect 59688 6372 59694 6384
rect 115198 6372 115204 6384
rect 59688 6344 115204 6372
rect 59688 6332 59694 6344
rect 115198 6332 115204 6344
rect 115256 6332 115262 6384
rect 229830 6332 229836 6384
rect 229888 6372 229894 6384
rect 408586 6372 408592 6384
rect 229888 6344 408592 6372
rect 229888 6332 229894 6344
rect 408586 6332 408592 6344
rect 408644 6332 408650 6384
rect 416682 6332 416688 6384
rect 416740 6372 416746 6384
rect 486142 6372 486148 6384
rect 416740 6344 486148 6372
rect 416740 6332 416746 6344
rect 486142 6332 486148 6344
rect 486200 6332 486206 6384
rect 56042 6264 56048 6316
rect 56100 6304 56106 6316
rect 116578 6304 116584 6316
rect 56100 6276 116584 6304
rect 56100 6264 56106 6276
rect 116578 6264 116584 6276
rect 116636 6264 116642 6316
rect 226426 6264 226432 6316
rect 226484 6304 226490 6316
rect 409966 6304 409972 6316
rect 226484 6276 409972 6304
rect 226484 6264 226490 6276
rect 409966 6264 409972 6276
rect 410024 6264 410030 6316
rect 442258 6264 442264 6316
rect 442316 6304 442322 6316
rect 569126 6304 569132 6316
rect 442316 6276 569132 6304
rect 442316 6264 442322 6276
rect 569126 6264 569132 6276
rect 569184 6264 569190 6316
rect 14734 6196 14740 6248
rect 14792 6236 14798 6248
rect 94498 6236 94504 6248
rect 14792 6208 94504 6236
rect 14792 6196 14798 6208
rect 94498 6196 94504 6208
rect 94556 6196 94562 6248
rect 222746 6196 222752 6248
rect 222804 6236 222810 6248
rect 411622 6236 411628 6248
rect 222804 6208 411628 6236
rect 222804 6196 222810 6208
rect 411622 6196 411628 6208
rect 411680 6196 411686 6248
rect 441062 6196 441068 6248
rect 441120 6236 441126 6248
rect 572714 6236 572720 6248
rect 441120 6208 572720 6236
rect 441120 6196 441126 6208
rect 572714 6196 572720 6208
rect 572772 6196 572778 6248
rect 8754 6128 8760 6180
rect 8812 6168 8818 6180
rect 129182 6168 129188 6180
rect 8812 6140 129188 6168
rect 8812 6128 8818 6140
rect 129182 6128 129188 6140
rect 129240 6128 129246 6180
rect 219250 6128 219256 6180
rect 219308 6168 219314 6180
rect 411438 6168 411444 6180
rect 219308 6140 411444 6168
rect 219308 6128 219314 6140
rect 411438 6128 411444 6140
rect 411496 6128 411502 6180
rect 440878 6128 440884 6180
rect 440936 6168 440942 6180
rect 576302 6168 576308 6180
rect 440936 6140 576308 6168
rect 440936 6128 440942 6140
rect 576302 6128 576308 6140
rect 576360 6128 576366 6180
rect 77202 5516 77208 5568
rect 77260 5556 77266 5568
rect 82078 5556 82084 5568
rect 77260 5528 82084 5556
rect 77260 5516 77266 5528
rect 82078 5516 82084 5528
rect 82136 5516 82142 5568
rect 86862 5244 86868 5296
rect 86920 5284 86926 5296
rect 141418 5284 141424 5296
rect 86920 5256 141424 5284
rect 86920 5244 86926 5256
rect 141418 5244 141424 5256
rect 141476 5244 141482 5296
rect 71498 5176 71504 5228
rect 71556 5216 71562 5228
rect 79318 5216 79324 5228
rect 71556 5188 79324 5216
rect 71556 5176 71562 5188
rect 79318 5176 79324 5188
rect 79376 5176 79382 5228
rect 83274 5176 83280 5228
rect 83332 5216 83338 5228
rect 141602 5216 141608 5228
rect 83332 5188 141608 5216
rect 83332 5176 83338 5188
rect 141602 5176 141608 5188
rect 141660 5176 141666 5228
rect 460198 5176 460204 5228
rect 460256 5216 460262 5228
rect 508866 5216 508872 5228
rect 460256 5188 508872 5216
rect 460256 5176 460262 5188
rect 508866 5176 508872 5188
rect 508924 5176 508930 5228
rect 79686 5108 79692 5160
rect 79744 5148 79750 5160
rect 142798 5148 142804 5160
rect 79744 5120 142804 5148
rect 79744 5108 79750 5120
rect 142798 5108 142804 5120
rect 142856 5108 142862 5160
rect 458818 5108 458824 5160
rect 458876 5148 458882 5160
rect 512454 5148 512460 5160
rect 458876 5120 512460 5148
rect 458876 5108 458882 5120
rect 512454 5108 512460 5120
rect 512512 5108 512518 5160
rect 76190 5040 76196 5092
rect 76248 5080 76254 5092
rect 144178 5080 144184 5092
rect 76248 5052 144184 5080
rect 76248 5040 76254 5052
rect 144178 5040 144184 5052
rect 144236 5040 144242 5092
rect 197906 5040 197912 5092
rect 197964 5080 197970 5092
rect 197964 5052 200114 5080
rect 197964 5040 197970 5052
rect 72602 4972 72608 5024
rect 72660 5012 72666 5024
rect 145558 5012 145564 5024
rect 72660 4984 145564 5012
rect 72660 4972 72666 4984
rect 145558 4972 145564 4984
rect 145616 4972 145622 5024
rect 69106 4904 69112 4956
rect 69164 4944 69170 4956
rect 145742 4944 145748 4956
rect 69164 4916 145748 4944
rect 69164 4904 69170 4916
rect 145742 4904 145748 4916
rect 145800 4904 145806 4956
rect 200086 4944 200114 5052
rect 212166 5040 212172 5092
rect 212224 5080 212230 5092
rect 414106 5080 414112 5092
rect 212224 5052 414112 5080
rect 212224 5040 212230 5052
rect 414106 5040 414112 5052
rect 414164 5040 414170 5092
rect 457438 5040 457444 5092
rect 457496 5080 457502 5092
rect 515950 5080 515956 5092
rect 457496 5052 515956 5080
rect 457496 5040 457502 5052
rect 515950 5040 515956 5052
rect 516008 5040 516014 5092
rect 201586 4972 201592 5024
rect 201644 5012 201650 5024
rect 416866 5012 416872 5024
rect 201644 4984 416872 5012
rect 201644 4972 201650 4984
rect 416866 4972 416872 4984
rect 416924 4972 416930 5024
rect 457622 4972 457628 5024
rect 457680 5012 457686 5024
rect 519538 5012 519544 5024
rect 457680 4984 519544 5012
rect 457680 4972 457686 4984
rect 519538 4972 519544 4984
rect 519596 4972 519602 5024
rect 418246 4944 418252 4956
rect 200086 4916 418252 4944
rect 418246 4904 418252 4916
rect 418304 4904 418310 4956
rect 454678 4904 454684 4956
rect 454736 4944 454742 4956
rect 526622 4944 526628 4956
rect 454736 4916 526628 4944
rect 454736 4904 454742 4916
rect 526622 4904 526628 4916
rect 526680 4904 526686 4956
rect 4062 4836 4068 4888
rect 4120 4876 4126 4888
rect 128998 4876 129004 4888
rect 4120 4848 129004 4876
rect 4120 4836 4126 4848
rect 128998 4836 129004 4848
rect 129056 4836 129062 4888
rect 187326 4836 187332 4888
rect 187384 4876 187390 4888
rect 421006 4876 421012 4888
rect 187384 4848 421012 4876
rect 187384 4836 187390 4848
rect 421006 4836 421012 4848
rect 421064 4836 421070 4888
rect 453390 4836 453396 4888
rect 453448 4876 453454 4888
rect 516778 4876 516784 4888
rect 453448 4848 516784 4876
rect 453448 4836 453454 4848
rect 516778 4836 516784 4848
rect 516836 4836 516842 4888
rect 516888 4848 521654 4876
rect 12342 4768 12348 4820
rect 12400 4808 12406 4820
rect 162118 4808 162124 4820
rect 12400 4780 162124 4808
rect 12400 4768 12406 4780
rect 162118 4768 162124 4780
rect 162176 4768 162182 4820
rect 183738 4768 183744 4820
rect 183796 4808 183802 4820
rect 422386 4808 422392 4820
rect 183796 4780 422392 4808
rect 183796 4768 183802 4780
rect 422386 4768 422392 4780
rect 422444 4768 422450 4820
rect 453482 4768 453488 4820
rect 453540 4808 453546 4820
rect 516888 4808 516916 4848
rect 453540 4780 516916 4808
rect 521626 4808 521654 4848
rect 533706 4808 533712 4820
rect 521626 4780 533712 4808
rect 453540 4768 453546 4780
rect 533706 4768 533712 4780
rect 533764 4768 533770 4820
rect 516778 4700 516784 4752
rect 516836 4740 516842 4752
rect 530118 4740 530124 4752
rect 516836 4712 530124 4740
rect 516836 4700 516842 4712
rect 530118 4700 530124 4712
rect 530176 4700 530182 4752
rect 74994 4156 75000 4208
rect 75052 4196 75058 4208
rect 77938 4196 77944 4208
rect 75052 4168 77944 4196
rect 75052 4156 75058 4168
rect 77938 4156 77944 4168
rect 77996 4156 78002 4208
rect 209774 4156 209780 4208
rect 209832 4196 209838 4208
rect 210970 4196 210976 4208
rect 209832 4168 210976 4196
rect 209832 4156 209838 4168
rect 210970 4156 210976 4168
rect 211028 4156 211034 4208
rect 251174 4156 251180 4208
rect 251232 4196 251238 4208
rect 252370 4196 252376 4208
rect 251232 4168 252376 4196
rect 251232 4156 251238 4168
rect 252370 4156 252376 4168
rect 252428 4156 252434 4208
rect 267734 4156 267740 4208
rect 267792 4196 267798 4208
rect 268470 4196 268476 4208
rect 267792 4168 268476 4196
rect 267792 4156 267798 4168
rect 268470 4156 268476 4168
rect 268528 4156 268534 4208
rect 292574 4156 292580 4208
rect 292632 4196 292638 4208
rect 293310 4196 293316 4208
rect 292632 4168 293316 4196
rect 292632 4156 292638 4168
rect 293310 4156 293316 4168
rect 293368 4156 293374 4208
rect 307846 4156 307852 4208
rect 307904 4196 307910 4208
rect 309042 4196 309048 4208
rect 307904 4168 309048 4196
rect 307904 4156 307910 4168
rect 309042 4156 309048 4168
rect 309100 4156 309106 4208
rect 68646 4088 68652 4140
rect 68704 4128 68710 4140
rect 110506 4128 110512 4140
rect 68704 4100 110512 4128
rect 68704 4088 68710 4100
rect 110506 4088 110512 4100
rect 110564 4088 110570 4140
rect 208026 4088 208032 4140
rect 208084 4128 208090 4140
rect 450906 4128 450912 4140
rect 208084 4100 450912 4128
rect 208084 4088 208090 4100
rect 450906 4088 450912 4100
rect 450964 4088 450970 4140
rect 566458 4088 566464 4140
rect 566516 4128 566522 4140
rect 568022 4128 568028 4140
rect 566516 4100 568028 4128
rect 566516 4088 566522 4100
rect 568022 4088 568028 4100
rect 568080 4088 568086 4140
rect 576118 4088 576124 4140
rect 576176 4128 576182 4140
rect 577406 4128 577412 4140
rect 576176 4100 577412 4128
rect 576176 4088 576182 4100
rect 577406 4088 577412 4100
rect 577464 4088 577470 4140
rect 43070 4020 43076 4072
rect 43128 4060 43134 4072
rect 87598 4060 87604 4072
rect 43128 4032 87604 4060
rect 43128 4020 43134 4032
rect 87598 4020 87604 4032
rect 87656 4020 87662 4072
rect 206922 4020 206928 4072
rect 206980 4060 206986 4072
rect 454494 4060 454500 4072
rect 206980 4032 454500 4060
rect 206980 4020 206986 4032
rect 454494 4020 454500 4032
rect 454552 4020 454558 4072
rect 67542 3952 67548 4004
rect 67600 3992 67606 4004
rect 114002 3992 114008 4004
rect 67600 3964 114008 3992
rect 67600 3952 67606 3964
rect 114002 3952 114008 3964
rect 114060 3952 114066 4004
rect 205542 3952 205548 4004
rect 205600 3992 205606 4004
rect 458082 3992 458088 4004
rect 205600 3964 458088 3992
rect 205600 3952 205606 3964
rect 458082 3952 458088 3964
rect 458140 3952 458146 4004
rect 547138 3952 547144 4004
rect 547196 3992 547202 4004
rect 550266 3992 550272 4004
rect 547196 3964 550272 3992
rect 547196 3952 547202 3964
rect 550266 3952 550272 3964
rect 550324 3952 550330 4004
rect 39574 3884 39580 3936
rect 39632 3924 39638 3936
rect 88978 3924 88984 3936
rect 39632 3896 88984 3924
rect 39632 3884 39638 3896
rect 88978 3884 88984 3896
rect 89036 3884 89042 3936
rect 203886 3884 203892 3936
rect 203944 3924 203950 3936
rect 461578 3924 461584 3936
rect 203944 3896 461584 3924
rect 203944 3884 203950 3896
rect 461578 3884 461584 3896
rect 461636 3884 461642 3936
rect 66162 3816 66168 3868
rect 66220 3856 66226 3868
rect 117590 3856 117596 3868
rect 66220 3828 117596 3856
rect 66220 3816 66226 3828
rect 117590 3816 117596 3828
rect 117648 3816 117654 3868
rect 204070 3816 204076 3868
rect 204128 3856 204134 3868
rect 465166 3856 465172 3868
rect 204128 3828 465172 3856
rect 204128 3816 204134 3828
rect 465166 3816 465172 3828
rect 465224 3816 465230 3868
rect 35986 3748 35992 3800
rect 36044 3788 36050 3800
rect 89254 3788 89260 3800
rect 36044 3760 89260 3788
rect 36044 3748 36050 3760
rect 89254 3748 89260 3760
rect 89312 3748 89318 3800
rect 100662 3748 100668 3800
rect 100720 3788 100726 3800
rect 112806 3788 112812 3800
rect 100720 3760 112812 3788
rect 100720 3748 100726 3760
rect 112806 3748 112812 3760
rect 112864 3748 112870 3800
rect 202782 3748 202788 3800
rect 202840 3788 202846 3800
rect 468662 3788 468668 3800
rect 202840 3760 468668 3788
rect 202840 3748 202846 3760
rect 468662 3748 468668 3760
rect 468720 3748 468726 3800
rect 15930 3680 15936 3732
rect 15988 3720 15994 3732
rect 61378 3720 61384 3732
rect 15988 3692 61384 3720
rect 15988 3680 15994 3692
rect 61378 3680 61384 3692
rect 61436 3680 61442 3732
rect 64690 3680 64696 3732
rect 64748 3720 64754 3732
rect 121086 3720 121092 3732
rect 64748 3692 121092 3720
rect 64748 3680 64754 3692
rect 121086 3680 121092 3692
rect 121144 3680 121150 3732
rect 201402 3680 201408 3732
rect 201460 3720 201466 3732
rect 472250 3720 472256 3732
rect 201460 3692 472256 3720
rect 201460 3680 201466 3692
rect 472250 3680 472256 3692
rect 472308 3680 472314 3732
rect 32398 3612 32404 3664
rect 32456 3652 32462 3664
rect 90358 3652 90364 3664
rect 32456 3624 90364 3652
rect 32456 3612 32462 3624
rect 90358 3612 90364 3624
rect 90416 3612 90422 3664
rect 99282 3612 99288 3664
rect 99340 3652 99346 3664
rect 116394 3652 116400 3664
rect 99340 3624 116400 3652
rect 99340 3612 99346 3624
rect 116394 3612 116400 3624
rect 116452 3612 116458 3664
rect 118786 3612 118792 3664
rect 118844 3652 118850 3664
rect 131758 3652 131764 3664
rect 118844 3624 131764 3652
rect 118844 3612 118850 3624
rect 131758 3612 131764 3624
rect 131816 3612 131822 3664
rect 168282 3612 168288 3664
rect 168340 3652 168346 3664
rect 168340 3624 171134 3652
rect 168340 3612 168346 3624
rect 11146 3544 11152 3596
rect 11204 3584 11210 3596
rect 62758 3584 62764 3596
rect 11204 3556 62764 3584
rect 11204 3544 11210 3556
rect 62758 3544 62764 3556
rect 62816 3544 62822 3596
rect 64506 3544 64512 3596
rect 64564 3584 64570 3596
rect 124674 3584 124680 3596
rect 64564 3556 124680 3584
rect 64564 3544 64570 3556
rect 124674 3544 124680 3556
rect 124732 3544 124738 3596
rect 130378 3544 130384 3596
rect 130436 3544 130442 3596
rect 135254 3544 135260 3596
rect 135312 3584 135318 3596
rect 136450 3584 136456 3596
rect 135312 3556 136456 3584
rect 135312 3544 135318 3556
rect 136450 3544 136456 3556
rect 136508 3544 136514 3596
rect 168374 3544 168380 3596
rect 168432 3584 168438 3596
rect 169570 3584 169576 3596
rect 168432 3556 169576 3584
rect 168432 3544 168438 3556
rect 169570 3544 169576 3556
rect 169628 3544 169634 3596
rect 171106 3584 171134 3624
rect 193214 3612 193220 3664
rect 193272 3652 193278 3664
rect 194410 3652 194416 3664
rect 193272 3624 194416 3652
rect 193272 3612 193278 3624
rect 194410 3612 194416 3624
rect 194468 3612 194474 3664
rect 199746 3612 199752 3664
rect 199804 3652 199810 3664
rect 475746 3652 475752 3664
rect 199804 3624 475752 3652
rect 199804 3612 199810 3624
rect 475746 3612 475752 3624
rect 475804 3612 475810 3664
rect 580994 3584 581000 3596
rect 171106 3556 581000 3584
rect 580994 3544 581000 3556
rect 581052 3544 581058 3596
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 10318 3516 10324 3528
rect 7708 3488 10324 3516
rect 7708 3476 7714 3488
rect 10318 3476 10324 3488
rect 10376 3476 10382 3528
rect 28902 3476 28908 3528
rect 28960 3516 28966 3528
rect 91738 3516 91744 3528
rect 28960 3488 91744 3516
rect 28960 3476 28966 3488
rect 91738 3476 91744 3488
rect 91796 3476 91802 3528
rect 97810 3476 97816 3528
rect 97868 3516 97874 3528
rect 119890 3516 119896 3528
rect 97868 3488 119896 3516
rect 97868 3476 97874 3488
rect 119890 3476 119896 3488
rect 119948 3476 119954 3528
rect 122282 3476 122288 3528
rect 122340 3516 122346 3528
rect 130396 3516 130424 3544
rect 122340 3488 130424 3516
rect 122340 3476 122346 3488
rect 160094 3476 160100 3528
rect 160152 3516 160158 3528
rect 161290 3516 161296 3528
rect 160152 3488 161296 3516
rect 160152 3476 160158 3488
rect 161290 3476 161296 3488
rect 161348 3476 161354 3528
rect 199930 3476 199936 3528
rect 199988 3516 199994 3528
rect 479334 3516 479340 3528
rect 199988 3488 479340 3516
rect 199988 3476 199994 3488
rect 479334 3476 479340 3488
rect 479392 3476 479398 3528
rect 498194 3476 498200 3528
rect 498252 3516 498258 3528
rect 499022 3516 499028 3528
rect 498252 3488 499028 3516
rect 498252 3476 498258 3488
rect 499022 3476 499028 3488
rect 499080 3476 499086 3528
rect 538858 3476 538864 3528
rect 538916 3516 538922 3528
rect 539594 3516 539600 3528
rect 538916 3488 539600 3516
rect 538916 3476 538922 3488
rect 539594 3476 539600 3488
rect 539652 3476 539658 3528
rect 564434 3476 564440 3528
rect 564492 3516 564498 3528
rect 565262 3516 565268 3528
rect 564492 3488 565268 3516
rect 564492 3476 564498 3488
rect 565262 3476 565268 3488
rect 565320 3476 565326 3528
rect 24210 3408 24216 3460
rect 24268 3448 24274 3460
rect 93302 3448 93308 3460
rect 24268 3420 93308 3448
rect 24268 3408 24274 3420
rect 93302 3408 93308 3420
rect 93360 3408 93366 3460
rect 97626 3408 97632 3460
rect 97684 3448 97690 3460
rect 123478 3448 123484 3460
rect 97684 3420 123484 3448
rect 97684 3408 97690 3420
rect 123478 3408 123484 3420
rect 123536 3408 123542 3460
rect 166626 3408 166632 3460
rect 166684 3448 166690 3460
rect 582190 3448 582196 3460
rect 166684 3420 582196 3448
rect 166684 3408 166690 3420
rect 582190 3408 582196 3420
rect 582248 3408 582254 3460
rect 46658 3340 46664 3392
rect 46716 3380 46722 3392
rect 86218 3380 86224 3392
rect 46716 3352 86224 3380
rect 46716 3340 46722 3352
rect 86218 3340 86224 3352
rect 86276 3340 86282 3392
rect 201494 3340 201500 3392
rect 201552 3380 201558 3392
rect 202690 3380 202696 3392
rect 201552 3352 202696 3380
rect 201552 3340 201558 3352
rect 202690 3340 202696 3352
rect 202748 3340 202754 3392
rect 208210 3340 208216 3392
rect 208268 3380 208274 3392
rect 447410 3380 447416 3392
rect 208268 3352 447416 3380
rect 208268 3340 208274 3352
rect 447410 3340 447416 3352
rect 447468 3340 447474 3392
rect 448606 3340 448612 3392
rect 448664 3380 448670 3392
rect 449802 3380 449808 3392
rect 448664 3352 449808 3380
rect 448664 3340 448670 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 2866 3272 2872 3324
rect 2924 3312 2930 3324
rect 7558 3312 7564 3324
rect 2924 3284 7564 3312
rect 2924 3272 2930 3284
rect 7558 3272 7564 3284
rect 7616 3272 7622 3324
rect 68830 3272 68836 3324
rect 68888 3312 68894 3324
rect 106918 3312 106924 3324
rect 68888 3284 106924 3312
rect 68888 3272 68894 3284
rect 106918 3272 106924 3284
rect 106976 3272 106982 3324
rect 209682 3272 209688 3324
rect 209740 3312 209746 3324
rect 443822 3312 443828 3324
rect 209740 3284 443828 3312
rect 209740 3272 209746 3284
rect 443822 3272 443828 3284
rect 443880 3272 443886 3324
rect 70210 3204 70216 3256
rect 70268 3244 70274 3256
rect 103330 3244 103336 3256
rect 70268 3216 103336 3244
rect 70268 3204 70274 3216
rect 103330 3204 103336 3216
rect 103388 3204 103394 3256
rect 160094 3204 160100 3256
rect 160152 3244 160158 3256
rect 291838 3244 291844 3256
rect 160152 3216 291844 3244
rect 160152 3204 160158 3216
rect 291838 3204 291844 3216
rect 291896 3204 291902 3256
rect 299474 3204 299480 3256
rect 299532 3244 299538 3256
rect 300762 3244 300768 3256
rect 299532 3216 300768 3244
rect 299532 3204 299538 3216
rect 300762 3204 300768 3216
rect 300820 3204 300826 3256
rect 316034 3204 316040 3256
rect 316092 3244 316098 3256
rect 317322 3244 317328 3256
rect 316092 3216 317328 3244
rect 316092 3204 316098 3216
rect 317322 3204 317328 3216
rect 317380 3204 317386 3256
rect 324406 3204 324412 3256
rect 324464 3244 324470 3256
rect 325602 3244 325608 3256
rect 324464 3216 325608 3244
rect 324464 3204 324470 3216
rect 325602 3204 325608 3216
rect 325660 3204 325666 3256
rect 332686 3204 332692 3256
rect 332744 3244 332750 3256
rect 333882 3244 333888 3256
rect 332744 3216 333888 3244
rect 332744 3204 332750 3216
rect 333882 3204 333888 3216
rect 333940 3204 333946 3256
rect 340966 3204 340972 3256
rect 341024 3244 341030 3256
rect 342162 3244 342168 3256
rect 341024 3216 342168 3244
rect 341024 3204 341030 3216
rect 342162 3204 342168 3216
rect 342220 3204 342226 3256
rect 349246 3204 349252 3256
rect 349304 3244 349310 3256
rect 350442 3244 350448 3256
rect 349304 3216 350448 3244
rect 349304 3204 349310 3216
rect 350442 3204 350448 3216
rect 350500 3204 350506 3256
rect 357526 3204 357532 3256
rect 357584 3244 357590 3256
rect 358722 3244 358728 3256
rect 357584 3216 358728 3244
rect 357584 3204 357590 3216
rect 358722 3204 358728 3216
rect 358780 3204 358786 3256
rect 365806 3204 365812 3256
rect 365864 3244 365870 3256
rect 367002 3244 367008 3256
rect 365864 3216 367008 3244
rect 365864 3204 365870 3216
rect 367002 3204 367008 3216
rect 367060 3204 367066 3256
rect 374086 3204 374092 3256
rect 374144 3244 374150 3256
rect 375282 3244 375288 3256
rect 374144 3216 375288 3244
rect 374144 3204 374150 3216
rect 375282 3204 375288 3216
rect 375340 3204 375346 3256
rect 382274 3204 382280 3256
rect 382332 3244 382338 3256
rect 383562 3244 383568 3256
rect 382332 3216 383568 3244
rect 382332 3204 382338 3216
rect 383562 3204 383568 3216
rect 383620 3204 383626 3256
rect 390646 3204 390652 3256
rect 390704 3244 390710 3256
rect 391842 3244 391848 3256
rect 390704 3216 391848 3244
rect 390704 3204 390710 3216
rect 391842 3204 391848 3216
rect 391900 3204 391906 3256
rect 398926 3204 398932 3256
rect 398984 3244 398990 3256
rect 400122 3244 400128 3256
rect 398984 3216 400128 3244
rect 398984 3204 398990 3216
rect 400122 3204 400128 3216
rect 400180 3204 400186 3256
rect 407114 3204 407120 3256
rect 407172 3244 407178 3256
rect 408402 3244 408408 3256
rect 407172 3216 408408 3244
rect 407172 3204 407178 3216
rect 408402 3204 408408 3216
rect 408460 3204 408466 3256
rect 431954 3204 431960 3256
rect 432012 3244 432018 3256
rect 433242 3244 433248 3256
rect 432012 3216 433248 3244
rect 432012 3204 432018 3216
rect 433242 3204 433248 3216
rect 433300 3204 433306 3256
rect 440326 3204 440332 3256
rect 440384 3244 440390 3256
rect 441522 3244 441528 3256
rect 440384 3216 441528 3244
rect 440384 3204 440390 3216
rect 441522 3204 441528 3216
rect 441580 3204 441586 3256
rect 566 3136 572 3188
rect 624 3176 630 3188
rect 3418 3176 3424 3188
rect 624 3148 3424 3176
rect 624 3136 630 3148
rect 3418 3136 3424 3148
rect 3476 3136 3482 3188
rect 226334 3136 226340 3188
rect 226392 3176 226398 3188
rect 227530 3176 227536 3188
rect 226392 3148 227536 3176
rect 226392 3136 226398 3148
rect 227530 3136 227536 3148
rect 227588 3136 227594 3188
rect 530578 3000 530584 3052
rect 530636 3040 530642 3052
rect 532510 3040 532516 3052
rect 530636 3012 532516 3040
rect 530636 3000 530642 3012
rect 532510 3000 532516 3012
rect 532568 3000 532574 3052
rect 9950 2932 9956 2984
rect 10008 2972 10014 2984
rect 11698 2972 11704 2984
rect 10008 2944 11704 2972
rect 10008 2932 10014 2944
rect 11698 2932 11704 2944
rect 11756 2932 11762 2984
<< via1 >>
rect 1400 386384 1452 386436
rect 57612 386384 57664 386436
rect 372160 59780 372212 59832
rect 373724 59780 373776 59832
rect 430120 59780 430172 59832
rect 431500 59780 431552 59832
rect 488080 59780 488132 59832
rect 489368 59780 489420 59832
rect 498476 59780 498528 59832
rect 499488 59780 499540 59832
rect 516968 59780 517020 59832
rect 518348 59780 518400 59832
rect 73068 59712 73120 59764
rect 74724 59712 74776 59764
rect 77944 59712 77996 59764
rect 79876 59712 79928 59764
rect 80704 59712 80756 59764
rect 83004 59712 83056 59764
rect 86224 59712 86276 59764
rect 87420 59712 87472 59764
rect 118608 59712 118660 59764
rect 120264 59712 120316 59764
rect 129004 59712 129056 59764
rect 131580 59712 131632 59764
rect 131764 59712 131816 59764
rect 132592 59712 132644 59764
rect 136548 59712 136600 59764
rect 137836 59712 137888 59764
rect 140044 59712 140096 59764
rect 141976 59712 142028 59764
rect 142804 59712 142856 59764
rect 145012 59712 145064 59764
rect 145748 59712 145800 59764
rect 148140 59712 148192 59764
rect 150348 59712 150400 59764
rect 152280 59712 152332 59764
rect 153844 59712 153896 59764
rect 156604 59712 156656 59764
rect 160744 59712 160796 59764
rect 162584 59712 162636 59764
rect 179236 59712 179288 59764
rect 181260 59712 181312 59764
rect 188896 59712 188948 59764
rect 190552 59712 190604 59764
rect 194508 59712 194560 59764
rect 195796 59712 195848 59764
rect 206928 59712 206980 59764
rect 208124 59712 208176 59764
rect 220452 59712 220504 59764
rect 222568 59712 222620 59764
rect 242808 59712 242860 59764
rect 244280 59712 244332 59764
rect 257896 59712 257948 59764
rect 259828 59712 259880 59764
rect 266268 59712 266320 59764
rect 268108 59712 268160 59764
rect 279424 59712 279476 59764
rect 280620 59712 280672 59764
rect 287704 59712 287756 59764
rect 289820 59712 289872 59764
rect 290648 59712 290700 59764
rect 292948 59712 293000 59764
rect 294604 59712 294656 59764
rect 297088 59712 297140 59764
rect 300124 59712 300176 59764
rect 302240 59712 302292 59764
rect 309048 59712 309100 59764
rect 310520 59712 310572 59764
rect 326712 59712 326764 59764
rect 329288 59712 329340 59764
rect 338028 59712 338080 59764
rect 339500 59712 339552 59764
rect 342168 59712 342220 59764
rect 344284 59712 344336 59764
rect 354680 59712 354732 59764
rect 356704 59712 356756 59764
rect 392860 59712 392912 59764
rect 394884 59712 394936 59764
rect 400128 59712 400180 59764
rect 401600 59712 401652 59764
rect 409512 59712 409564 59764
rect 411628 59712 411680 59764
rect 412640 59712 412692 59764
rect 414112 59712 414164 59764
rect 418712 59712 418764 59764
rect 419816 59712 419868 59764
rect 446680 59712 446732 59764
rect 449348 59712 449400 59764
rect 454960 59712 455012 59764
rect 457628 59712 457680 59764
rect 467288 59712 467340 59764
rect 468484 59712 468536 59764
rect 512828 59712 512880 59764
rect 514852 59712 514904 59764
rect 525248 59712 525300 59764
rect 527364 59712 527416 59764
rect 533712 59712 533764 59764
rect 535644 59712 535696 59764
rect 537668 59712 537720 59764
rect 539784 59712 539836 59764
rect 554320 59712 554372 59764
rect 556344 59712 556396 59764
rect 560392 59712 560444 59764
rect 561772 59712 561824 59764
rect 24860 59576 24912 59628
rect 60556 59576 60608 59628
rect 89168 59576 89220 59628
rect 91284 59576 91336 59628
rect 116584 59576 116636 59628
rect 118148 59576 118200 59628
rect 123484 59576 123536 59628
rect 125416 59576 125468 59628
rect 284944 59576 284996 59628
rect 286692 59576 286744 59628
rect 322204 59576 322256 59628
rect 325148 59576 325200 59628
rect 328736 59576 328788 59628
rect 330484 59576 330536 59628
rect 345296 59576 345348 59628
rect 347044 59576 347096 59628
rect 461124 59576 461176 59628
rect 462964 59576 463016 59628
rect 541808 59576 541860 59628
rect 544016 59576 544068 59628
rect 561496 59576 561548 59628
rect 563060 59576 563112 59628
rect 19340 59508 19392 59560
rect 62304 59508 62356 59560
rect 5540 59440 5592 59492
rect 57796 59440 57848 59492
rect 114008 59440 114060 59492
rect 116124 59440 116176 59492
rect 175096 59440 175148 59492
rect 177120 59440 177172 59492
rect 191748 59440 191800 59492
rect 193680 59440 193732 59492
rect 203892 59440 203944 59492
rect 206100 59440 206152 59492
rect 224868 59440 224920 59492
rect 226708 59440 226760 59492
rect 233056 59440 233108 59492
rect 234988 59440 235040 59492
rect 249708 59440 249760 59492
rect 251548 59440 251600 59492
rect 253756 59440 253808 59492
rect 255688 59440 255740 59492
rect 256608 59440 256660 59492
rect 257804 59440 257856 59492
rect 282184 59440 282236 59492
rect 284668 59440 284720 59492
rect 405280 59440 405332 59492
rect 407304 59440 407356 59492
rect 420828 59440 420880 59492
rect 422392 59440 422444 59492
rect 443552 59440 443604 59492
rect 444380 59440 444432 59492
rect 492128 59440 492180 59492
rect 494244 59440 494296 59492
rect 504548 59440 504600 59492
rect 506664 59440 506716 59492
rect 4160 59372 4212 59424
rect 58164 59372 58216 59424
rect 365812 59372 365864 59424
rect 366548 59372 366600 59424
rect 384488 59372 384540 59424
rect 385224 59372 385276 59424
rect 101956 59304 102008 59356
rect 103428 59304 103480 59356
rect 262220 59304 262272 59356
rect 263968 59304 264020 59356
rect 362224 59032 362276 59084
rect 389180 59032 389232 59084
rect 328460 58964 328512 59016
rect 376760 58964 376812 59016
rect 217968 58896 218020 58948
rect 425060 58896 425112 58948
rect 449716 58896 449768 58948
rect 536840 58896 536892 58948
rect 306196 58828 306248 58880
rect 572720 58828 572772 58880
rect 259460 58760 259512 58812
rect 529020 58760 529072 58812
rect 53840 58692 53892 58744
rect 150348 58692 150400 58744
rect 188988 58692 189040 58744
rect 524420 58692 524472 58744
rect 49700 58624 49752 58676
rect 85488 58624 85540 58676
rect 109868 58624 109920 58676
rect 110880 58624 110932 58676
rect 146300 58624 146352 58676
rect 561864 58624 561916 58676
rect 246948 58556 247000 58608
rect 248420 58556 248472 58608
rect 322112 58488 322164 58540
rect 323584 58488 323636 58540
rect 245292 58352 245344 58404
rect 246764 58352 246816 58404
rect 320456 58352 320508 58404
rect 322204 58352 322256 58404
rect 384120 58352 384172 58404
rect 385040 58352 385092 58404
rect 342260 57536 342312 57588
rect 374000 57536 374052 57588
rect 242716 57468 242768 57520
rect 340880 57468 340932 57520
rect 374092 57468 374144 57520
rect 495624 57468 495676 57520
rect 251180 57400 251232 57452
rect 266084 57400 266136 57452
rect 339500 57400 339552 57452
rect 466460 57400 466512 57452
rect 204260 57332 204312 57384
rect 413192 57332 413244 57384
rect 161480 57264 161532 57316
rect 425336 57264 425388 57316
rect 444564 57264 444616 57316
rect 557540 57264 557592 57316
rect 7564 57196 7616 57248
rect 164148 57196 164200 57248
rect 263600 57196 263652 57248
rect 528652 57196 528704 57248
rect 353300 56176 353352 56228
rect 420920 56176 420972 56228
rect 430580 56176 430632 56228
rect 481640 56176 481692 56228
rect 267740 56108 267792 56160
rect 394700 56108 394752 56160
rect 248420 56040 248472 56092
rect 266268 56040 266320 56092
rect 335360 56040 335412 56092
rect 481640 56040 481692 56092
rect 229008 55972 229060 56024
rect 379520 55972 379572 56024
rect 103520 55904 103572 55956
rect 136548 55904 136600 55956
rect 168380 55904 168432 55956
rect 423680 55904 423732 55956
rect 444380 55904 444432 55956
rect 561680 55904 561732 55956
rect 48320 55836 48372 55888
rect 118608 55836 118660 55888
rect 135260 55836 135312 55888
rect 567292 55836 567344 55888
rect 261944 54952 261996 55004
rect 266360 54952 266412 55004
rect 303620 54816 303672 54868
rect 386420 54816 386472 54868
rect 233056 54748 233108 54800
rect 361580 54748 361632 54800
rect 362132 54748 362184 54800
rect 391940 54748 391992 54800
rect 216496 54680 216548 54732
rect 418160 54680 418212 54732
rect 458180 54680 458232 54732
rect 473360 54680 473412 54732
rect 162860 54612 162912 54664
rect 290648 54612 290700 54664
rect 309048 54612 309100 54664
rect 556160 54612 556212 54664
rect 274640 54544 274692 54596
rect 527180 54544 527232 54596
rect 10324 54476 10376 54528
rect 162584 54476 162636 54528
rect 168472 54476 168524 54528
rect 556620 54476 556672 54528
rect 311624 53320 311676 53372
rect 545212 53320 545264 53372
rect 288440 53252 288492 53304
rect 523040 53252 523092 53304
rect 140780 53184 140832 53236
rect 434720 53184 434772 53236
rect 469220 53184 469272 53236
rect 476120 53184 476172 53236
rect 183468 53116 183520 53168
rect 530584 53116 530636 53168
rect 57980 53048 58032 53100
rect 149704 53048 149756 53100
rect 200120 53048 200172 53100
rect 549260 53048 549312 53100
rect 332600 51960 332652 52012
rect 488540 51960 488592 52012
rect 313280 51892 313332 51944
rect 516140 51892 516192 51944
rect 133880 51824 133932 51876
rect 436192 51824 436244 51876
rect 188896 51756 188948 51808
rect 514760 51756 514812 51808
rect 44180 51688 44232 51740
rect 154028 51688 154080 51740
rect 213920 51688 213972 51740
rect 545120 51688 545172 51740
rect 355324 50668 355376 50720
rect 414020 50668 414072 50720
rect 292580 50600 292632 50652
rect 390652 50600 390704 50652
rect 321008 50532 321060 50584
rect 531412 50532 531464 50584
rect 218060 50464 218112 50516
rect 543832 50464 543884 50516
rect 40040 50396 40092 50448
rect 153844 50396 153896 50448
rect 179236 50396 179288 50448
rect 546592 50396 546644 50448
rect 139400 50328 139452 50380
rect 567200 50328 567252 50380
rect 258080 49240 258132 49292
rect 400220 49240 400272 49292
rect 325148 49172 325200 49224
rect 520280 49172 520332 49224
rect 151820 49104 151872 49156
rect 294788 49104 294840 49156
rect 316040 49104 316092 49156
rect 515036 49104 515088 49156
rect 110512 49036 110564 49088
rect 133328 49036 133380 49088
rect 143540 49036 143592 49088
rect 433340 49036 433392 49088
rect 52460 48968 52512 49020
rect 117964 48968 118016 49020
rect 209780 48968 209832 49020
rect 546500 48968 546552 49020
rect 276020 47880 276072 47932
rect 394792 47880 394844 47932
rect 341708 47812 341760 47864
rect 463700 47812 463752 47864
rect 219348 47744 219400 47796
rect 411260 47744 411312 47796
rect 201500 47676 201552 47728
rect 279424 47676 279476 47728
rect 323584 47676 323636 47728
rect 523040 47676 523092 47728
rect 93860 47608 93912 47660
rect 138664 47608 138716 47660
rect 207020 47608 207072 47660
rect 547880 47608 547932 47660
rect 11704 47540 11756 47592
rect 95884 47540 95936 47592
rect 143632 47540 143684 47592
rect 565820 47540 565872 47592
rect 364340 47064 364392 47116
rect 369952 47064 370004 47116
rect 338120 46520 338172 46572
rect 509240 46520 509292 46572
rect 222108 46452 222160 46504
rect 400220 46452 400272 46504
rect 325700 46384 325752 46436
rect 513380 46384 513432 46436
rect 208400 46316 208452 46368
rect 415584 46316 415636 46368
rect 469864 46316 469916 46368
rect 473360 46316 473412 46368
rect 198648 46248 198700 46300
rect 481732 46248 481784 46300
rect 3424 46180 3476 46232
rect 164884 46180 164936 46232
rect 195980 46180 196032 46232
rect 550640 46180 550692 46232
rect 337568 45160 337620 45212
rect 473452 45160 473504 45212
rect 244188 45092 244240 45144
rect 325700 45092 325752 45144
rect 334624 45092 334676 45144
rect 484400 45092 484452 45144
rect 138020 45024 138072 45076
rect 298928 45024 298980 45076
rect 349160 45024 349212 45076
rect 506664 45024 506716 45076
rect 193220 44956 193272 45008
rect 419632 44956 419684 45008
rect 211068 44888 211120 44940
rect 440240 44888 440292 44940
rect 62120 44820 62172 44872
rect 114008 44820 114060 44872
rect 128360 44820 128412 44872
rect 569960 44820 570012 44872
rect 338764 43732 338816 43784
rect 470600 43732 470652 43784
rect 233240 43664 233292 43716
rect 407120 43664 407172 43716
rect 331220 43596 331272 43648
rect 510712 43596 510764 43648
rect 324964 43528 325016 43580
rect 516140 43528 516192 43580
rect 193312 43460 193364 43512
rect 552112 43460 552164 43512
rect 46940 43392 46992 43444
rect 152464 43392 152516 43444
rect 173808 43392 173860 43444
rect 566464 43392 566516 43444
rect 226248 42372 226300 42424
rect 386420 42372 386472 42424
rect 345020 42304 345072 42356
rect 506480 42304 506532 42356
rect 331864 42236 331916 42288
rect 495440 42236 495492 42288
rect 197268 42168 197320 42220
rect 485780 42168 485832 42220
rect 129740 42100 129792 42152
rect 437480 42100 437532 42152
rect 80060 42032 80112 42084
rect 109868 42032 109920 42084
rect 189080 42032 189132 42084
rect 552296 42032 552348 42084
rect 241336 40944 241388 40996
rect 336740 40944 336792 40996
rect 337384 40944 337436 40996
rect 477500 40944 477552 40996
rect 333980 40876 334032 40928
rect 510896 40876 510948 40928
rect 131120 40808 131172 40860
rect 300124 40808 300176 40860
rect 329288 40808 329340 40860
rect 506480 40808 506532 40860
rect 215300 40740 215352 40792
rect 412640 40740 412692 40792
rect 27620 40672 27672 40724
rect 125048 40672 125100 40724
rect 182180 40672 182232 40724
rect 554780 40672 554832 40724
rect 251272 39652 251324 39704
rect 402980 39652 403032 39704
rect 224684 39584 224736 39636
rect 393320 39584 393372 39636
rect 327724 39516 327776 39568
rect 509240 39516 509292 39568
rect 327080 39448 327132 39500
rect 512000 39448 512052 39500
rect 151912 39380 151964 39432
rect 431960 39380 432012 39432
rect 52552 39312 52604 39364
rect 84844 39312 84896 39364
rect 178040 39312 178092 39364
rect 556344 39312 556396 39364
rect 253940 38224 253992 38276
rect 401600 38224 401652 38276
rect 220636 38156 220688 38208
rect 407120 38156 407172 38208
rect 324320 38088 324372 38140
rect 513472 38088 513524 38140
rect 322204 38020 322256 38072
rect 527180 38020 527232 38072
rect 158720 37952 158772 38004
rect 429200 37952 429252 38004
rect 448520 37952 448572 38004
rect 477776 37952 477828 38004
rect 20720 37884 20772 37936
rect 159364 37884 159416 37936
rect 175280 37884 175332 37936
rect 556528 37884 556580 37936
rect 230388 36796 230440 36848
rect 372620 36796 372672 36848
rect 292672 36728 292724 36780
rect 523224 36728 523276 36780
rect 249616 36660 249668 36712
rect 305000 36660 305052 36712
rect 310428 36660 310480 36712
rect 552020 36660 552072 36712
rect 136640 36592 136692 36644
rect 436376 36592 436428 36644
rect 444380 36592 444432 36644
rect 477592 36592 477644 36644
rect 171140 36524 171192 36576
rect 557632 36524 557684 36576
rect 364984 35572 365036 35624
rect 382556 35572 382608 35624
rect 332600 35504 332652 35556
rect 378232 35504 378284 35556
rect 352564 35436 352616 35488
rect 423956 35436 424008 35488
rect 231768 35368 231820 35420
rect 368480 35368 368532 35420
rect 423772 35368 423824 35420
rect 484492 35368 484544 35420
rect 179420 35300 179472 35352
rect 423680 35300 423732 35352
rect 446404 35300 446456 35352
rect 554780 35300 554832 35352
rect 256700 35232 256752 35284
rect 532700 35232 532752 35284
rect 153200 35164 153252 35216
rect 563060 35164 563112 35216
rect 358268 34076 358320 34128
rect 402980 34076 403032 34128
rect 317420 34008 317472 34060
rect 382280 34008 382332 34060
rect 190460 33940 190512 33992
rect 419816 33940 419868 33992
rect 447784 33940 447836 33992
rect 550640 33940 550692 33992
rect 252560 33872 252612 33924
rect 534080 33872 534132 33924
rect 51080 33804 51132 33856
rect 151084 33804 151136 33856
rect 180708 33804 180760 33856
rect 542360 33804 542412 33856
rect 150440 33736 150492 33788
rect 564624 33736 564676 33788
rect 289820 32716 289872 32768
rect 390836 32716 390888 32768
rect 356704 32648 356756 32700
rect 409880 32648 409932 32700
rect 224868 32580 224920 32632
rect 390560 32580 390612 32632
rect 437480 32580 437532 32632
rect 480260 32580 480312 32632
rect 212540 32512 212592 32564
rect 276664 32512 276716 32564
rect 277400 32512 277452 32564
rect 527364 32512 527416 32564
rect 184940 32444 184992 32496
rect 284944 32444 284996 32496
rect 307576 32444 307628 32496
rect 563060 32444 563112 32496
rect 26240 32376 26292 32428
rect 158168 32376 158220 32428
rect 164240 32376 164292 32428
rect 560392 32376 560444 32428
rect 296720 31288 296772 31340
rect 389272 31288 389324 31340
rect 398840 31288 398892 31340
rect 491300 31288 491352 31340
rect 149060 31220 149112 31272
rect 294604 31220 294656 31272
rect 303344 31220 303396 31272
rect 576124 31220 576176 31272
rect 242900 31152 242952 31204
rect 536932 31152 536984 31204
rect 126980 31084 127032 31136
rect 438860 31084 438912 31136
rect 449348 31084 449400 31136
rect 547880 31084 547932 31136
rect 41420 31016 41472 31068
rect 120908 31016 120960 31068
rect 179052 31016 179104 31068
rect 547144 31016 547196 31068
rect 394700 29928 394752 29980
rect 492680 29928 492732 29980
rect 260840 29860 260892 29912
rect 399116 29860 399168 29912
rect 330484 29792 330536 29844
rect 498200 29792 498252 29844
rect 165620 29724 165672 29776
rect 428004 29724 428056 29776
rect 449164 29724 449216 29776
rect 543740 29724 543792 29776
rect 224960 29656 225012 29708
rect 542452 29656 542504 29708
rect 34520 29588 34572 29640
rect 122104 29588 122156 29640
rect 183192 29588 183244 29640
rect 535460 29588 535512 29640
rect 387800 28568 387852 28620
rect 494060 28568 494112 28620
rect 271880 28500 271932 28552
rect 396080 28500 396132 28552
rect 329104 28432 329156 28484
rect 502340 28432 502392 28484
rect 172520 28364 172572 28416
rect 425152 28364 425204 28416
rect 450544 28364 450596 28416
rect 539876 28364 539928 28416
rect 220820 28296 220872 28348
rect 544016 28296 544068 28348
rect 16580 28228 16632 28280
rect 160744 28228 160796 28280
rect 182088 28228 182140 28280
rect 538864 28228 538916 28280
rect 187700 27208 187752 27260
rect 283564 27208 283616 27260
rect 353944 27208 353996 27260
rect 416780 27208 416832 27260
rect 282920 27140 282972 27192
rect 393412 27140 393464 27192
rect 217968 27072 218020 27124
rect 415400 27072 415452 27124
rect 433340 27072 433392 27124
rect 481824 27072 481876 27124
rect 270500 27004 270552 27056
rect 528560 27004 528612 27056
rect 135352 26936 135404 26988
rect 298744 26936 298796 26988
rect 306288 26936 306340 26988
rect 565820 26936 565872 26988
rect 17960 26868 18012 26920
rect 126244 26868 126296 26920
rect 160100 26868 160152 26920
rect 560576 26868 560628 26920
rect 307760 25848 307812 25900
rect 386604 25848 386656 25900
rect 383660 25780 383712 25832
rect 495532 25780 495584 25832
rect 236000 25712 236052 25764
rect 407304 25712 407356 25764
rect 461768 25712 461820 25764
rect 500960 25712 501012 25764
rect 202880 25644 202932 25696
rect 548064 25644 548116 25696
rect 29000 25576 29052 25628
rect 157984 25576 158036 25628
rect 177948 25576 178000 25628
rect 553492 25576 553544 25628
rect 157340 25508 157392 25560
rect 561772 25508 561824 25560
rect 278780 24420 278832 24472
rect 394884 24420 394936 24472
rect 376760 24352 376812 24404
rect 498384 24352 498436 24404
rect 333244 24284 333296 24336
rect 491300 24284 491352 24336
rect 176660 24216 176712 24268
rect 423864 24216 423916 24268
rect 464344 24216 464396 24268
rect 494060 24216 494112 24268
rect 184848 24148 184900 24200
rect 528560 24148 528612 24200
rect 74448 24080 74500 24132
rect 88340 24080 88392 24132
rect 185032 24080 185084 24132
rect 553400 24080 553452 24132
rect 98000 23808 98052 23860
rect 104164 23808 104216 23860
rect 194600 23060 194652 23112
rect 282368 23060 282420 23112
rect 357440 23060 357492 23112
rect 371240 23060 371292 23112
rect 264980 22992 265032 23044
rect 398932 22992 398984 23044
rect 223488 22924 223540 22976
rect 397460 22924 397512 22976
rect 426440 22924 426492 22976
rect 483020 22924 483072 22976
rect 267832 22856 267884 22908
rect 529940 22856 529992 22908
rect 144920 22788 144972 22840
rect 295984 22788 296036 22840
rect 304908 22788 304960 22840
rect 569960 22788 570012 22840
rect 77300 22720 77352 22772
rect 109684 22720 109736 22772
rect 125600 22720 125652 22772
rect 571340 22720 571392 22772
rect 349252 21700 349304 21752
rect 374092 21700 374144 21752
rect 220452 21632 220504 21684
rect 404360 21632 404412 21684
rect 408500 21632 408552 21684
rect 488632 21632 488684 21684
rect 216312 21564 216364 21616
rect 422300 21564 422352 21616
rect 213828 21496 213880 21548
rect 429200 21496 429252 21548
rect 462320 21496 462372 21548
rect 473544 21496 473596 21548
rect 212356 21428 212408 21480
rect 431960 21428 432012 21480
rect 465908 21428 465960 21480
rect 490196 21428 490248 21480
rect 35900 21360 35952 21412
rect 155224 21360 155276 21412
rect 212172 21360 212224 21412
rect 436100 21360 436152 21412
rect 443644 21360 443696 21412
rect 564440 21360 564492 21412
rect 228732 20408 228784 20460
rect 375380 20408 375432 20460
rect 227628 20340 227680 20392
rect 382372 20340 382424 20392
rect 176568 20272 176620 20324
rect 556252 20272 556304 20324
rect 175096 20204 175148 20256
rect 560300 20204 560352 20256
rect 174912 20136 174964 20188
rect 564532 20136 564584 20188
rect 172428 20068 172480 20120
rect 571340 20068 571392 20120
rect 170772 20000 170824 20052
rect 574100 20000 574152 20052
rect 33140 19932 33192 19984
rect 156604 19932 156656 19984
rect 170956 19932 171008 19984
rect 578240 19932 578292 19984
rect 195796 19116 195848 19168
rect 490012 19116 490064 19168
rect 195612 19048 195664 19100
rect 492680 19048 492732 19100
rect 194508 18980 194560 19032
rect 496912 18980 496964 19032
rect 193128 18912 193180 18964
rect 499580 18912 499632 18964
rect 191656 18844 191708 18896
rect 503720 18844 503772 18896
rect 191472 18776 191524 18828
rect 506572 18776 506624 18828
rect 190368 18708 190420 18760
rect 510620 18708 510672 18760
rect 187516 18640 187568 18692
rect 517520 18640 517572 18692
rect 67640 18572 67692 18624
rect 80888 18572 80940 18624
rect 86960 18572 87012 18624
rect 106924 18572 106976 18624
rect 107660 18572 107712 18624
rect 134524 18572 134576 18624
rect 187332 18572 187384 18624
rect 521660 18572 521712 18624
rect 351184 17824 351236 17876
rect 427820 17824 427872 17876
rect 349804 17756 349856 17808
rect 432052 17756 432104 17808
rect 349988 17688 350040 17740
rect 434720 17688 434772 17740
rect 348424 17620 348476 17672
rect 438860 17620 438912 17672
rect 440332 17620 440384 17672
rect 478880 17620 478932 17672
rect 347044 17552 347096 17604
rect 441620 17552 441672 17604
rect 251088 17484 251140 17536
rect 300860 17484 300912 17536
rect 345664 17484 345716 17536
rect 445760 17484 445812 17536
rect 209872 17416 209924 17468
rect 278228 17416 278280 17468
rect 345848 17416 345900 17468
rect 448612 17416 448664 17468
rect 451280 17416 451332 17468
rect 476212 17416 476264 17468
rect 241152 17348 241204 17400
rect 332692 17348 332744 17400
rect 344284 17348 344336 17400
rect 452660 17348 452712 17400
rect 63500 17280 63552 17332
rect 80704 17280 80756 17332
rect 169760 17280 169812 17332
rect 289084 17280 289136 17332
rect 342904 17280 342956 17332
rect 456892 17280 456944 17332
rect 465724 17280 465776 17332
rect 487160 17280 487212 17332
rect 72884 17212 72936 17264
rect 95240 17212 95292 17264
rect 100760 17212 100812 17264
rect 137468 17212 137520 17264
rect 154580 17212 154632 17264
rect 430672 17212 430724 17264
rect 456064 17212 456116 17264
rect 523132 17212 523184 17264
rect 238668 16192 238720 16244
rect 344560 16192 344612 16244
rect 366548 16192 366600 16244
rect 374092 16192 374144 16244
rect 237196 16124 237248 16176
rect 348056 16124 348108 16176
rect 363604 16124 363656 16176
rect 385960 16124 386012 16176
rect 237012 16056 237064 16108
rect 351184 16056 351236 16108
rect 360844 16056 360896 16108
rect 396080 16056 396132 16108
rect 467104 16056 467156 16108
rect 484032 16056 484084 16108
rect 234528 15988 234580 16040
rect 357532 15988 357584 16040
rect 358084 15988 358136 16040
rect 407212 15988 407264 16040
rect 420184 15988 420236 16040
rect 485964 15988 486016 16040
rect 232872 15920 232924 15972
rect 365720 15920 365772 15972
rect 366364 15920 366416 15972
rect 378324 15920 378376 15972
rect 381176 15920 381228 15972
rect 496820 15920 496872 15972
rect 73344 15852 73396 15904
rect 111064 15852 111116 15904
rect 114744 15852 114796 15904
rect 133144 15852 133196 15904
rect 147864 15852 147916 15904
rect 432144 15852 432196 15904
rect 461584 15852 461636 15904
rect 505376 15852 505428 15904
rect 367744 15308 367796 15360
rect 371240 15308 371292 15360
rect 260748 14696 260800 14748
rect 270040 14696 270092 14748
rect 320824 14696 320876 14748
rect 534448 14696 534500 14748
rect 249432 14628 249484 14680
rect 307852 14628 307904 14680
rect 319444 14628 319496 14680
rect 538220 14628 538272 14680
rect 198740 14560 198792 14612
rect 280804 14560 280856 14612
rect 318064 14560 318116 14612
rect 541992 14560 542044 14612
rect 101956 14492 102008 14544
rect 105636 14492 105688 14544
rect 167184 14492 167236 14544
rect 290464 14492 290516 14544
rect 311808 14492 311860 14544
rect 548616 14492 548668 14544
rect 66720 14424 66772 14476
rect 113824 14424 113876 14476
rect 128176 14424 128228 14476
rect 301504 14424 301556 14476
rect 307392 14424 307444 14476
rect 559288 14424 559340 14476
rect 469864 13744 469916 13796
rect 470692 13744 470744 13796
rect 248328 13472 248380 13524
rect 312176 13472 312228 13524
rect 353576 13472 353628 13524
rect 372712 13472 372764 13524
rect 246948 13404 247000 13456
rect 316224 13404 316276 13456
rect 359464 13404 359516 13456
rect 398932 13404 398984 13456
rect 245292 13336 245344 13388
rect 319720 13336 319772 13388
rect 322112 13336 322164 13388
rect 382464 13336 382516 13388
rect 311440 13268 311492 13320
rect 385040 13268 385092 13320
rect 468484 13268 468536 13320
rect 480536 13268 480588 13320
rect 245476 13200 245528 13252
rect 322940 13200 322992 13252
rect 336280 13200 336332 13252
rect 378416 13200 378468 13252
rect 402520 13200 402572 13252
rect 489920 13200 489972 13252
rect 73068 13132 73120 13184
rect 92480 13132 92532 13184
rect 94412 13132 94464 13184
rect 105728 13132 105780 13184
rect 242808 13132 242860 13184
rect 330392 13132 330444 13184
rect 341524 13132 341576 13184
rect 459928 13132 459980 13184
rect 462964 13132 463016 13184
rect 498292 13132 498344 13184
rect 60832 13064 60884 13116
rect 82084 13064 82136 13116
rect 97448 13064 97500 13116
rect 137284 13064 137336 13116
rect 156144 13064 156196 13116
rect 293224 13064 293276 13116
rect 320456 13064 320508 13116
rect 514852 13064 514904 13116
rect 465816 12928 465868 12980
rect 471980 12928 472032 12980
rect 259368 12248 259420 12300
rect 273260 12248 273312 12300
rect 257896 12180 257948 12232
rect 276664 12180 276716 12232
rect 257712 12112 257764 12164
rect 280712 12112 280764 12164
rect 255228 12044 255280 12096
rect 287336 12044 287388 12096
rect 346952 12044 347004 12096
rect 374276 12044 374328 12096
rect 253756 11976 253808 12028
rect 291384 11976 291436 12028
rect 339500 11976 339552 12028
rect 376852 11976 376904 12028
rect 253572 11908 253624 11960
rect 294880 11908 294932 11960
rect 324412 11908 324464 11960
rect 380992 11908 381044 11960
rect 455696 11908 455748 11960
rect 474740 11908 474792 11960
rect 252468 11840 252520 11892
rect 298100 11840 298152 11892
rect 314660 11840 314712 11892
rect 383752 11840 383804 11892
rect 412640 11840 412692 11892
rect 487252 11840 487304 11892
rect 71688 11772 71740 11824
rect 99840 11772 99892 11824
rect 102048 11772 102100 11824
rect 109040 11772 109092 11824
rect 256608 11772 256660 11824
rect 284300 11772 284352 11824
rect 286600 11772 286652 11824
rect 392032 11772 392084 11824
rect 405740 11772 405792 11824
rect 490104 11772 490156 11824
rect 56784 11704 56836 11756
rect 83464 11704 83516 11756
rect 89904 11704 89956 11756
rect 140044 11704 140096 11756
rect 143540 11704 143592 11756
rect 144736 11704 144788 11756
rect 142160 11636 142212 11688
rect 297364 11704 297416 11756
rect 299480 11704 299532 11756
rect 387892 11704 387944 11756
rect 390652 11704 390704 11756
rect 494244 11704 494296 11756
rect 259460 11636 259512 11688
rect 260656 11636 260708 11688
rect 259460 10956 259512 11008
rect 262864 10956 262916 11008
rect 361120 10820 361172 10872
rect 370136 10820 370188 10872
rect 245200 10684 245252 10736
rect 267004 10684 267056 10736
rect 370136 10684 370188 10736
rect 499672 10684 499724 10736
rect 237656 10616 237708 10668
rect 269948 10616 270000 10668
rect 365812 10616 365864 10668
rect 501052 10616 501104 10668
rect 234620 10548 234672 10600
rect 269764 10548 269816 10600
rect 363512 10548 363564 10600
rect 502524 10548 502576 10600
rect 226340 10480 226392 10532
rect 272524 10480 272576 10532
rect 359464 10480 359516 10532
rect 502708 10480 502760 10532
rect 235908 10412 235960 10464
rect 355232 10412 355284 10464
rect 356336 10412 356388 10464
rect 503812 10412 503864 10464
rect 91560 10344 91612 10396
rect 105544 10344 105596 10396
rect 223580 10344 223632 10396
rect 274088 10344 274140 10396
rect 352840 10344 352892 10396
rect 505192 10344 505244 10396
rect 65064 10276 65116 10328
rect 146944 10276 146996 10328
rect 219992 10276 220044 10328
rect 273904 10276 273956 10328
rect 340972 10276 341024 10328
rect 507860 10276 507912 10328
rect 77024 9596 77076 9648
rect 78588 9596 78640 9648
rect 151728 9596 151780 9648
rect 153016 9596 153068 9648
rect 255872 9460 255924 9512
rect 264244 9460 264296 9512
rect 241704 9392 241756 9444
rect 268384 9392 268436 9444
rect 231032 9324 231084 9376
rect 271144 9324 271196 9376
rect 310244 9324 310296 9376
rect 517612 9324 517664 9376
rect 216864 9256 216916 9308
rect 275284 9256 275336 9308
rect 306748 9256 306800 9308
rect 518992 9256 519044 9308
rect 181444 9188 181496 9240
rect 286508 9188 286560 9240
rect 303160 9188 303212 9240
rect 519176 9188 519228 9240
rect 177856 9120 177908 9172
rect 286324 9120 286376 9172
rect 299664 9120 299716 9172
rect 520372 9120 520424 9172
rect 174268 9052 174320 9104
rect 287704 9052 287756 9104
rect 296076 9052 296128 9104
rect 521752 9052 521804 9104
rect 84476 8984 84528 9036
rect 108304 8984 108356 9036
rect 192024 8984 192076 9036
rect 282184 8984 282236 9036
rect 285404 8984 285456 9036
rect 524512 8984 524564 9036
rect 62028 8916 62080 8968
rect 148324 8916 148376 8968
rect 206192 8916 206244 8968
rect 278044 8916 278096 8968
rect 281908 8916 281960 8968
rect 525800 8916 525852 8968
rect 249984 7964 250036 8016
rect 535644 7964 535696 8016
rect 246396 7896 246448 7948
rect 535828 7896 535880 7948
rect 45468 7828 45520 7880
rect 119344 7828 119396 7880
rect 239312 7828 239364 7880
rect 538312 7828 538364 7880
rect 38384 7760 38436 7812
rect 120724 7760 120776 7812
rect 235816 7760 235868 7812
rect 539784 7760 539836 7812
rect 31300 7692 31352 7744
rect 123484 7692 123536 7744
rect 232228 7692 232280 7744
rect 539600 7692 539652 7744
rect 23020 7624 23072 7676
rect 124864 7624 124916 7676
rect 228732 7624 228784 7676
rect 541072 7624 541124 7676
rect 13544 7556 13596 7608
rect 127624 7556 127676 7608
rect 132960 7556 133012 7608
rect 568856 7556 568908 7608
rect 523040 7488 523092 7540
rect 523868 7488 523920 7540
rect 247592 6536 247644 6588
rect 403164 6536 403216 6588
rect 75828 6468 75880 6520
rect 85672 6468 85724 6520
rect 244096 6468 244148 6520
rect 404452 6468 404504 6520
rect 70308 6400 70360 6452
rect 112444 6400 112496 6452
rect 240508 6400 240560 6452
rect 405832 6400 405884 6452
rect 59636 6332 59688 6384
rect 115204 6332 115256 6384
rect 229836 6332 229888 6384
rect 408592 6332 408644 6384
rect 416688 6332 416740 6384
rect 486148 6332 486200 6384
rect 56048 6264 56100 6316
rect 116584 6264 116636 6316
rect 226432 6264 226484 6316
rect 409972 6264 410024 6316
rect 442264 6264 442316 6316
rect 569132 6264 569184 6316
rect 14740 6196 14792 6248
rect 94504 6196 94556 6248
rect 222752 6196 222804 6248
rect 411628 6196 411680 6248
rect 441068 6196 441120 6248
rect 572720 6196 572772 6248
rect 8760 6128 8812 6180
rect 129188 6128 129240 6180
rect 219256 6128 219308 6180
rect 411444 6128 411496 6180
rect 440884 6128 440936 6180
rect 576308 6128 576360 6180
rect 77208 5516 77260 5568
rect 82084 5516 82136 5568
rect 86868 5244 86920 5296
rect 141424 5244 141476 5296
rect 71504 5176 71556 5228
rect 79324 5176 79376 5228
rect 83280 5176 83332 5228
rect 141608 5176 141660 5228
rect 460204 5176 460256 5228
rect 508872 5176 508924 5228
rect 79692 5108 79744 5160
rect 142804 5108 142856 5160
rect 458824 5108 458876 5160
rect 512460 5108 512512 5160
rect 76196 5040 76248 5092
rect 144184 5040 144236 5092
rect 197912 5040 197964 5092
rect 72608 4972 72660 5024
rect 145564 4972 145616 5024
rect 69112 4904 69164 4956
rect 145748 4904 145800 4956
rect 212172 5040 212224 5092
rect 414112 5040 414164 5092
rect 457444 5040 457496 5092
rect 515956 5040 516008 5092
rect 201592 4972 201644 5024
rect 416872 4972 416924 5024
rect 457628 4972 457680 5024
rect 519544 4972 519596 5024
rect 418252 4904 418304 4956
rect 454684 4904 454736 4956
rect 526628 4904 526680 4956
rect 4068 4836 4120 4888
rect 129004 4836 129056 4888
rect 187332 4836 187384 4888
rect 421012 4836 421064 4888
rect 453396 4836 453448 4888
rect 516784 4836 516836 4888
rect 12348 4768 12400 4820
rect 162124 4768 162176 4820
rect 183744 4768 183796 4820
rect 422392 4768 422444 4820
rect 453488 4768 453540 4820
rect 533712 4768 533764 4820
rect 516784 4700 516836 4752
rect 530124 4700 530176 4752
rect 75000 4156 75052 4208
rect 77944 4156 77996 4208
rect 209780 4156 209832 4208
rect 210976 4156 211028 4208
rect 251180 4156 251232 4208
rect 252376 4156 252428 4208
rect 267740 4156 267792 4208
rect 268476 4156 268528 4208
rect 292580 4156 292632 4208
rect 293316 4156 293368 4208
rect 307852 4156 307904 4208
rect 309048 4156 309100 4208
rect 68652 4088 68704 4140
rect 110512 4088 110564 4140
rect 208032 4088 208084 4140
rect 450912 4088 450964 4140
rect 566464 4088 566516 4140
rect 568028 4088 568080 4140
rect 576124 4088 576176 4140
rect 577412 4088 577464 4140
rect 43076 4020 43128 4072
rect 87604 4020 87656 4072
rect 206928 4020 206980 4072
rect 454500 4020 454552 4072
rect 67548 3952 67600 4004
rect 114008 3952 114060 4004
rect 205548 3952 205600 4004
rect 458088 3952 458140 4004
rect 547144 3952 547196 4004
rect 550272 3952 550324 4004
rect 39580 3884 39632 3936
rect 88984 3884 89036 3936
rect 203892 3884 203944 3936
rect 461584 3884 461636 3936
rect 66168 3816 66220 3868
rect 117596 3816 117648 3868
rect 204076 3816 204128 3868
rect 465172 3816 465224 3868
rect 35992 3748 36044 3800
rect 89260 3748 89312 3800
rect 100668 3748 100720 3800
rect 112812 3748 112864 3800
rect 202788 3748 202840 3800
rect 468668 3748 468720 3800
rect 15936 3680 15988 3732
rect 61384 3680 61436 3732
rect 64696 3680 64748 3732
rect 121092 3680 121144 3732
rect 201408 3680 201460 3732
rect 472256 3680 472308 3732
rect 32404 3612 32456 3664
rect 90364 3612 90416 3664
rect 99288 3612 99340 3664
rect 116400 3612 116452 3664
rect 118792 3612 118844 3664
rect 131764 3612 131816 3664
rect 168288 3612 168340 3664
rect 11152 3544 11204 3596
rect 62764 3544 62816 3596
rect 64512 3544 64564 3596
rect 124680 3544 124732 3596
rect 130384 3544 130436 3596
rect 135260 3544 135312 3596
rect 136456 3544 136508 3596
rect 168380 3544 168432 3596
rect 169576 3544 169628 3596
rect 193220 3612 193272 3664
rect 194416 3612 194468 3664
rect 199752 3612 199804 3664
rect 475752 3612 475804 3664
rect 581000 3544 581052 3596
rect 7656 3476 7708 3528
rect 10324 3476 10376 3528
rect 28908 3476 28960 3528
rect 91744 3476 91796 3528
rect 97816 3476 97868 3528
rect 119896 3476 119948 3528
rect 122288 3476 122340 3528
rect 160100 3476 160152 3528
rect 161296 3476 161348 3528
rect 199936 3476 199988 3528
rect 479340 3476 479392 3528
rect 498200 3476 498252 3528
rect 499028 3476 499080 3528
rect 538864 3476 538916 3528
rect 539600 3476 539652 3528
rect 564440 3476 564492 3528
rect 565268 3476 565320 3528
rect 24216 3408 24268 3460
rect 93308 3408 93360 3460
rect 97632 3408 97684 3460
rect 123484 3408 123536 3460
rect 166632 3408 166684 3460
rect 582196 3408 582248 3460
rect 46664 3340 46716 3392
rect 86224 3340 86276 3392
rect 201500 3340 201552 3392
rect 202696 3340 202748 3392
rect 208216 3340 208268 3392
rect 447416 3340 447468 3392
rect 448612 3340 448664 3392
rect 449808 3340 449860 3392
rect 2872 3272 2924 3324
rect 7564 3272 7616 3324
rect 68836 3272 68888 3324
rect 106924 3272 106976 3324
rect 209688 3272 209740 3324
rect 443828 3272 443880 3324
rect 70216 3204 70268 3256
rect 103336 3204 103388 3256
rect 160100 3204 160152 3256
rect 291844 3204 291896 3256
rect 299480 3204 299532 3256
rect 300768 3204 300820 3256
rect 316040 3204 316092 3256
rect 317328 3204 317380 3256
rect 324412 3204 324464 3256
rect 325608 3204 325660 3256
rect 332692 3204 332744 3256
rect 333888 3204 333940 3256
rect 340972 3204 341024 3256
rect 342168 3204 342220 3256
rect 349252 3204 349304 3256
rect 350448 3204 350500 3256
rect 357532 3204 357584 3256
rect 358728 3204 358780 3256
rect 365812 3204 365864 3256
rect 367008 3204 367060 3256
rect 374092 3204 374144 3256
rect 375288 3204 375340 3256
rect 382280 3204 382332 3256
rect 383568 3204 383620 3256
rect 390652 3204 390704 3256
rect 391848 3204 391900 3256
rect 398932 3204 398984 3256
rect 400128 3204 400180 3256
rect 407120 3204 407172 3256
rect 408408 3204 408460 3256
rect 431960 3204 432012 3256
rect 433248 3204 433300 3256
rect 440332 3204 440384 3256
rect 441528 3204 441580 3256
rect 572 3136 624 3188
rect 3424 3136 3476 3188
rect 226340 3136 226392 3188
rect 227536 3136 227588 3188
rect 530584 3000 530636 3052
rect 532516 3000 532568 3052
rect 9956 2932 10008 2984
rect 11704 2932 11756 2984
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 57610 387696 57666 387705
rect 57610 387631 57666 387640
rect 57624 386442 57652 387631
rect 1400 386436 1452 386442
rect 1400 386378 1452 386384
rect 57612 386436 57664 386442
rect 57612 386378 57664 386384
rect 572 3188 624 3194
rect 572 3130 624 3136
rect 584 480 612 3130
rect 542 -960 654 480
rect 1412 354 1440 386378
rect 372160 59832 372212 59838
rect 60646 59800 60702 59809
rect 66442 59800 66498 59809
rect 60646 59735 60702 59744
rect 65996 59758 66442 59786
rect 60554 59664 60610 59673
rect 24860 59628 24912 59634
rect 60554 59599 60556 59608
rect 24860 59570 24912 59576
rect 60608 59599 60610 59608
rect 60556 59570 60608 59576
rect 19340 59560 19392 59566
rect 19340 59502 19392 59508
rect 5540 59492 5592 59498
rect 5540 59434 5592 59440
rect 4160 59424 4212 59430
rect 4160 59366 4212 59372
rect 3424 46232 3476 46238
rect 3424 46174 3476 46180
rect 2872 3324 2924 3330
rect 2872 3266 2924 3272
rect 2884 480 2912 3266
rect 3436 3194 3464 46174
rect 4172 16574 4200 59366
rect 5552 16574 5580 59434
rect 7564 57248 7616 57254
rect 7564 57190 7616 57196
rect 4172 16546 5304 16574
rect 5552 16546 6040 16574
rect 4068 4888 4120 4894
rect 4068 4830 4120 4836
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 4080 480 4108 4830
rect 5276 480 5304 16546
rect 1646 354 1758 480
rect 1412 326 1758 354
rect 1646 -960 1758 326
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6012 354 6040 16546
rect 7576 3330 7604 57190
rect 10324 54528 10376 54534
rect 10324 54470 10376 54476
rect 8760 6180 8812 6186
rect 8760 6122 8812 6128
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7564 3324 7616 3330
rect 7564 3266 7616 3272
rect 7668 480 7696 3470
rect 8772 480 8800 6122
rect 10336 3534 10364 54470
rect 11704 47592 11756 47598
rect 11704 47534 11756 47540
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 9956 2984 10008 2990
rect 9956 2926 10008 2932
rect 9968 480 9996 2926
rect 11164 480 11192 3538
rect 11716 2990 11744 47534
rect 16580 28280 16632 28286
rect 16580 28222 16632 28228
rect 16592 16574 16620 28222
rect 17960 26920 18012 26926
rect 17960 26862 18012 26868
rect 16592 16546 17080 16574
rect 13544 7608 13596 7614
rect 13544 7550 13596 7556
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 11704 2984 11756 2990
rect 11704 2926 11756 2932
rect 12360 480 12388 4762
rect 13556 480 13584 7550
rect 14740 6248 14792 6254
rect 14740 6190 14792 6196
rect 14752 480 14780 6190
rect 15936 3732 15988 3738
rect 15936 3674 15988 3680
rect 15948 480 15976 3674
rect 17052 480 17080 16546
rect 6430 354 6542 480
rect 6012 326 6542 354
rect 6430 -960 6542 326
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 26862
rect 19352 16574 19380 59502
rect 20720 37936 20772 37942
rect 20720 37878 20772 37884
rect 20732 16574 20760 37878
rect 24872 16574 24900 59570
rect 57794 59528 57850 59537
rect 57794 59463 57796 59472
rect 57848 59463 57850 59472
rect 57796 59434 57848 59440
rect 58164 59424 58216 59430
rect 58162 59392 58164 59401
rect 60660 59401 60688 59735
rect 62302 59664 62358 59673
rect 62302 59599 62358 59608
rect 62316 59566 62344 59599
rect 62304 59560 62356 59566
rect 61382 59528 61438 59537
rect 62304 59502 62356 59508
rect 64510 59528 64566 59537
rect 61382 59463 61438 59472
rect 64510 59463 64566 59472
rect 58216 59392 58218 59401
rect 58162 59327 58218 59336
rect 60646 59392 60702 59401
rect 60646 59327 60702 59336
rect 53840 58744 53892 58750
rect 53840 58686 53892 58692
rect 49700 58676 49752 58682
rect 49700 58618 49752 58624
rect 48320 55888 48372 55894
rect 48320 55830 48372 55836
rect 44180 51740 44232 51746
rect 44180 51682 44232 51688
rect 40040 50448 40092 50454
rect 40040 50390 40092 50396
rect 27620 40724 27672 40730
rect 27620 40666 27672 40672
rect 26240 32428 26292 32434
rect 26240 32370 26292 32376
rect 19352 16546 20208 16574
rect 20732 16546 21864 16574
rect 24872 16546 25360 16574
rect 19430 3360 19486 3369
rect 19430 3295 19486 3304
rect 19444 480 19472 3295
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20180 354 20208 16546
rect 21836 480 21864 16546
rect 23020 7676 23072 7682
rect 23020 7618 23072 7624
rect 23032 480 23060 7618
rect 24216 3460 24268 3466
rect 24216 3402 24268 3408
rect 24228 480 24256 3402
rect 25332 480 25360 16546
rect 20598 354 20710 480
rect 20180 326 20710 354
rect 20598 -960 20710 326
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 32370
rect 27632 16574 27660 40666
rect 34520 29640 34572 29646
rect 34520 29582 34572 29588
rect 29000 25628 29052 25634
rect 29000 25570 29052 25576
rect 29012 16574 29040 25570
rect 33140 19984 33192 19990
rect 33140 19926 33192 19932
rect 33152 16574 33180 19926
rect 27632 16546 27752 16574
rect 29012 16546 30144 16574
rect 33152 16546 33640 16574
rect 27724 480 27752 16546
rect 28908 3528 28960 3534
rect 28908 3470 28960 3476
rect 28920 480 28948 3470
rect 30116 480 30144 16546
rect 31300 7744 31352 7750
rect 31300 7686 31352 7692
rect 31312 480 31340 7686
rect 32404 3664 32456 3670
rect 32404 3606 32456 3612
rect 32416 480 32444 3606
rect 33612 480 33640 16546
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34532 354 34560 29582
rect 35900 21412 35952 21418
rect 35900 21354 35952 21360
rect 35912 16574 35940 21354
rect 40052 16574 40080 50390
rect 41420 31068 41472 31074
rect 41420 31010 41472 31016
rect 41432 16574 41460 31010
rect 44192 16574 44220 51682
rect 46940 43444 46992 43450
rect 46940 43386 46992 43392
rect 46952 16574 46980 43386
rect 48332 16574 48360 55830
rect 49712 16574 49740 58618
rect 52460 49020 52512 49026
rect 52460 48962 52512 48968
rect 51080 33856 51132 33862
rect 51080 33798 51132 33804
rect 35912 16546 36768 16574
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 44192 16546 44312 16574
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 35992 3800 36044 3806
rect 35992 3742 36044 3748
rect 36004 480 36032 3742
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 38384 7812 38436 7818
rect 38384 7754 38436 7760
rect 38396 480 38424 7754
rect 39580 3936 39632 3942
rect 39580 3878 39632 3884
rect 39592 480 39620 3878
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40236 354 40264 16546
rect 41892 480 41920 16546
rect 43076 4072 43128 4078
rect 43076 4014 43128 4020
rect 43088 480 43116 4014
rect 44284 480 44312 16546
rect 45468 7880 45520 7886
rect 45468 7822 45520 7828
rect 45480 480 45508 7822
rect 46664 3392 46716 3398
rect 46664 3334 46716 3340
rect 46676 480 46704 3334
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51092 354 51120 33798
rect 52472 6914 52500 48962
rect 52552 39364 52604 39370
rect 52552 39306 52604 39312
rect 52564 16574 52592 39306
rect 53852 16574 53880 58686
rect 57980 53100 58032 53106
rect 57980 53042 58032 53048
rect 57992 16574 58020 53042
rect 52564 16546 53328 16574
rect 53852 16546 54984 16574
rect 57992 16546 58480 16574
rect 52472 6886 52592 6914
rect 52564 480 52592 6886
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53300 354 53328 16546
rect 54956 480 54984 16546
rect 56784 11756 56836 11762
rect 56784 11698 56836 11704
rect 56048 6316 56100 6322
rect 56048 6258 56100 6264
rect 56060 480 56088 6258
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 11698
rect 58452 480 58480 16546
rect 60832 13116 60884 13122
rect 60832 13058 60884 13064
rect 59636 6384 59688 6390
rect 59636 6326 59688 6332
rect 59648 480 59676 6326
rect 60844 480 60872 13058
rect 61396 3738 61424 59463
rect 62762 59392 62818 59401
rect 62762 59327 62818 59336
rect 62120 44872 62172 44878
rect 62120 44814 62172 44820
rect 62132 16574 62160 44814
rect 62132 16546 62712 16574
rect 62028 8968 62080 8974
rect 62028 8910 62080 8916
rect 61384 3732 61436 3738
rect 61384 3674 61436 3680
rect 62040 480 62068 8910
rect 62684 3482 62712 16546
rect 62776 3602 62804 59327
rect 63500 17332 63552 17338
rect 63500 17274 63552 17280
rect 63512 16574 63540 17274
rect 63512 16546 64368 16574
rect 62764 3596 62816 3602
rect 62764 3538 62816 3544
rect 62684 3454 63264 3482
rect 63236 480 63264 3454
rect 64340 480 64368 16546
rect 64524 3602 64552 59463
rect 65996 59401 66024 59758
rect 70582 59800 70638 59809
rect 66442 59735 66498 59744
rect 70136 59758 70582 59786
rect 67546 59664 67602 59673
rect 67546 59599 67602 59608
rect 64694 59392 64750 59401
rect 64694 59327 64750 59336
rect 65982 59392 66038 59401
rect 65982 59327 66038 59336
rect 66166 59392 66222 59401
rect 66166 59327 66222 59336
rect 64708 3738 64736 59327
rect 65064 10328 65116 10334
rect 65064 10270 65116 10276
rect 64696 3732 64748 3738
rect 64696 3674 64748 3680
rect 64512 3596 64564 3602
rect 64512 3538 64564 3544
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 10270
rect 66180 3874 66208 59327
rect 66720 14476 66772 14482
rect 66720 14418 66772 14424
rect 66168 3868 66220 3874
rect 66168 3810 66220 3816
rect 66732 480 66760 14418
rect 67560 4010 67588 59599
rect 68650 59528 68706 59537
rect 68650 59463 68706 59472
rect 67640 18624 67692 18630
rect 67640 18566 67692 18572
rect 67548 4004 67600 4010
rect 67548 3946 67600 3952
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 18566
rect 68664 4146 68692 59463
rect 70136 59401 70164 59758
rect 70582 59735 70638 59744
rect 71594 59800 71650 59809
rect 74722 59800 74778 59809
rect 71594 59735 71650 59744
rect 73068 59764 73120 59770
rect 71608 59401 71636 59735
rect 79874 59800 79930 59809
rect 74722 59735 74724 59744
rect 73068 59706 73120 59712
rect 74776 59735 74778 59744
rect 77944 59764 77996 59770
rect 74724 59706 74776 59712
rect 83002 59800 83058 59809
rect 79874 59735 79876 59744
rect 77944 59706 77996 59712
rect 79928 59735 79930 59744
rect 80704 59764 80756 59770
rect 79876 59706 79928 59712
rect 87418 59800 87474 59809
rect 83002 59735 83004 59744
rect 80704 59706 80756 59712
rect 83056 59735 83058 59744
rect 86224 59764 86276 59770
rect 83004 59706 83056 59712
rect 87418 59735 87420 59744
rect 86224 59706 86276 59712
rect 87472 59735 87474 59744
rect 94502 59800 94558 59809
rect 94502 59735 94558 59744
rect 97170 59800 97226 59809
rect 97538 59800 97594 59809
rect 97226 59758 97538 59786
rect 97170 59735 97226 59744
rect 97538 59735 97594 59744
rect 98458 59800 98514 59809
rect 98458 59735 98514 59744
rect 104806 59800 104862 59809
rect 108210 59800 108266 59809
rect 104806 59735 104862 59744
rect 107948 59758 108210 59786
rect 87420 59706 87472 59712
rect 71686 59664 71742 59673
rect 71686 59599 71742 59608
rect 68834 59392 68890 59401
rect 68834 59327 68890 59336
rect 70122 59392 70178 59401
rect 70122 59327 70178 59336
rect 70306 59392 70362 59401
rect 70306 59327 70362 59336
rect 71594 59392 71650 59401
rect 71594 59327 71650 59336
rect 68652 4140 68704 4146
rect 68652 4082 68704 4088
rect 68848 3330 68876 59327
rect 70320 6914 70348 59327
rect 71700 11830 71728 59599
rect 72882 59528 72938 59537
rect 72882 59463 72938 59472
rect 72896 17270 72924 59463
rect 72884 17264 72936 17270
rect 72884 17206 72936 17212
rect 73080 13190 73108 59706
rect 75826 59664 75882 59673
rect 75826 59599 75882 59608
rect 74446 59392 74502 59401
rect 74446 59327 74502 59336
rect 74460 24138 74488 59327
rect 74448 24132 74500 24138
rect 74448 24074 74500 24080
rect 73344 15904 73396 15910
rect 73344 15846 73396 15852
rect 73068 13184 73120 13190
rect 73068 13126 73120 13132
rect 71688 11824 71740 11830
rect 71688 11766 71740 11772
rect 70228 6886 70348 6914
rect 69112 4956 69164 4962
rect 69112 4898 69164 4904
rect 68836 3324 68888 3330
rect 68836 3266 68888 3272
rect 69124 480 69152 4898
rect 70228 3262 70256 6886
rect 70308 6452 70360 6458
rect 70308 6394 70360 6400
rect 70216 3256 70268 3262
rect 70216 3198 70268 3204
rect 70320 480 70348 6394
rect 71504 5228 71556 5234
rect 71504 5170 71556 5176
rect 71516 480 71544 5170
rect 72608 5024 72660 5030
rect 72608 4966 72660 4972
rect 72620 480 72648 4966
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 15846
rect 75840 6526 75868 59599
rect 77206 59528 77262 59537
rect 77206 59463 77262 59472
rect 77022 59392 77078 59401
rect 77022 59327 77078 59336
rect 77036 9654 77064 59327
rect 77024 9648 77076 9654
rect 77024 9590 77076 9596
rect 75828 6520 75880 6526
rect 75828 6462 75880 6468
rect 77220 5574 77248 59463
rect 77300 22772 77352 22778
rect 77300 22714 77352 22720
rect 77312 16574 77340 22714
rect 77312 16546 77432 16574
rect 77208 5568 77260 5574
rect 77208 5510 77260 5516
rect 76196 5092 76248 5098
rect 76196 5034 76248 5040
rect 75000 4208 75052 4214
rect 75000 4150 75052 4156
rect 75012 480 75040 4150
rect 76208 480 76236 5034
rect 77404 480 77432 16546
rect 77956 4214 77984 59706
rect 79874 59664 79930 59673
rect 79874 59599 79930 59608
rect 79888 51074 79916 59599
rect 79336 51046 79916 51074
rect 78588 9648 78640 9654
rect 78588 9590 78640 9596
rect 77944 4208 77996 4214
rect 77944 4150 77996 4156
rect 78600 480 78628 9590
rect 79336 5234 79364 51046
rect 80060 42084 80112 42090
rect 80060 42026 80112 42032
rect 80072 16574 80100 42026
rect 80716 17338 80744 59706
rect 80886 59528 80942 59537
rect 80886 59463 80942 59472
rect 83462 59528 83518 59537
rect 83462 59463 83518 59472
rect 80900 18630 80928 59463
rect 82082 59392 82138 59401
rect 82082 59327 82138 59336
rect 80888 18624 80940 18630
rect 80888 18566 80940 18572
rect 80704 17332 80756 17338
rect 80704 17274 80756 17280
rect 80072 16546 80928 16574
rect 79324 5228 79376 5234
rect 79324 5170 79376 5176
rect 79692 5160 79744 5166
rect 79692 5102 79744 5108
rect 79704 480 79732 5102
rect 80900 480 80928 16546
rect 82096 13122 82124 59327
rect 82084 13116 82136 13122
rect 82084 13058 82136 13064
rect 83476 11762 83504 59463
rect 84842 59392 84898 59401
rect 84842 59327 84898 59336
rect 84856 39370 84884 59327
rect 85486 59256 85542 59265
rect 85486 59191 85542 59200
rect 85500 58682 85528 59191
rect 85488 58676 85540 58682
rect 85488 58618 85540 58624
rect 84844 39364 84896 39370
rect 84844 39306 84896 39312
rect 83464 11756 83516 11762
rect 83464 11698 83516 11704
rect 84476 9036 84528 9042
rect 84476 8978 84528 8984
rect 82084 5568 82136 5574
rect 82084 5510 82136 5516
rect 82096 480 82124 5510
rect 83280 5228 83332 5234
rect 83280 5170 83332 5176
rect 83292 480 83320 5170
rect 84488 480 84516 8978
rect 85672 6520 85724 6526
rect 85672 6462 85724 6468
rect 85684 480 85712 6462
rect 86236 3398 86264 59706
rect 87602 59664 87658 59673
rect 91282 59664 91338 59673
rect 87602 59599 87658 59608
rect 89168 59628 89220 59634
rect 86960 18624 87012 18630
rect 86960 18566 87012 18572
rect 86972 16574 87000 18566
rect 86972 16546 87552 16574
rect 86868 5296 86920 5302
rect 86868 5238 86920 5244
rect 86224 3392 86276 3398
rect 86224 3334 86276 3340
rect 86880 480 86908 5238
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87524 354 87552 16546
rect 87616 4078 87644 59599
rect 93306 59664 93362 59673
rect 91282 59599 91284 59608
rect 89168 59570 89220 59576
rect 91336 59599 91338 59608
rect 92952 59622 93306 59650
rect 91284 59570 91336 59576
rect 88982 59528 89038 59537
rect 88982 59463 89038 59472
rect 88340 24132 88392 24138
rect 88340 24074 88392 24080
rect 88352 16574 88380 24074
rect 88352 16546 88932 16574
rect 87604 4072 87656 4078
rect 87604 4014 87656 4020
rect 88904 3482 88932 16546
rect 88996 3942 89024 59463
rect 89180 16574 89208 59570
rect 92952 59401 92980 59622
rect 93306 59599 93362 59608
rect 94318 59664 94374 59673
rect 94318 59599 94374 59608
rect 93306 59528 93362 59537
rect 93306 59463 93362 59472
rect 90362 59392 90418 59401
rect 90362 59327 90418 59336
rect 91742 59392 91798 59401
rect 91742 59327 91798 59336
rect 92938 59392 92994 59401
rect 92938 59327 92994 59336
rect 93122 59392 93178 59401
rect 93122 59327 93178 59336
rect 89180 16546 89300 16574
rect 88984 3936 89036 3942
rect 88984 3878 89036 3884
rect 89272 3806 89300 16546
rect 89904 11756 89956 11762
rect 89904 11698 89956 11704
rect 89260 3800 89312 3806
rect 89260 3742 89312 3748
rect 88904 3454 89208 3482
rect 89180 480 89208 3454
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 11698
rect 90376 3670 90404 59327
rect 91560 10396 91612 10402
rect 91560 10338 91612 10344
rect 90364 3664 90416 3670
rect 90364 3606 90416 3612
rect 91572 480 91600 10338
rect 91756 3534 91784 59327
rect 92480 13184 92532 13190
rect 92480 13126 92532 13132
rect 91744 3528 91796 3534
rect 91744 3470 91796 3476
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 13126
rect 93136 3369 93164 59327
rect 93320 3466 93348 59463
rect 94332 59401 94360 59599
rect 94516 59537 94544 59735
rect 97814 59664 97870 59673
rect 97814 59599 97870 59608
rect 94502 59528 94558 59537
rect 94502 59463 94558 59472
rect 95882 59528 95938 59537
rect 95882 59463 95938 59472
rect 97630 59528 97686 59537
rect 97630 59463 97686 59472
rect 94318 59392 94374 59401
rect 94318 59327 94374 59336
rect 94502 59392 94558 59401
rect 94502 59327 94558 59336
rect 93860 47660 93912 47666
rect 93860 47602 93912 47608
rect 93872 16574 93900 47602
rect 93872 16546 93992 16574
rect 93308 3460 93360 3466
rect 93308 3402 93360 3408
rect 93122 3360 93178 3369
rect 93122 3295 93178 3304
rect 93964 480 93992 16546
rect 94412 13184 94464 13190
rect 94412 13126 94464 13132
rect 94424 490 94452 13126
rect 94516 6254 94544 59327
rect 95896 47598 95924 59463
rect 95884 47592 95936 47598
rect 95884 47534 95936 47540
rect 95240 17264 95292 17270
rect 95240 17206 95292 17212
rect 95252 16574 95280 17206
rect 95252 16546 95832 16574
rect 94504 6248 94556 6254
rect 94504 6190 94556 6196
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94424 462 94820 490
rect 94792 354 94820 462
rect 95118 354 95230 480
rect 94792 326 95230 354
rect 95804 354 95832 16546
rect 97448 13116 97500 13122
rect 97448 13058 97500 13064
rect 97460 480 97488 13058
rect 97644 3466 97672 59463
rect 97828 3534 97856 59599
rect 98472 59537 98500 59735
rect 104714 59664 104770 59673
rect 104714 59599 104770 59608
rect 98458 59528 98514 59537
rect 102598 59528 102654 59537
rect 98458 59463 98514 59472
rect 102060 59486 102598 59514
rect 99286 59392 99342 59401
rect 99286 59327 99342 59336
rect 101956 59356 102008 59362
rect 98000 23860 98052 23866
rect 98000 23802 98052 23808
rect 98012 16574 98040 23802
rect 98012 16546 98224 16574
rect 97816 3528 97868 3534
rect 97816 3470 97868 3476
rect 97632 3460 97684 3466
rect 97632 3402 97684 3408
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99300 3670 99328 59327
rect 101956 59298 102008 59304
rect 100666 59256 100722 59265
rect 100666 59191 100722 59200
rect 99840 11824 99892 11830
rect 99840 11766 99892 11772
rect 99288 3664 99340 3670
rect 99288 3606 99340 3612
rect 99852 480 99880 11766
rect 100680 3806 100708 59191
rect 100760 17264 100812 17270
rect 100760 17206 100812 17212
rect 100668 3800 100720 3806
rect 100668 3742 100720 3748
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 17206
rect 101968 14550 101996 59298
rect 101956 14544 102008 14550
rect 101956 14486 102008 14492
rect 102060 11830 102088 59486
rect 102598 59463 102654 59472
rect 102230 59392 102286 59401
rect 102230 59327 102286 59336
rect 103426 59392 103482 59401
rect 103426 59327 103428 59336
rect 102048 11824 102100 11830
rect 102048 11766 102100 11772
rect 102244 480 102272 59327
rect 103480 59327 103482 59336
rect 103428 59298 103480 59304
rect 103520 55956 103572 55962
rect 103520 55898 103572 55904
rect 103532 16574 103560 55898
rect 104728 45554 104756 59599
rect 104820 59401 104848 59735
rect 105726 59528 105782 59537
rect 105726 59463 105782 59472
rect 104806 59392 104862 59401
rect 104806 59327 104862 59336
rect 105542 59392 105598 59401
rect 105542 59327 105598 59336
rect 104176 45526 104756 45554
rect 104176 23866 104204 45526
rect 104164 23860 104216 23866
rect 104164 23802 104216 23808
rect 103532 16546 104112 16574
rect 103336 3256 103388 3262
rect 103336 3198 103388 3204
rect 103348 480 103376 3198
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105556 10402 105584 59327
rect 105636 14544 105688 14550
rect 105636 14486 105688 14492
rect 105544 10396 105596 10402
rect 105544 10338 105596 10344
rect 105648 6914 105676 14486
rect 105740 13190 105768 59463
rect 107948 59401 107976 59758
rect 108210 59735 108266 59744
rect 112534 59800 112590 59809
rect 120262 59800 120318 59809
rect 112534 59735 112590 59744
rect 118608 59764 118660 59770
rect 108302 59664 108358 59673
rect 108302 59599 108358 59608
rect 110878 59664 110934 59673
rect 110878 59599 110934 59608
rect 112442 59664 112498 59673
rect 112442 59599 112498 59608
rect 106922 59392 106978 59401
rect 106922 59327 106978 59336
rect 107934 59392 107990 59401
rect 107934 59327 107990 59336
rect 106936 18630 106964 59327
rect 106924 18624 106976 18630
rect 106924 18566 106976 18572
rect 107660 18624 107712 18630
rect 107660 18566 107712 18572
rect 107672 16574 107700 18566
rect 107672 16546 108160 16574
rect 105728 13184 105780 13190
rect 105728 13126 105780 13132
rect 105648 6886 105768 6914
rect 105740 480 105768 6886
rect 106924 3324 106976 3330
rect 106924 3266 106976 3272
rect 106936 480 106964 3266
rect 108132 480 108160 16546
rect 108316 9042 108344 59599
rect 109682 59528 109738 59537
rect 109682 59463 109738 59472
rect 109696 22778 109724 59463
rect 110892 58682 110920 59599
rect 111062 59392 111118 59401
rect 111062 59327 111118 59336
rect 109868 58676 109920 58682
rect 109868 58618 109920 58624
rect 110880 58676 110932 58682
rect 110880 58618 110932 58624
rect 109880 42090 109908 58618
rect 110512 49088 110564 49094
rect 110512 49030 110564 49036
rect 109868 42084 109920 42090
rect 109868 42026 109920 42032
rect 109684 22772 109736 22778
rect 109684 22714 109736 22720
rect 109040 11824 109092 11830
rect 109040 11766 109092 11772
rect 108304 9036 108356 9042
rect 108304 8978 108356 8984
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109052 354 109080 11766
rect 110524 6914 110552 49030
rect 111076 15910 111104 59327
rect 111064 15904 111116 15910
rect 111064 15846 111116 15852
rect 110524 6886 111656 6914
rect 110512 4140 110564 4146
rect 110512 4082 110564 4088
rect 110524 480 110552 4082
rect 111628 480 111656 6886
rect 112456 6458 112484 59599
rect 112548 59401 112576 59735
rect 120262 59735 120264 59744
rect 118608 59706 118660 59712
rect 120316 59735 120318 59744
rect 121274 59800 121330 59809
rect 128450 59800 128506 59809
rect 121274 59735 121330 59744
rect 128096 59758 128450 59786
rect 120264 59706 120316 59712
rect 118146 59664 118202 59673
rect 116584 59628 116636 59634
rect 118146 59599 118148 59608
rect 116584 59570 116636 59576
rect 118200 59599 118202 59608
rect 118148 59570 118200 59576
rect 113822 59528 113878 59537
rect 116122 59528 116178 59537
rect 113822 59463 113878 59472
rect 114008 59492 114060 59498
rect 112534 59392 112590 59401
rect 112534 59327 112590 59336
rect 113836 14482 113864 59463
rect 116122 59463 116124 59472
rect 114008 59434 114060 59440
rect 116176 59463 116178 59472
rect 116124 59434 116176 59440
rect 114020 44878 114048 59434
rect 115202 59392 115258 59401
rect 115202 59327 115258 59336
rect 114008 44872 114060 44878
rect 114008 44814 114060 44820
rect 114744 15904 114796 15910
rect 114744 15846 114796 15852
rect 113824 14476 113876 14482
rect 113824 14418 113876 14424
rect 112444 6452 112496 6458
rect 112444 6394 112496 6400
rect 114008 4004 114060 4010
rect 114008 3946 114060 3952
rect 112812 3800 112864 3806
rect 112812 3742 112864 3748
rect 112824 480 112852 3742
rect 114020 480 114048 3946
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 114756 354 114784 15846
rect 115216 6390 115244 59327
rect 115204 6384 115256 6390
rect 115204 6326 115256 6332
rect 116596 6322 116624 59570
rect 118146 59528 118202 59537
rect 118146 59463 118202 59472
rect 118160 51074 118188 59463
rect 118620 55894 118648 59706
rect 120906 59664 120962 59673
rect 120906 59599 120962 59608
rect 119342 59392 119398 59401
rect 119342 59327 119398 59336
rect 120722 59392 120778 59401
rect 120722 59327 120778 59336
rect 118608 55888 118660 55894
rect 118608 55830 118660 55836
rect 117976 51046 118188 51074
rect 117976 49026 118004 51046
rect 117964 49020 118016 49026
rect 117964 48962 118016 48968
rect 119356 7886 119384 59327
rect 119344 7880 119396 7886
rect 119344 7822 119396 7828
rect 120736 7818 120764 59327
rect 120920 31074 120948 59599
rect 121288 59537 121316 59735
rect 125414 59664 125470 59673
rect 123484 59628 123536 59634
rect 125414 59599 125416 59608
rect 123484 59570 123536 59576
rect 125468 59599 125470 59608
rect 125416 59570 125468 59576
rect 121274 59528 121330 59537
rect 121274 59463 121330 59472
rect 122102 59392 122158 59401
rect 122102 59327 122158 59336
rect 122838 59392 122894 59401
rect 122838 59327 122894 59336
rect 120908 31068 120960 31074
rect 120908 31010 120960 31016
rect 122116 29646 122144 59327
rect 122852 59242 122880 59327
rect 123114 59256 123170 59265
rect 122852 59214 123114 59242
rect 123114 59191 123170 59200
rect 122104 29640 122156 29646
rect 122104 29582 122156 29588
rect 120724 7812 120776 7818
rect 120724 7754 120776 7760
rect 123496 7750 123524 59570
rect 128096 59537 128124 59758
rect 131578 59800 131634 59809
rect 128450 59735 128506 59744
rect 129004 59764 129056 59770
rect 137834 59800 137890 59809
rect 131578 59735 131580 59744
rect 129004 59706 129056 59712
rect 131632 59735 131634 59744
rect 131764 59764 131816 59770
rect 131580 59706 131632 59712
rect 131764 59706 131816 59712
rect 132592 59764 132644 59770
rect 132592 59706 132644 59712
rect 136548 59764 136600 59770
rect 137834 59735 137836 59744
rect 136548 59706 136600 59712
rect 137888 59735 137890 59744
rect 138938 59800 138994 59809
rect 141974 59800 142030 59809
rect 138938 59735 138994 59744
rect 140044 59764 140096 59770
rect 137836 59706 137888 59712
rect 125414 59528 125470 59537
rect 125414 59463 125470 59472
rect 128082 59528 128138 59537
rect 128082 59463 128138 59472
rect 124862 59256 124918 59265
rect 124862 59191 124918 59200
rect 123484 7744 123536 7750
rect 123484 7686 123536 7692
rect 124876 7682 124904 59191
rect 125428 45554 125456 59463
rect 126242 59392 126298 59401
rect 126242 59327 126298 59336
rect 125060 45526 125456 45554
rect 125060 40730 125088 45526
rect 125048 40724 125100 40730
rect 125048 40666 125100 40672
rect 126256 26926 126284 59327
rect 127714 59256 127770 59265
rect 127714 59191 127770 59200
rect 127728 45554 127756 59191
rect 127636 45526 127756 45554
rect 126980 31136 127032 31142
rect 126980 31078 127032 31084
rect 126244 26920 126296 26926
rect 126244 26862 126296 26868
rect 125600 22772 125652 22778
rect 125600 22714 125652 22720
rect 124864 7676 124916 7682
rect 124864 7618 124916 7624
rect 116584 6316 116636 6322
rect 116584 6258 116636 6264
rect 117596 3868 117648 3874
rect 117596 3810 117648 3816
rect 116400 3664 116452 3670
rect 116400 3606 116452 3612
rect 116412 480 116440 3606
rect 117608 480 117636 3810
rect 121092 3732 121144 3738
rect 121092 3674 121144 3680
rect 118792 3664 118844 3670
rect 118792 3606 118844 3612
rect 118804 480 118832 3606
rect 119896 3528 119948 3534
rect 119896 3470 119948 3476
rect 119908 480 119936 3470
rect 121104 480 121132 3674
rect 124680 3596 124732 3602
rect 124680 3538 124732 3544
rect 122288 3528 122340 3534
rect 122288 3470 122340 3476
rect 122300 480 122328 3470
rect 123484 3460 123536 3466
rect 123484 3402 123536 3408
rect 123496 480 123524 3402
rect 124692 480 124720 3538
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125612 354 125640 22714
rect 126992 480 127020 31078
rect 127636 7614 127664 45526
rect 128360 44872 128412 44878
rect 128360 44814 128412 44820
rect 128372 16574 128400 44814
rect 128372 16546 128952 16574
rect 128176 14476 128228 14482
rect 128176 14418 128228 14424
rect 127624 7608 127676 7614
rect 127624 7550 127676 7556
rect 128188 480 128216 14418
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 129016 4894 129044 59706
rect 129186 59528 129242 59537
rect 129186 59463 129242 59472
rect 129200 6186 129228 59463
rect 130382 59392 130438 59401
rect 130382 59327 130438 59336
rect 129740 42152 129792 42158
rect 129740 42094 129792 42100
rect 129752 16574 129780 42094
rect 129752 16546 130332 16574
rect 129188 6180 129240 6186
rect 129188 6122 129240 6128
rect 129004 4888 129056 4894
rect 129004 4830 129056 4836
rect 130304 3482 130332 16546
rect 130396 3602 130424 59327
rect 131120 40860 131172 40866
rect 131120 40802 131172 40808
rect 131132 16574 131160 40802
rect 131132 16546 131344 16574
rect 130384 3596 130436 3602
rect 130384 3538 130436 3544
rect 130304 3454 130608 3482
rect 130580 480 130608 3454
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 131776 3670 131804 59706
rect 132604 59673 132632 59706
rect 132590 59664 132646 59673
rect 132590 59599 132646 59608
rect 133142 59528 133198 59537
rect 133142 59463 133198 59472
rect 133156 15910 133184 59463
rect 133326 59392 133382 59401
rect 133326 59327 133382 59336
rect 133340 49094 133368 59327
rect 134522 59256 134578 59265
rect 134522 59191 134578 59200
rect 133880 51876 133932 51882
rect 133880 51818 133932 51824
rect 133328 49088 133380 49094
rect 133328 49030 133380 49036
rect 133144 15904 133196 15910
rect 133144 15846 133196 15852
rect 132960 7608 133012 7614
rect 132960 7550 133012 7556
rect 131764 3664 131816 3670
rect 131764 3606 131816 3612
rect 132972 480 133000 7550
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 133892 354 133920 51818
rect 134536 18630 134564 59191
rect 136560 55962 136588 59706
rect 137834 59664 137890 59673
rect 137834 59599 137890 59608
rect 137466 59528 137522 59537
rect 137466 59463 137522 59472
rect 137282 59392 137338 59401
rect 137282 59327 137338 59336
rect 136548 55956 136600 55962
rect 136548 55898 136600 55904
rect 135260 55888 135312 55894
rect 135260 55830 135312 55836
rect 134524 18624 134576 18630
rect 134524 18566 134576 18572
rect 135272 3602 135300 55830
rect 136640 36644 136692 36650
rect 136640 36586 136692 36592
rect 135352 26988 135404 26994
rect 135352 26930 135404 26936
rect 135260 3596 135312 3602
rect 135260 3538 135312 3544
rect 135364 3482 135392 26930
rect 136652 16574 136680 36586
rect 136652 16546 137232 16574
rect 136456 3596 136508 3602
rect 136456 3538 136508 3544
rect 135272 3454 135392 3482
rect 135272 480 135300 3454
rect 136468 480 136496 3538
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 137296 13122 137324 59327
rect 137480 17270 137508 59463
rect 137848 59401 137876 59599
rect 138952 59537 138980 59735
rect 145010 59800 145066 59809
rect 141974 59735 141976 59744
rect 140044 59706 140096 59712
rect 142028 59735 142030 59744
rect 142804 59764 142856 59770
rect 141976 59706 142028 59712
rect 148138 59800 148194 59809
rect 145010 59735 145012 59744
rect 142804 59706 142856 59712
rect 145064 59735 145066 59744
rect 145748 59764 145800 59770
rect 145012 59706 145064 59712
rect 148138 59735 148140 59744
rect 145748 59706 145800 59712
rect 148192 59735 148194 59744
rect 150254 59800 150310 59809
rect 152278 59800 152334 59809
rect 150254 59735 150310 59744
rect 150348 59764 150400 59770
rect 148140 59706 148192 59712
rect 138938 59528 138994 59537
rect 138938 59463 138994 59472
rect 137834 59392 137890 59401
rect 137834 59327 137890 59336
rect 138662 59392 138718 59401
rect 138662 59327 138718 59336
rect 138676 47666 138704 59327
rect 139400 50380 139452 50386
rect 139400 50322 139452 50328
rect 138664 47660 138716 47666
rect 138664 47602 138716 47608
rect 138020 45076 138072 45082
rect 138020 45018 138072 45024
rect 137468 17264 137520 17270
rect 137468 17206 137520 17212
rect 138032 16574 138060 45018
rect 139412 16574 139440 50322
rect 138032 16546 138888 16574
rect 139412 16546 139624 16574
rect 137284 13116 137336 13122
rect 137284 13058 137336 13064
rect 138860 480 138888 16546
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 140056 11762 140084 59706
rect 141422 59528 141478 59537
rect 141422 59463 141478 59472
rect 140780 53236 140832 53242
rect 140780 53178 140832 53184
rect 140792 16574 140820 53178
rect 140792 16546 141280 16574
rect 140044 11756 140096 11762
rect 140044 11698 140096 11704
rect 141252 480 141280 16546
rect 141436 5302 141464 59463
rect 141606 59392 141662 59401
rect 141606 59327 141662 59336
rect 141424 5296 141476 5302
rect 141424 5238 141476 5244
rect 141620 5234 141648 59327
rect 142160 11688 142212 11694
rect 142160 11630 142212 11636
rect 141608 5228 141660 5234
rect 141608 5170 141660 5176
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142172 354 142200 11630
rect 142816 5166 142844 59706
rect 145562 59528 145618 59537
rect 145562 59463 145618 59472
rect 144182 59256 144238 59265
rect 144182 59191 144238 59200
rect 143540 49088 143592 49094
rect 143540 49030 143592 49036
rect 143552 11762 143580 49030
rect 143632 47592 143684 47598
rect 143632 47534 143684 47540
rect 143540 11756 143592 11762
rect 143540 11698 143592 11704
rect 143644 6914 143672 47534
rect 143552 6886 143672 6914
rect 142804 5160 142856 5166
rect 142804 5102 142856 5108
rect 143552 480 143580 6886
rect 144196 5098 144224 59191
rect 144920 22840 144972 22846
rect 144920 22782 144972 22788
rect 144932 16574 144960 22782
rect 144932 16546 145512 16574
rect 144736 11756 144788 11762
rect 144736 11698 144788 11704
rect 144184 5092 144236 5098
rect 144184 5034 144236 5040
rect 144748 480 144776 11698
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 145576 5030 145604 59463
rect 145564 5024 145616 5030
rect 145564 4966 145616 4972
rect 145760 4962 145788 59706
rect 149702 59664 149758 59673
rect 149702 59599 149758 59608
rect 148322 59528 148378 59537
rect 148322 59463 148378 59472
rect 146942 59392 146998 59401
rect 146942 59327 146998 59336
rect 146300 58676 146352 58682
rect 146300 58618 146352 58624
rect 146312 6914 146340 58618
rect 146956 10334 146984 59327
rect 147864 15904 147916 15910
rect 147864 15846 147916 15852
rect 146944 10328 146996 10334
rect 146944 10270 146996 10276
rect 146312 6886 147168 6914
rect 145748 4956 145800 4962
rect 145748 4898 145800 4904
rect 147140 480 147168 6886
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 15846
rect 148336 8974 148364 59463
rect 149716 53106 149744 59599
rect 150268 59537 150296 59735
rect 156602 59800 156658 59809
rect 152278 59735 152280 59744
rect 150348 59706 150400 59712
rect 152332 59735 152334 59744
rect 153844 59764 153896 59770
rect 152280 59706 152332 59712
rect 156602 59735 156604 59744
rect 153844 59706 153896 59712
rect 156656 59735 156658 59744
rect 157430 59800 157486 59809
rect 157430 59735 157486 59744
rect 159546 59800 159602 59809
rect 162582 59800 162638 59809
rect 159546 59735 159602 59744
rect 160744 59764 160796 59770
rect 156604 59706 156656 59712
rect 150254 59528 150310 59537
rect 150254 59463 150310 59472
rect 150360 58750 150388 59706
rect 151082 59392 151138 59401
rect 151082 59327 151138 59336
rect 150348 58744 150400 58750
rect 150348 58686 150400 58692
rect 149704 53100 149756 53106
rect 149704 53042 149756 53048
rect 151096 33862 151124 59327
rect 152462 59256 152518 59265
rect 152462 59191 152518 59200
rect 151820 49156 151872 49162
rect 151820 49098 151872 49104
rect 151084 33856 151136 33862
rect 151084 33798 151136 33804
rect 150440 33788 150492 33794
rect 150440 33730 150492 33736
rect 149060 31272 149112 31278
rect 149060 31214 149112 31220
rect 149072 16574 149100 31214
rect 150452 16574 150480 33730
rect 149072 16546 149560 16574
rect 150452 16546 150664 16574
rect 148324 8968 148376 8974
rect 148324 8910 148376 8916
rect 149532 480 149560 16546
rect 150636 480 150664 16546
rect 151832 9674 151860 49098
rect 152476 43450 152504 59191
rect 153856 50454 153884 59706
rect 154302 59664 154358 59673
rect 154302 59599 154358 59608
rect 156602 59664 156658 59673
rect 156602 59599 156658 59608
rect 154026 59528 154082 59537
rect 154026 59463 154082 59472
rect 154040 51746 154068 59463
rect 154316 59401 154344 59599
rect 154302 59392 154358 59401
rect 154302 59327 154358 59336
rect 155222 59392 155278 59401
rect 155222 59327 155278 59336
rect 154028 51740 154080 51746
rect 154028 51682 154080 51688
rect 153844 50448 153896 50454
rect 153844 50390 153896 50396
rect 152464 43444 152516 43450
rect 152464 43386 152516 43392
rect 151912 39432 151964 39438
rect 151912 39374 151964 39380
rect 151740 9654 151860 9674
rect 151728 9648 151860 9654
rect 151780 9646 151860 9648
rect 151728 9590 151780 9596
rect 151924 6914 151952 39374
rect 153200 35216 153252 35222
rect 153200 35158 153252 35164
rect 153212 16574 153240 35158
rect 155236 21418 155264 59327
rect 155224 21412 155276 21418
rect 155224 21354 155276 21360
rect 156616 19990 156644 59599
rect 157444 59401 157472 59735
rect 158626 59664 158682 59673
rect 158626 59599 158682 59608
rect 157982 59528 158038 59537
rect 157982 59463 158038 59472
rect 157430 59392 157486 59401
rect 157430 59327 157486 59336
rect 157996 25634 158024 59463
rect 158640 45554 158668 59599
rect 159560 59537 159588 59735
rect 162582 59735 162584 59744
rect 160744 59706 160796 59712
rect 162636 59735 162638 59744
rect 165710 59800 165766 59809
rect 165710 59735 165766 59744
rect 170954 59800 171010 59809
rect 170954 59735 171010 59744
rect 178222 59800 178278 59809
rect 181258 59800 181314 59809
rect 178222 59735 178278 59744
rect 179236 59764 179288 59770
rect 162584 59706 162636 59712
rect 159546 59528 159602 59537
rect 159546 59463 159602 59472
rect 159362 59392 159418 59401
rect 159362 59327 159418 59336
rect 158180 45526 158668 45554
rect 158180 32434 158208 45526
rect 158720 38004 158772 38010
rect 158720 37946 158772 37952
rect 158168 32428 158220 32434
rect 158168 32370 158220 32376
rect 157984 25628 158036 25634
rect 157984 25570 158036 25576
rect 157340 25560 157392 25566
rect 157340 25502 157392 25508
rect 156604 19984 156656 19990
rect 156604 19926 156656 19932
rect 154580 17264 154632 17270
rect 154580 17206 154632 17212
rect 154592 16574 154620 17206
rect 157352 16574 157380 25502
rect 158732 16574 158760 37946
rect 159376 37942 159404 59327
rect 159364 37936 159416 37942
rect 159364 37878 159416 37884
rect 160756 28286 160784 59706
rect 164882 59664 164938 59673
rect 164882 59599 164938 59608
rect 162582 59528 162638 59537
rect 162136 59486 162582 59514
rect 161480 57316 161532 57322
rect 161480 57258 161532 57264
rect 160744 28280 160796 28286
rect 160744 28222 160796 28228
rect 160100 26920 160152 26926
rect 160100 26862 160152 26868
rect 153212 16546 153792 16574
rect 154592 16546 155448 16574
rect 157352 16546 157840 16574
rect 158732 16546 158944 16574
rect 153016 9648 153068 9654
rect 153016 9590 153068 9596
rect 151832 6886 151952 6914
rect 151832 480 151860 6886
rect 153028 480 153056 9590
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16546
rect 155420 480 155448 16546
rect 156144 13116 156196 13122
rect 156144 13058 156196 13064
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156156 354 156184 13058
rect 157812 480 157840 16546
rect 158916 480 158944 16546
rect 160112 3534 160140 26862
rect 161492 16574 161520 57258
rect 161492 16546 162072 16574
rect 160100 3528 160152 3534
rect 160100 3470 160152 3476
rect 161296 3528 161348 3534
rect 161296 3470 161348 3476
rect 160100 3256 160152 3262
rect 160100 3198 160152 3204
rect 160112 480 160140 3198
rect 161308 480 161336 3470
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 16546
rect 162136 4826 162164 59486
rect 162582 59463 162638 59472
rect 162582 59392 162638 59401
rect 162582 59327 162638 59336
rect 162596 54534 162624 59327
rect 164146 59256 164202 59265
rect 164146 59191 164202 59200
rect 164160 57254 164188 59191
rect 164148 57248 164200 57254
rect 164148 57190 164200 57196
rect 162860 54664 162912 54670
rect 162860 54606 162912 54612
rect 162584 54528 162636 54534
rect 162584 54470 162636 54476
rect 162872 16574 162900 54606
rect 164896 46238 164924 59599
rect 165724 59401 165752 59735
rect 170862 59664 170918 59673
rect 170862 59599 170918 59608
rect 166814 59528 166870 59537
rect 166814 59463 166870 59472
rect 165710 59392 165766 59401
rect 165710 59327 165766 59336
rect 166630 59392 166686 59401
rect 166630 59327 166686 59336
rect 164884 46232 164936 46238
rect 164884 46174 164936 46180
rect 164240 32428 164292 32434
rect 164240 32370 164292 32376
rect 164252 16574 164280 32370
rect 165620 29776 165672 29782
rect 165620 29718 165672 29724
rect 165632 16574 165660 29718
rect 162872 16546 163728 16574
rect 164252 16546 164464 16574
rect 165632 16546 166120 16574
rect 162124 4820 162176 4826
rect 162124 4762 162176 4768
rect 163700 480 163728 16546
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164436 354 164464 16546
rect 166092 480 166120 16546
rect 166644 3466 166672 59327
rect 166632 3460 166684 3466
rect 166632 3402 166684 3408
rect 166828 3369 166856 59463
rect 168286 59256 168342 59265
rect 168286 59191 168342 59200
rect 167184 14544 167236 14550
rect 167184 14486 167236 14492
rect 166814 3360 166870 3369
rect 166814 3295 166870 3304
rect 167196 480 167224 14486
rect 168300 3670 168328 59191
rect 168380 55956 168432 55962
rect 168380 55898 168432 55904
rect 168288 3664 168340 3670
rect 168288 3606 168340 3612
rect 168392 3602 168420 55898
rect 168472 54528 168524 54534
rect 168472 54470 168524 54476
rect 168380 3596 168432 3602
rect 168380 3538 168432 3544
rect 168484 3482 168512 54470
rect 170876 45554 170904 59599
rect 170784 45526 170904 45554
rect 170784 20058 170812 45526
rect 170772 20052 170824 20058
rect 170772 19994 170824 20000
rect 170968 19990 170996 59735
rect 178130 59664 178186 59673
rect 177960 59622 178130 59650
rect 177118 59528 177174 59537
rect 175096 59492 175148 59498
rect 177118 59463 177120 59472
rect 175096 59434 175148 59440
rect 177172 59463 177174 59472
rect 177120 59434 177172 59440
rect 172426 59392 172482 59401
rect 172426 59327 172482 59336
rect 171140 36576 171192 36582
rect 171140 36518 171192 36524
rect 170956 19984 171008 19990
rect 170956 19926 171008 19932
rect 169760 17332 169812 17338
rect 169760 17274 169812 17280
rect 169772 16574 169800 17274
rect 171152 16574 171180 36518
rect 172440 20126 172468 59327
rect 173806 59256 173862 59265
rect 173806 59191 173862 59200
rect 173820 43450 173848 59191
rect 174910 59120 174966 59129
rect 174910 59055 174966 59064
rect 173808 43444 173860 43450
rect 173808 43386 173860 43392
rect 172520 28416 172572 28422
rect 172520 28358 172572 28364
rect 172428 20120 172480 20126
rect 172428 20062 172480 20068
rect 172532 16574 172560 28358
rect 174924 20194 174952 59055
rect 175108 20262 175136 59434
rect 176566 59392 176622 59401
rect 176566 59327 176622 59336
rect 175280 37936 175332 37942
rect 175280 37878 175332 37884
rect 175096 20256 175148 20262
rect 175096 20198 175148 20204
rect 174912 20188 174964 20194
rect 174912 20130 174964 20136
rect 175292 16574 175320 37878
rect 176580 20330 176608 59327
rect 177960 25634 177988 59622
rect 178130 59599 178186 59608
rect 178236 59401 178264 59735
rect 190550 59800 190606 59809
rect 181258 59735 181260 59744
rect 179236 59706 179288 59712
rect 181312 59735 181314 59744
rect 188896 59764 188948 59770
rect 181260 59706 181312 59712
rect 195794 59800 195850 59809
rect 190550 59735 190552 59744
rect 188896 59706 188948 59712
rect 190604 59735 190606 59744
rect 194508 59764 194560 59770
rect 190552 59706 190604 59712
rect 195794 59735 195796 59744
rect 194508 59706 194560 59712
rect 195848 59735 195850 59744
rect 196806 59800 196862 59809
rect 196806 59735 196862 59744
rect 198830 59800 198886 59809
rect 208122 59800 208178 59809
rect 198830 59735 198886 59744
rect 206928 59764 206980 59770
rect 195796 59706 195848 59712
rect 179142 59528 179198 59537
rect 179142 59463 179198 59472
rect 178222 59392 178278 59401
rect 178222 59327 178278 59336
rect 179156 45554 179184 59463
rect 179248 50454 179276 59706
rect 182086 59664 182142 59673
rect 182086 59599 182142 59608
rect 180706 59392 180762 59401
rect 180706 59327 180762 59336
rect 179236 50448 179288 50454
rect 179236 50390 179288 50396
rect 179064 45526 179184 45554
rect 178040 39364 178092 39370
rect 178040 39306 178092 39312
rect 177948 25628 178000 25634
rect 177948 25570 178000 25576
rect 176660 24268 176712 24274
rect 176660 24210 176712 24216
rect 176568 20324 176620 20330
rect 176568 20266 176620 20272
rect 169772 16546 170352 16574
rect 171152 16546 172008 16574
rect 172532 16546 172744 16574
rect 175292 16546 175504 16574
rect 169576 3596 169628 3602
rect 169576 3538 169628 3544
rect 168392 3454 168512 3482
rect 168392 480 168420 3454
rect 169588 480 169616 3538
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 16546
rect 171980 480 172008 16546
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 174268 9104 174320 9110
rect 174268 9046 174320 9052
rect 174280 480 174308 9046
rect 175476 480 175504 16546
rect 176672 480 176700 24210
rect 178052 16574 178080 39306
rect 179064 31074 179092 45526
rect 179420 35352 179472 35358
rect 179420 35294 179472 35300
rect 179052 31068 179104 31074
rect 179052 31010 179104 31016
rect 179432 16574 179460 35294
rect 180720 33862 180748 59327
rect 180708 33856 180760 33862
rect 180708 33798 180760 33804
rect 182100 28286 182128 59599
rect 183190 59528 183246 59537
rect 183190 59463 183246 59472
rect 187422 59528 187478 59537
rect 187422 59463 187478 59472
rect 182180 40724 182232 40730
rect 182180 40666 182232 40672
rect 182088 28280 182140 28286
rect 182088 28222 182140 28228
rect 178052 16546 178632 16574
rect 179432 16546 180288 16574
rect 177856 9172 177908 9178
rect 177856 9114 177908 9120
rect 177868 480 177896 9114
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173134 -960 173246 326
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 180260 480 180288 16546
rect 181444 9240 181496 9246
rect 181444 9182 181496 9188
rect 181456 480 181484 9182
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182192 354 182220 40666
rect 183204 29646 183232 59463
rect 183466 59392 183522 59401
rect 183466 59327 183522 59336
rect 183480 53174 183508 59327
rect 184846 59256 184902 59265
rect 184846 59191 184902 59200
rect 183468 53168 183520 53174
rect 183468 53110 183520 53116
rect 183192 29640 183244 29646
rect 183192 29582 183244 29588
rect 184860 24206 184888 59191
rect 187436 45554 187464 59463
rect 187514 59392 187570 59401
rect 187514 59327 187570 59336
rect 187344 45526 187464 45554
rect 184940 32496 184992 32502
rect 184940 32438 184992 32444
rect 184848 24200 184900 24206
rect 184848 24142 184900 24148
rect 183744 4820 183796 4826
rect 183744 4762 183796 4768
rect 183756 480 183784 4762
rect 184952 480 184980 32438
rect 185032 24132 185084 24138
rect 185032 24074 185084 24080
rect 185044 16574 185072 24074
rect 187344 18630 187372 45526
rect 187528 18698 187556 59327
rect 188908 51814 188936 59706
rect 188986 59664 189042 59673
rect 190550 59664 190606 59673
rect 188986 59599 189042 59608
rect 190380 59622 190550 59650
rect 189000 58750 189028 59599
rect 188988 58744 189040 58750
rect 188988 58686 189040 58692
rect 188896 51808 188948 51814
rect 188896 51750 188948 51756
rect 189080 42084 189132 42090
rect 189080 42026 189132 42032
rect 187700 27260 187752 27266
rect 187700 27202 187752 27208
rect 187516 18692 187568 18698
rect 187516 18634 187568 18640
rect 187332 18624 187384 18630
rect 187332 18566 187384 18572
rect 187712 16574 187740 27202
rect 189092 16574 189120 42026
rect 190380 18766 190408 59622
rect 190550 59599 190606 59608
rect 191470 59528 191526 59537
rect 193678 59528 193734 59537
rect 191470 59463 191526 59472
rect 191748 59492 191800 59498
rect 190460 33992 190512 33998
rect 190460 33934 190512 33940
rect 190368 18760 190420 18766
rect 190368 18702 190420 18708
rect 185044 16546 186176 16574
rect 187712 16546 188568 16574
rect 189092 16546 189304 16574
rect 186148 480 186176 16546
rect 187332 4888 187384 4894
rect 187332 4830 187384 4836
rect 187344 480 187372 4830
rect 188540 480 188568 16546
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189276 354 189304 16546
rect 189694 354 189806 480
rect 189276 326 189806 354
rect 190472 354 190500 33934
rect 191484 18834 191512 59463
rect 193678 59463 193680 59472
rect 191748 59434 191800 59440
rect 193732 59463 193734 59472
rect 193680 59434 193732 59440
rect 191760 45554 191788 59434
rect 193126 59392 193182 59401
rect 193126 59327 193182 59336
rect 191668 45526 191788 45554
rect 191668 18902 191696 45526
rect 193140 18970 193168 59327
rect 193220 45008 193272 45014
rect 193220 44950 193272 44956
rect 193128 18964 193180 18970
rect 193128 18906 193180 18912
rect 191656 18896 191708 18902
rect 191656 18838 191708 18844
rect 191472 18828 191524 18834
rect 191472 18770 191524 18776
rect 192024 9036 192076 9042
rect 192024 8978 192076 8984
rect 192036 480 192064 8978
rect 193232 3670 193260 44950
rect 193312 43512 193364 43518
rect 193312 43454 193364 43460
rect 193220 3664 193272 3670
rect 193220 3606 193272 3612
rect 193324 3482 193352 43454
rect 194520 19038 194548 59706
rect 195794 59664 195850 59673
rect 195794 59599 195850 59608
rect 195702 59528 195758 59537
rect 195702 59463 195758 59472
rect 195716 51074 195744 59463
rect 195624 51046 195744 51074
rect 194600 23112 194652 23118
rect 194600 23054 194652 23060
rect 194508 19032 194560 19038
rect 194508 18974 194560 18980
rect 194612 16574 194640 23054
rect 195624 19106 195652 51046
rect 195808 19174 195836 59599
rect 196820 59537 196848 59735
rect 196806 59528 196862 59537
rect 196806 59463 196862 59472
rect 198646 59528 198702 59537
rect 198646 59463 198702 59472
rect 197266 59392 197322 59401
rect 197266 59327 197322 59336
rect 195980 46232 196032 46238
rect 195980 46174 196032 46180
rect 195796 19168 195848 19174
rect 195796 19110 195848 19116
rect 195612 19100 195664 19106
rect 195612 19042 195664 19048
rect 195992 16574 196020 46174
rect 197280 42226 197308 59327
rect 198660 46306 198688 59463
rect 198844 59401 198872 59735
rect 208122 59735 208124 59744
rect 206928 59706 206980 59712
rect 208176 59735 208178 59744
rect 209962 59800 210018 59809
rect 210330 59800 210386 59809
rect 210018 59758 210330 59786
rect 209962 59735 210018 59744
rect 210330 59735 210386 59744
rect 211250 59800 211306 59809
rect 222566 59800 222622 59809
rect 211250 59735 211306 59744
rect 220452 59764 220504 59770
rect 208124 59706 208176 59712
rect 200026 59664 200082 59673
rect 200026 59599 200082 59608
rect 199842 59528 199898 59537
rect 199842 59463 199898 59472
rect 198830 59392 198886 59401
rect 198830 59327 198886 59336
rect 198648 46300 198700 46306
rect 198648 46242 198700 46248
rect 199856 45554 199884 59463
rect 200040 51074 200068 59599
rect 206098 59528 206154 59537
rect 203892 59492 203944 59498
rect 206098 59463 206100 59472
rect 203892 59434 203944 59440
rect 206152 59463 206154 59472
rect 206100 59434 206152 59440
rect 201406 59392 201462 59401
rect 201406 59327 201462 59336
rect 200120 53100 200172 53106
rect 200120 53042 200172 53048
rect 199764 45526 199884 45554
rect 199948 51046 200068 51074
rect 197268 42220 197320 42226
rect 197268 42162 197320 42168
rect 194612 16546 195192 16574
rect 195992 16546 196848 16574
rect 194416 3664 194468 3670
rect 194416 3606 194468 3612
rect 193232 3454 193352 3482
rect 193232 480 193260 3454
rect 194428 480 194456 3606
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 189694 -960 189806 326
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 196820 480 196848 16546
rect 198740 14612 198792 14618
rect 198740 14554 198792 14560
rect 197912 5092 197964 5098
rect 197912 5034 197964 5040
rect 197924 480 197952 5034
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 14554
rect 199764 3670 199792 45526
rect 199752 3664 199804 3670
rect 199752 3606 199804 3612
rect 199948 3534 199976 51046
rect 200132 16574 200160 53042
rect 200132 16546 200344 16574
rect 199936 3528 199988 3534
rect 199936 3470 199988 3476
rect 200316 480 200344 16546
rect 201420 3738 201448 59327
rect 202786 59256 202842 59265
rect 202786 59191 202842 59200
rect 201500 47728 201552 47734
rect 201500 47670 201552 47676
rect 201408 3732 201460 3738
rect 201408 3674 201460 3680
rect 201512 3398 201540 47670
rect 201592 5024 201644 5030
rect 201592 4966 201644 4972
rect 201500 3392 201552 3398
rect 201500 3334 201552 3340
rect 201604 2530 201632 4966
rect 202800 3806 202828 59191
rect 202880 25696 202932 25702
rect 202880 25638 202932 25644
rect 202892 16574 202920 25638
rect 202892 16546 203472 16574
rect 202788 3800 202840 3806
rect 202788 3742 202840 3748
rect 202696 3392 202748 3398
rect 202696 3334 202748 3340
rect 201512 2502 201632 2530
rect 201512 480 201540 2502
rect 202708 480 202736 3334
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 16546
rect 203904 3942 203932 59434
rect 205546 59392 205602 59401
rect 205546 59327 205602 59336
rect 204074 59256 204130 59265
rect 204074 59191 204130 59200
rect 203892 3936 203944 3942
rect 203892 3878 203944 3884
rect 204088 3874 204116 59191
rect 204260 57384 204312 57390
rect 204260 57326 204312 57332
rect 204272 16574 204300 57326
rect 204272 16546 205128 16574
rect 204076 3868 204128 3874
rect 204076 3810 204128 3816
rect 205100 480 205128 16546
rect 205560 4010 205588 59327
rect 206192 8968 206244 8974
rect 206192 8910 206244 8916
rect 205548 4004 205600 4010
rect 205548 3946 205600 3952
rect 206204 480 206232 8910
rect 206940 4078 206968 59706
rect 208214 59664 208270 59673
rect 208214 59599 208270 59608
rect 211066 59664 211122 59673
rect 211066 59599 211122 59608
rect 208122 59528 208178 59537
rect 208122 59463 208178 59472
rect 207020 47660 207072 47666
rect 207020 47602 207072 47608
rect 206928 4072 206980 4078
rect 206928 4014 206980 4020
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 47602
rect 208136 45554 208164 59463
rect 208044 45526 208164 45554
rect 208044 4146 208072 45526
rect 208032 4140 208084 4146
rect 208032 4082 208084 4088
rect 208228 3398 208256 59599
rect 209686 59392 209742 59401
rect 209686 59327 209742 59336
rect 208400 46368 208452 46374
rect 208400 46310 208452 46316
rect 208412 16574 208440 46310
rect 208412 16546 208624 16574
rect 208216 3392 208268 3398
rect 208216 3334 208268 3340
rect 208596 480 208624 16546
rect 209700 3330 209728 59327
rect 209780 49020 209832 49026
rect 209780 48962 209832 48968
rect 209792 4214 209820 48962
rect 211080 44946 211108 59599
rect 211264 59401 211292 59735
rect 222566 59735 222568 59744
rect 220452 59706 220504 59712
rect 222620 59735 222622 59744
rect 223670 59800 223726 59809
rect 223670 59735 223726 59744
rect 227902 59800 227958 59809
rect 227902 59735 227958 59744
rect 238758 59800 238814 59809
rect 244278 59800 244334 59809
rect 238758 59735 238814 59744
rect 242808 59764 242860 59770
rect 222568 59706 222620 59712
rect 217966 59664 218022 59673
rect 217966 59599 218022 59608
rect 219898 59664 219954 59673
rect 219898 59599 219954 59608
rect 212262 59528 212318 59537
rect 212262 59463 212318 59472
rect 216402 59528 216458 59537
rect 216402 59463 216458 59472
rect 211250 59392 211306 59401
rect 211250 59327 211306 59336
rect 212276 51074 212304 59463
rect 212354 59392 212410 59401
rect 212354 59327 212410 59336
rect 212184 51046 212304 51074
rect 211068 44940 211120 44946
rect 211068 44882 211120 44888
rect 212184 21418 212212 51046
rect 212368 21486 212396 59327
rect 213826 59256 213882 59265
rect 213826 59191 213882 59200
rect 212540 32564 212592 32570
rect 212540 32506 212592 32512
rect 212356 21480 212408 21486
rect 212356 21422 212408 21428
rect 212172 21412 212224 21418
rect 212172 21354 212224 21360
rect 209872 17468 209924 17474
rect 209872 17410 209924 17416
rect 209780 4208 209832 4214
rect 209780 4150 209832 4156
rect 209884 3482 209912 17410
rect 212552 16574 212580 32506
rect 213840 21554 213868 59191
rect 213920 51740 213972 51746
rect 213920 51682 213972 51688
rect 213828 21548 213880 21554
rect 213828 21490 213880 21496
rect 213932 16574 213960 51682
rect 216416 45554 216444 59463
rect 216494 59392 216550 59401
rect 216494 59327 216550 59336
rect 216508 54738 216536 59327
rect 217874 59256 217930 59265
rect 217874 59191 217930 59200
rect 217888 55214 217916 59191
rect 217980 58954 218008 59599
rect 219346 59528 219402 59537
rect 219346 59463 219402 59472
rect 217968 58948 218020 58954
rect 217968 58890 218020 58896
rect 217888 55186 218008 55214
rect 216496 54732 216548 54738
rect 216496 54674 216548 54680
rect 216324 45526 216444 45554
rect 215300 40792 215352 40798
rect 215300 40734 215352 40740
rect 212552 16546 213408 16574
rect 213932 16546 214512 16574
rect 212172 5092 212224 5098
rect 212172 5034 212224 5040
rect 210976 4208 211028 4214
rect 210976 4150 211028 4156
rect 209792 3454 209912 3482
rect 209688 3324 209740 3330
rect 209688 3266 209740 3272
rect 209792 480 209820 3454
rect 210988 480 211016 4150
rect 212184 480 212212 5034
rect 213380 480 213408 16546
rect 214484 480 214512 16546
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 40734
rect 216324 21622 216352 45526
rect 217980 27130 218008 55186
rect 218060 50516 218112 50522
rect 218060 50458 218112 50464
rect 217968 27124 218020 27130
rect 217968 27066 218020 27072
rect 216312 21616 216364 21622
rect 216312 21558 216364 21564
rect 216864 9308 216916 9314
rect 216864 9250 216916 9256
rect 216876 480 216904 9250
rect 218072 480 218100 50458
rect 219360 47802 219388 59463
rect 219912 59401 219940 59599
rect 219898 59392 219954 59401
rect 219898 59327 219954 59336
rect 219348 47796 219400 47802
rect 219348 47738 219400 47744
rect 220464 21690 220492 59706
rect 223486 59664 223542 59673
rect 223486 59599 223542 59608
rect 220634 59392 220690 59401
rect 220634 59327 220690 59336
rect 220648 38214 220676 59327
rect 222106 59256 222162 59265
rect 222106 59191 222162 59200
rect 222120 46510 222148 59191
rect 222108 46504 222160 46510
rect 222108 46446 222160 46452
rect 220636 38208 220688 38214
rect 220636 38150 220688 38156
rect 220820 28348 220872 28354
rect 220820 28290 220872 28296
rect 220452 21684 220504 21690
rect 220452 21626 220504 21632
rect 220832 16574 220860 28290
rect 223500 22982 223528 59599
rect 223684 59401 223712 59735
rect 227810 59664 227866 59673
rect 227640 59622 227810 59650
rect 224682 59528 224738 59537
rect 226706 59528 226762 59537
rect 224682 59463 224738 59472
rect 224868 59492 224920 59498
rect 223670 59392 223726 59401
rect 223670 59327 223726 59336
rect 224696 39642 224724 59463
rect 226706 59463 226708 59472
rect 224868 59434 224920 59440
rect 226760 59463 226762 59472
rect 226708 59434 226760 59440
rect 224684 39636 224736 39642
rect 224684 39578 224736 39584
rect 224880 32638 224908 59434
rect 226246 59392 226302 59401
rect 226246 59327 226302 59336
rect 226260 42430 226288 59327
rect 226248 42424 226300 42430
rect 226248 42366 226300 42372
rect 224868 32632 224920 32638
rect 224868 32574 224920 32580
rect 224960 29708 225012 29714
rect 224960 29650 225012 29656
rect 223488 22976 223540 22982
rect 223488 22918 223540 22924
rect 224972 16574 225000 29650
rect 227640 20398 227668 59622
rect 227810 59599 227866 59608
rect 227916 59401 227944 59735
rect 232962 59664 233018 59673
rect 232962 59599 233018 59608
rect 229006 59528 229062 59537
rect 229006 59463 229062 59472
rect 232870 59528 232926 59537
rect 232870 59463 232926 59472
rect 227902 59392 227958 59401
rect 227902 59327 227958 59336
rect 228822 59392 228878 59401
rect 228822 59327 228878 59336
rect 228836 45554 228864 59327
rect 229020 56030 229048 59463
rect 230386 59392 230442 59401
rect 230386 59327 230442 59336
rect 231766 59392 231822 59401
rect 231766 59327 231822 59336
rect 229008 56024 229060 56030
rect 229008 55966 229060 55972
rect 228744 45526 228864 45554
rect 228744 20466 228772 45526
rect 230400 36854 230428 59327
rect 230388 36848 230440 36854
rect 230388 36790 230440 36796
rect 231780 35426 231808 59327
rect 231768 35420 231820 35426
rect 231768 35362 231820 35368
rect 228732 20460 228784 20466
rect 228732 20402 228784 20408
rect 227628 20392 227680 20398
rect 227628 20334 227680 20340
rect 220832 16546 221136 16574
rect 224972 16546 225184 16574
rect 219992 10328 220044 10334
rect 219992 10270 220044 10276
rect 219256 6180 219308 6186
rect 219256 6122 219308 6128
rect 219268 480 219296 6122
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 10270
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 16546
rect 223580 10396 223632 10402
rect 223580 10338 223632 10344
rect 222752 6248 222804 6254
rect 222752 6190 222804 6196
rect 222764 480 222792 6190
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 10338
rect 225156 480 225184 16546
rect 232884 15978 232912 59463
rect 232976 59401 233004 59599
rect 238772 59537 238800 59735
rect 244278 59735 244280 59744
rect 242808 59706 242860 59712
rect 244332 59735 244334 59744
rect 246762 59800 246818 59809
rect 246762 59735 246818 59744
rect 248418 59800 248474 59809
rect 248418 59735 248474 59744
rect 252650 59800 252706 59809
rect 259826 59800 259882 59809
rect 252650 59735 252706 59744
rect 257896 59764 257948 59770
rect 244280 59706 244332 59712
rect 242714 59664 242770 59673
rect 242714 59599 242770 59608
rect 234986 59528 235042 59537
rect 233056 59492 233108 59498
rect 234986 59463 234988 59472
rect 233056 59434 233108 59440
rect 235040 59463 235042 59472
rect 238758 59528 238814 59537
rect 238758 59463 238814 59472
rect 241334 59528 241390 59537
rect 241334 59463 241390 59472
rect 234988 59434 235040 59440
rect 232962 59392 233018 59401
rect 232962 59327 233018 59336
rect 233068 54806 233096 59434
rect 234526 59392 234582 59401
rect 234526 59327 234582 59336
rect 238666 59392 238722 59401
rect 238666 59327 238722 59336
rect 241242 59392 241298 59401
rect 241242 59327 241298 59336
rect 233056 54800 233108 54806
rect 233056 54742 233108 54748
rect 233240 43716 233292 43722
rect 233240 43658 233292 43664
rect 233252 16574 233280 43658
rect 233252 16546 233464 16574
rect 232872 15972 232924 15978
rect 232872 15914 232924 15920
rect 226340 10532 226392 10538
rect 226340 10474 226392 10480
rect 226352 3194 226380 10474
rect 231032 9376 231084 9382
rect 231032 9318 231084 9324
rect 228732 7676 228784 7682
rect 228732 7618 228784 7624
rect 226432 6316 226484 6322
rect 226432 6258 226484 6264
rect 226340 3188 226392 3194
rect 226340 3130 226392 3136
rect 226444 2122 226472 6258
rect 227536 3188 227588 3194
rect 227536 3130 227588 3136
rect 226352 2094 226472 2122
rect 226352 480 226380 2094
rect 227548 480 227576 3130
rect 228744 480 228772 7618
rect 229836 6384 229888 6390
rect 229836 6326 229888 6332
rect 229848 480 229876 6326
rect 231044 480 231072 9318
rect 232228 7744 232280 7750
rect 232228 7686 232280 7692
rect 232240 480 232268 7686
rect 233436 480 233464 16546
rect 234540 16046 234568 59327
rect 235906 59256 235962 59265
rect 235906 59191 235962 59200
rect 237194 59256 237250 59265
rect 237194 59191 237250 59200
rect 234528 16040 234580 16046
rect 234528 15982 234580 15988
rect 234620 10600 234672 10606
rect 234620 10542 234672 10548
rect 234632 480 234660 10542
rect 235920 10470 235948 59191
rect 237010 59120 237066 59129
rect 237010 59055 237066 59064
rect 236000 25764 236052 25770
rect 236000 25706 236052 25712
rect 236012 16574 236040 25706
rect 236012 16546 236592 16574
rect 235908 10464 235960 10470
rect 235908 10406 235960 10412
rect 235816 7812 235868 7818
rect 235816 7754 235868 7760
rect 235828 480 235856 7754
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 237024 16114 237052 59055
rect 237208 16182 237236 59191
rect 238680 16250 238708 59327
rect 241256 45554 241284 59327
rect 241164 45526 241284 45554
rect 241164 17406 241192 45526
rect 241348 41002 241376 59463
rect 242728 57526 242756 59599
rect 242716 57520 242768 57526
rect 242716 57462 242768 57468
rect 241336 40996 241388 41002
rect 241336 40938 241388 40944
rect 241152 17400 241204 17406
rect 241152 17342 241204 17348
rect 238668 16244 238720 16250
rect 238668 16186 238720 16192
rect 237196 16176 237248 16182
rect 237196 16118 237248 16124
rect 237012 16108 237064 16114
rect 237012 16050 237064 16056
rect 242820 13190 242848 59706
rect 245474 59664 245530 59673
rect 245474 59599 245530 59608
rect 244186 59528 244242 59537
rect 244186 59463 244242 59472
rect 244200 45150 244228 59463
rect 245292 58404 245344 58410
rect 245292 58346 245344 58352
rect 244188 45144 244240 45150
rect 244188 45086 244240 45092
rect 242900 31204 242952 31210
rect 242900 31146 242952 31152
rect 242808 13184 242860 13190
rect 242808 13126 242860 13132
rect 237656 10668 237708 10674
rect 237656 10610 237708 10616
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 10610
rect 241704 9444 241756 9450
rect 241704 9386 241756 9392
rect 239312 7880 239364 7886
rect 239312 7822 239364 7828
rect 239324 480 239352 7822
rect 240508 6452 240560 6458
rect 240508 6394 240560 6400
rect 240520 480 240548 6394
rect 241716 480 241744 9386
rect 242912 480 242940 31146
rect 245304 13394 245332 58346
rect 245292 13388 245344 13394
rect 245292 13330 245344 13336
rect 245488 13258 245516 59599
rect 246776 58410 246804 59735
rect 248326 59528 248382 59537
rect 248326 59463 248382 59472
rect 246948 58608 247000 58614
rect 246948 58550 247000 58556
rect 246764 58404 246816 58410
rect 246764 58346 246816 58352
rect 246960 13462 246988 58550
rect 248340 13530 248368 59463
rect 248432 58614 248460 59735
rect 252558 59664 252614 59673
rect 252480 59622 252558 59650
rect 249430 59528 249486 59537
rect 251546 59528 251602 59537
rect 249430 59463 249486 59472
rect 249708 59492 249760 59498
rect 248420 58608 248472 58614
rect 248420 58550 248472 58556
rect 248420 56092 248472 56098
rect 248420 56034 248472 56040
rect 248328 13524 248380 13530
rect 248328 13466 248380 13472
rect 246948 13456 247000 13462
rect 246948 13398 247000 13404
rect 245476 13252 245528 13258
rect 245476 13194 245528 13200
rect 245200 10736 245252 10742
rect 245200 10678 245252 10684
rect 244096 6520 244148 6526
rect 244096 6462 244148 6468
rect 244108 480 244136 6462
rect 245212 480 245240 10678
rect 246396 7948 246448 7954
rect 246396 7890 246448 7896
rect 246408 480 246436 7890
rect 247592 6588 247644 6594
rect 247592 6530 247644 6536
rect 247604 480 247632 6530
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248432 354 248460 56034
rect 249444 14686 249472 59463
rect 251546 59463 251548 59472
rect 249708 59434 249760 59440
rect 251600 59463 251602 59472
rect 251548 59434 251600 59440
rect 249720 45554 249748 59434
rect 251086 59392 251142 59401
rect 251086 59327 251142 59336
rect 249628 45526 249748 45554
rect 249628 36718 249656 45526
rect 249616 36712 249668 36718
rect 249616 36654 249668 36660
rect 251100 17542 251128 59327
rect 251180 57452 251232 57458
rect 251180 57394 251232 57400
rect 251088 17536 251140 17542
rect 251088 17478 251140 17484
rect 249432 14680 249484 14686
rect 249432 14622 249484 14628
rect 249984 8016 250036 8022
rect 249984 7958 250036 7964
rect 249996 480 250024 7958
rect 251192 4214 251220 57394
rect 251272 39704 251324 39710
rect 251272 39646 251324 39652
rect 251180 4208 251232 4214
rect 251180 4150 251232 4156
rect 251284 3482 251312 39646
rect 252480 11898 252508 59622
rect 252558 59599 252614 59608
rect 252664 59401 252692 59735
rect 259826 59735 259828 59744
rect 257896 59706 257948 59712
rect 259880 59735 259882 59744
rect 263966 59800 264022 59809
rect 263966 59735 264022 59744
rect 266174 59800 266230 59809
rect 268106 59800 268162 59809
rect 266174 59735 266230 59744
rect 266268 59764 266320 59770
rect 259828 59706 259880 59712
rect 253662 59528 253718 59537
rect 255686 59528 255742 59537
rect 253662 59463 253718 59472
rect 253756 59492 253808 59498
rect 252650 59392 252706 59401
rect 252650 59327 252706 59336
rect 253676 51074 253704 59463
rect 257802 59528 257858 59537
rect 255686 59463 255688 59472
rect 253756 59434 253808 59440
rect 255740 59463 255742 59472
rect 256608 59492 256660 59498
rect 255688 59434 255740 59440
rect 257802 59463 257804 59472
rect 256608 59434 256660 59440
rect 257856 59463 257858 59472
rect 257804 59434 257856 59440
rect 253584 51046 253704 51074
rect 252560 33924 252612 33930
rect 252560 33866 252612 33872
rect 252572 16574 252600 33866
rect 252572 16546 253520 16574
rect 252468 11892 252520 11898
rect 252468 11834 252520 11840
rect 252376 4208 252428 4214
rect 252376 4150 252428 4156
rect 251192 3454 251312 3482
rect 251192 480 251220 3454
rect 252388 480 252416 4150
rect 253492 480 253520 16546
rect 253584 11966 253612 51046
rect 253768 12034 253796 59434
rect 255226 59392 255282 59401
rect 255226 59327 255282 59336
rect 253940 38276 253992 38282
rect 253940 38218 253992 38224
rect 253952 16574 253980 38218
rect 253952 16546 254256 16574
rect 253756 12028 253808 12034
rect 253756 11970 253808 11976
rect 253572 11960 253624 11966
rect 253572 11902 253624 11908
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 255240 12102 255268 59327
rect 255228 12096 255280 12102
rect 255228 12038 255280 12044
rect 256620 11830 256648 59434
rect 257802 59392 257858 59401
rect 257802 59327 257858 59336
rect 257816 45554 257844 59327
rect 257724 45526 257844 45554
rect 256700 35284 256752 35290
rect 256700 35226 256752 35232
rect 256608 11824 256660 11830
rect 256608 11766 256660 11772
rect 255872 9512 255924 9518
rect 255872 9454 255924 9460
rect 255884 480 255912 9454
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 256712 354 256740 35226
rect 257724 12170 257752 45526
rect 257908 12238 257936 59706
rect 260746 59528 260802 59537
rect 260746 59463 260802 59472
rect 259366 59256 259422 59265
rect 259366 59191 259422 59200
rect 258080 49292 258132 49298
rect 258080 49234 258132 49240
rect 258092 16574 258120 49234
rect 258092 16546 258304 16574
rect 257896 12232 257948 12238
rect 257896 12174 257948 12180
rect 257712 12164 257764 12170
rect 257712 12106 257764 12112
rect 258276 480 258304 16546
rect 259380 12306 259408 59191
rect 259460 58812 259512 58818
rect 259460 58754 259512 58760
rect 259368 12300 259420 12306
rect 259368 12242 259420 12248
rect 259472 11694 259500 58754
rect 260760 14754 260788 59463
rect 261942 59392 261998 59401
rect 263980 59362 264008 59735
rect 266082 59664 266138 59673
rect 266082 59599 266138 59608
rect 264242 59528 264298 59537
rect 264242 59463 264298 59472
rect 261942 59327 261998 59336
rect 262220 59356 262272 59362
rect 261956 55010 261984 59327
rect 262220 59298 262272 59304
rect 263968 59356 264020 59362
rect 263968 59298 264020 59304
rect 261944 55004 261996 55010
rect 261944 54946 261996 54952
rect 260840 29912 260892 29918
rect 260840 29854 260892 29860
rect 260852 16574 260880 29854
rect 262232 16574 262260 59298
rect 262862 59256 262918 59265
rect 262862 59191 262918 59200
rect 260852 16546 261800 16574
rect 262232 16546 262536 16574
rect 260748 14748 260800 14754
rect 260748 14690 260800 14696
rect 259460 11688 259512 11694
rect 259460 11630 259512 11636
rect 260656 11688 260708 11694
rect 260656 11630 260708 11636
rect 259460 11008 259512 11014
rect 259460 10950 259512 10956
rect 259472 480 259500 10950
rect 260668 480 260696 11630
rect 261772 480 261800 16546
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 262876 11014 262904 59191
rect 263600 57248 263652 57254
rect 263600 57190 263652 57196
rect 263612 16574 263640 57190
rect 263612 16546 264192 16574
rect 262864 11008 262916 11014
rect 262864 10950 262916 10956
rect 264164 480 264192 16546
rect 264256 9518 264284 59463
rect 266096 57458 266124 59599
rect 266188 59537 266216 59735
rect 272522 59800 272578 59809
rect 268106 59735 268108 59744
rect 266268 59706 266320 59712
rect 268160 59735 268162 59744
rect 272260 59758 272522 59786
rect 268108 59706 268160 59712
rect 266174 59528 266230 59537
rect 266174 59463 266230 59472
rect 266084 57452 266136 57458
rect 266084 57394 266136 57400
rect 266280 56098 266308 59706
rect 270222 59664 270278 59673
rect 270222 59599 270278 59608
rect 269946 59528 270002 59537
rect 269946 59463 270002 59472
rect 267002 59392 267058 59401
rect 267002 59327 267058 59336
rect 266268 56092 266320 56098
rect 266268 56034 266320 56040
rect 266360 55004 266412 55010
rect 266360 54946 266412 54952
rect 264980 23044 265032 23050
rect 264980 22986 265032 22992
rect 264244 9512 264296 9518
rect 264244 9454 264296 9460
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 264992 354 265020 22986
rect 266372 16574 266400 54946
rect 266372 16546 266584 16574
rect 266556 480 266584 16546
rect 267016 10742 267044 59327
rect 268382 59256 268438 59265
rect 268382 59191 268438 59200
rect 269762 59256 269818 59265
rect 269762 59191 269818 59200
rect 267740 56160 267792 56166
rect 267740 56102 267792 56108
rect 267004 10736 267056 10742
rect 267004 10678 267056 10684
rect 267752 4214 267780 56102
rect 267832 22908 267884 22914
rect 267832 22850 267884 22856
rect 267740 4208 267792 4214
rect 267740 4150 267792 4156
rect 267844 3482 267872 22850
rect 268396 9450 268424 59191
rect 269776 10606 269804 59191
rect 269960 10674 269988 59463
rect 270236 59401 270264 59599
rect 272260 59401 272288 59758
rect 272522 59735 272578 59744
rect 275466 59800 275522 59809
rect 275466 59735 275522 59744
rect 276386 59800 276442 59809
rect 280618 59800 280674 59809
rect 276386 59735 276442 59744
rect 279424 59764 279476 59770
rect 272522 59664 272578 59673
rect 272522 59599 272578 59608
rect 275374 59664 275430 59673
rect 275374 59599 275430 59608
rect 270222 59392 270278 59401
rect 270222 59327 270278 59336
rect 271142 59392 271198 59401
rect 271142 59327 271198 59336
rect 272246 59392 272302 59401
rect 272246 59327 272302 59336
rect 270500 27056 270552 27062
rect 270500 26998 270552 27004
rect 270512 16574 270540 26998
rect 270512 16546 270816 16574
rect 270040 14748 270092 14754
rect 270040 14690 270092 14696
rect 269948 10668 270000 10674
rect 269948 10610 270000 10616
rect 269764 10600 269816 10606
rect 269764 10542 269816 10548
rect 268384 9444 268436 9450
rect 268384 9386 268436 9392
rect 268476 4208 268528 4214
rect 268476 4150 268528 4156
rect 267752 3454 267872 3482
rect 267752 480 267780 3454
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268488 354 268516 4150
rect 270052 480 270080 14690
rect 268814 354 268926 480
rect 268488 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 270788 354 270816 16546
rect 271156 9382 271184 59327
rect 271880 28552 271932 28558
rect 271880 28494 271932 28500
rect 271892 16574 271920 28494
rect 271892 16546 272472 16574
rect 271144 9376 271196 9382
rect 271144 9318 271196 9324
rect 272444 480 272472 16546
rect 272536 10538 272564 59599
rect 274086 59528 274142 59537
rect 274086 59463 274142 59472
rect 273902 59392 273958 59401
rect 273902 59327 273958 59336
rect 273260 12300 273312 12306
rect 273260 12242 273312 12248
rect 272524 10532 272576 10538
rect 272524 10474 272576 10480
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273272 354 273300 12242
rect 273916 10334 273944 59327
rect 274100 10402 274128 59463
rect 274640 54596 274692 54602
rect 274640 54538 274692 54544
rect 274652 16574 274680 54538
rect 275388 45554 275416 59599
rect 275480 59537 275508 59735
rect 275466 59528 275522 59537
rect 275466 59463 275522 59472
rect 276400 59401 276428 59735
rect 289818 59800 289874 59809
rect 280618 59735 280620 59744
rect 279424 59706 279476 59712
rect 280672 59735 280674 59744
rect 287704 59764 287756 59770
rect 280620 59706 280672 59712
rect 292946 59800 293002 59809
rect 289818 59735 289820 59744
rect 287704 59706 287756 59712
rect 289872 59735 289874 59744
rect 290648 59764 290700 59770
rect 289820 59706 289872 59712
rect 297086 59800 297142 59809
rect 292946 59735 292948 59744
rect 290648 59706 290700 59712
rect 293000 59735 293002 59744
rect 294604 59764 294656 59770
rect 292948 59706 293000 59712
rect 302238 59800 302294 59809
rect 297086 59735 297088 59744
rect 294604 59706 294656 59712
rect 297140 59735 297142 59744
rect 300124 59764 300176 59770
rect 297088 59706 297140 59712
rect 302238 59735 302240 59744
rect 300124 59706 300176 59712
rect 302292 59735 302294 59744
rect 306194 59800 306250 59809
rect 310518 59800 310574 59809
rect 306194 59735 306250 59744
rect 309048 59764 309100 59770
rect 302240 59706 302292 59712
rect 276386 59392 276442 59401
rect 276386 59327 276442 59336
rect 276662 59256 276718 59265
rect 276662 59191 276718 59200
rect 278226 59256 278282 59265
rect 278226 59191 278282 59200
rect 276020 47932 276072 47938
rect 276020 47874 276072 47880
rect 275296 45526 275416 45554
rect 274652 16546 274864 16574
rect 274088 10396 274140 10402
rect 274088 10338 274140 10344
rect 273904 10328 273956 10334
rect 273904 10270 273956 10276
rect 274836 480 274864 16546
rect 275296 9314 275324 45526
rect 275284 9308 275336 9314
rect 275284 9250 275336 9256
rect 276032 480 276060 47874
rect 276676 32570 276704 59191
rect 278042 59120 278098 59129
rect 278042 59055 278098 59064
rect 276664 32564 276716 32570
rect 276664 32506 276716 32512
rect 277400 32564 277452 32570
rect 277400 32506 277452 32512
rect 276664 12232 276716 12238
rect 276664 12174 276716 12180
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276676 354 276704 12174
rect 277412 6914 277440 32506
rect 278056 8974 278084 59055
rect 278240 17474 278268 59191
rect 279436 47734 279464 59706
rect 280802 59664 280858 59673
rect 286690 59664 286746 59673
rect 280802 59599 280858 59608
rect 284944 59628 284996 59634
rect 279424 47728 279476 47734
rect 279424 47670 279476 47676
rect 278780 24472 278832 24478
rect 278780 24414 278832 24420
rect 278228 17468 278280 17474
rect 278228 17410 278280 17416
rect 278792 16574 278820 24414
rect 278792 16546 279096 16574
rect 278044 8968 278096 8974
rect 278044 8910 278096 8916
rect 277412 6886 278360 6914
rect 278332 480 278360 6886
rect 277094 354 277206 480
rect 276676 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280816 14618 280844 59599
rect 286690 59599 286692 59608
rect 284944 59570 284996 59576
rect 286744 59599 286746 59608
rect 286692 59570 286744 59576
rect 282366 59528 282422 59537
rect 282184 59492 282236 59498
rect 282366 59463 282422 59472
rect 284666 59528 284722 59537
rect 284666 59463 284668 59472
rect 282184 59434 282236 59440
rect 280804 14612 280856 14618
rect 280804 14554 280856 14560
rect 280712 12164 280764 12170
rect 280712 12106 280764 12112
rect 280724 480 280752 12106
rect 282196 9042 282224 59434
rect 282380 23118 282408 59463
rect 284720 59463 284722 59472
rect 284668 59434 284720 59440
rect 283562 59392 283618 59401
rect 283562 59327 283618 59336
rect 283576 27266 283604 59327
rect 284956 32502 284984 59570
rect 286690 59528 286746 59537
rect 286690 59463 286746 59472
rect 286322 59256 286378 59265
rect 286322 59191 286378 59200
rect 284944 32496 284996 32502
rect 284944 32438 284996 32444
rect 283564 27260 283616 27266
rect 283564 27202 283616 27208
rect 282920 27192 282972 27198
rect 282920 27134 282972 27140
rect 282368 23112 282420 23118
rect 282368 23054 282420 23060
rect 282932 16574 282960 27134
rect 282932 16546 283144 16574
rect 282184 9036 282236 9042
rect 282184 8978 282236 8984
rect 281908 8968 281960 8974
rect 281908 8910 281960 8916
rect 281920 480 281948 8910
rect 283116 480 283144 16546
rect 284300 11824 284352 11830
rect 284300 11766 284352 11772
rect 284312 480 284340 11766
rect 286336 9178 286364 59191
rect 286704 45554 286732 59463
rect 286520 45526 286732 45554
rect 286520 9246 286548 45526
rect 287336 12096 287388 12102
rect 287336 12038 287388 12044
rect 286600 11824 286652 11830
rect 286600 11766 286652 11772
rect 286508 9240 286560 9246
rect 286508 9182 286560 9188
rect 286324 9172 286376 9178
rect 286324 9114 286376 9120
rect 285404 9036 285456 9042
rect 285404 8978 285456 8984
rect 285416 480 285444 8978
rect 286612 480 286640 11766
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 354 287376 12038
rect 287716 9110 287744 59706
rect 290462 59528 290518 59537
rect 290462 59463 290518 59472
rect 289082 59256 289138 59265
rect 289082 59191 289138 59200
rect 288440 53304 288492 53310
rect 288440 53246 288492 53252
rect 288452 16574 288480 53246
rect 289096 17338 289124 59191
rect 289820 32768 289872 32774
rect 289820 32710 289872 32716
rect 289084 17332 289136 17338
rect 289084 17274 289136 17280
rect 288452 16546 289032 16574
rect 287704 9104 287756 9110
rect 287704 9046 287756 9052
rect 289004 480 289032 16546
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 289832 354 289860 32710
rect 290476 14550 290504 59463
rect 290660 54670 290688 59706
rect 293222 59528 293278 59537
rect 293222 59463 293278 59472
rect 291842 59392 291898 59401
rect 291842 59327 291898 59336
rect 290648 54664 290700 54670
rect 290648 54606 290700 54612
rect 290464 14544 290516 14550
rect 290464 14486 290516 14492
rect 291384 12028 291436 12034
rect 291384 11970 291436 11976
rect 291396 480 291424 11970
rect 291856 3262 291884 59327
rect 292580 50652 292632 50658
rect 292580 50594 292632 50600
rect 292592 4214 292620 50594
rect 292672 36780 292724 36786
rect 292672 36722 292724 36728
rect 292580 4208 292632 4214
rect 292580 4150 292632 4156
rect 292684 3482 292712 36722
rect 293236 13122 293264 59463
rect 294616 31278 294644 59706
rect 299110 59664 299166 59673
rect 299110 59599 299166 59608
rect 296074 59528 296130 59537
rect 295812 59486 296074 59514
rect 295812 59401 295840 59486
rect 296074 59463 296130 59472
rect 298926 59528 298982 59537
rect 298926 59463 298982 59472
rect 294786 59392 294842 59401
rect 294786 59327 294842 59336
rect 295798 59392 295854 59401
rect 295798 59327 295854 59336
rect 295982 59392 296038 59401
rect 295982 59327 296038 59336
rect 294800 49162 294828 59327
rect 294788 49156 294840 49162
rect 294788 49098 294840 49104
rect 294604 31272 294656 31278
rect 294604 31214 294656 31220
rect 295996 22846 296024 59327
rect 297362 59256 297418 59265
rect 297362 59191 297418 59200
rect 298742 59256 298798 59265
rect 298742 59191 298798 59200
rect 296720 31340 296772 31346
rect 296720 31282 296772 31288
rect 295984 22840 296036 22846
rect 295984 22782 296036 22788
rect 296732 16574 296760 31282
rect 296732 16546 297312 16574
rect 293224 13116 293276 13122
rect 293224 13058 293276 13064
rect 294880 11960 294932 11966
rect 294880 11902 294932 11908
rect 293316 4208 293368 4214
rect 293316 4150 293368 4156
rect 292592 3454 292712 3482
rect 291844 3256 291896 3262
rect 291844 3198 291896 3204
rect 292592 480 292620 3454
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293328 354 293356 4150
rect 294892 480 294920 11902
rect 296076 9104 296128 9110
rect 296076 9046 296128 9052
rect 296088 480 296116 9046
rect 297284 480 297312 16546
rect 297376 11762 297404 59191
rect 298756 26994 298784 59191
rect 298940 45082 298968 59463
rect 299124 59401 299152 59599
rect 299110 59392 299166 59401
rect 299110 59327 299166 59336
rect 298928 45076 298980 45082
rect 298928 45018 298980 45024
rect 300136 40866 300164 59706
rect 303342 59528 303398 59537
rect 303342 59463 303398 59472
rect 301594 59256 301650 59265
rect 301594 59191 301650 59200
rect 301608 45554 301636 59191
rect 301516 45526 301636 45554
rect 300124 40860 300176 40866
rect 300124 40802 300176 40808
rect 298744 26988 298796 26994
rect 298744 26930 298796 26936
rect 300860 17536 300912 17542
rect 300860 17478 300912 17484
rect 298100 11892 298152 11898
rect 298100 11834 298152 11840
rect 297364 11756 297416 11762
rect 297364 11698 297416 11704
rect 293654 354 293766 480
rect 293328 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 354 298140 11834
rect 299480 11756 299532 11762
rect 299480 11698 299532 11704
rect 299492 3262 299520 11698
rect 299664 9172 299716 9178
rect 299664 9114 299716 9120
rect 299480 3256 299532 3262
rect 299480 3198 299532 3204
rect 299676 480 299704 9114
rect 300872 6914 300900 17478
rect 301516 14482 301544 45526
rect 303356 31278 303384 59463
rect 304906 59392 304962 59401
rect 304906 59327 304962 59336
rect 303620 54868 303672 54874
rect 303620 54810 303672 54816
rect 303344 31272 303396 31278
rect 303344 31214 303396 31220
rect 303632 16574 303660 54810
rect 304920 22846 304948 59327
rect 306208 58886 306236 59735
rect 310518 59735 310520 59744
rect 309048 59706 309100 59712
rect 310572 59735 310574 59744
rect 318430 59800 318486 59809
rect 318430 59735 318486 59744
rect 322202 59800 322258 59809
rect 322202 59735 322258 59744
rect 326710 59800 326766 59809
rect 338026 59800 338082 59809
rect 326710 59735 326712 59744
rect 310520 59706 310572 59712
rect 306286 59392 306342 59401
rect 306286 59327 306342 59336
rect 307574 59392 307630 59401
rect 307574 59327 307630 59336
rect 306196 58880 306248 58886
rect 306196 58822 306248 58828
rect 305000 36712 305052 36718
rect 305000 36654 305052 36660
rect 304908 22840 304960 22846
rect 304908 22782 304960 22788
rect 305012 16574 305040 36654
rect 306300 26994 306328 59327
rect 307390 59120 307446 59129
rect 307390 59055 307446 59064
rect 306288 26988 306340 26994
rect 306288 26930 306340 26936
rect 303632 16546 303936 16574
rect 305012 16546 305592 16574
rect 301504 14476 301556 14482
rect 301504 14418 301556 14424
rect 303160 9240 303212 9246
rect 303160 9182 303212 9188
rect 300872 6886 301544 6914
rect 300768 3256 300820 3262
rect 300768 3198 300820 3204
rect 300780 480 300808 3198
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 6886
rect 303172 480 303200 9182
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305564 480 305592 16546
rect 307404 14482 307432 59055
rect 307588 32502 307616 59327
rect 309060 54670 309088 59706
rect 310426 59528 310482 59537
rect 310426 59463 310482 59472
rect 311806 59528 311862 59537
rect 311806 59463 311862 59472
rect 318062 59528 318118 59537
rect 318062 59463 318118 59472
rect 309048 54664 309100 54670
rect 309048 54606 309100 54612
rect 310440 36718 310468 59463
rect 311622 59392 311678 59401
rect 311622 59327 311678 59336
rect 311636 53378 311664 59327
rect 311624 53372 311676 53378
rect 311624 53314 311676 53320
rect 310428 36712 310480 36718
rect 310428 36654 310480 36660
rect 307576 32496 307628 32502
rect 307576 32438 307628 32444
rect 307760 25900 307812 25906
rect 307760 25842 307812 25848
rect 307392 14476 307444 14482
rect 307392 14418 307444 14424
rect 306748 9308 306800 9314
rect 306748 9250 306800 9256
rect 306760 480 306788 9250
rect 307772 3482 307800 25842
rect 307852 14680 307904 14686
rect 307852 14622 307904 14628
rect 307864 4214 307892 14622
rect 311820 14550 311848 59463
rect 313280 51944 313332 51950
rect 313280 51886 313332 51892
rect 313292 16574 313320 51886
rect 316040 49156 316092 49162
rect 316040 49098 316092 49104
rect 313292 16546 313872 16574
rect 311808 14544 311860 14550
rect 311808 14486 311860 14492
rect 312176 13524 312228 13530
rect 312176 13466 312228 13472
rect 311440 13320 311492 13326
rect 311440 13262 311492 13268
rect 310244 9376 310296 9382
rect 310244 9318 310296 9324
rect 307852 4208 307904 4214
rect 307852 4150 307904 4156
rect 309048 4208 309100 4214
rect 309048 4150 309100 4156
rect 307772 3454 307984 3482
rect 307956 480 307984 3454
rect 309060 480 309088 4150
rect 310256 480 310284 9318
rect 311452 480 311480 13262
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 354 312216 13466
rect 313844 480 313872 16546
rect 314660 11892 314712 11898
rect 314660 11834 314712 11840
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314672 354 314700 11834
rect 316052 3262 316080 49098
rect 317420 34060 317472 34066
rect 317420 34002 317472 34008
rect 316224 13456 316276 13462
rect 316224 13398 316276 13404
rect 316040 3256 316092 3262
rect 316040 3198 316092 3204
rect 316236 480 316264 13398
rect 317432 6914 317460 34002
rect 318076 14618 318104 59463
rect 318444 59401 318472 59735
rect 320454 59664 320510 59673
rect 320454 59599 320510 59608
rect 322110 59664 322166 59673
rect 322216 59634 322244 59735
rect 326764 59735 326766 59744
rect 329288 59764 329340 59770
rect 326712 59706 326764 59712
rect 342166 59800 342222 59809
rect 338026 59735 338028 59744
rect 329288 59706 329340 59712
rect 338080 59735 338082 59744
rect 339500 59764 339552 59770
rect 338028 59706 338080 59712
rect 351182 59800 351238 59809
rect 342166 59735 342168 59744
rect 339500 59706 339552 59712
rect 342220 59735 342222 59744
rect 344284 59764 344336 59770
rect 342168 59706 342220 59712
rect 354678 59800 354734 59809
rect 351238 59758 351500 59786
rect 351182 59735 351238 59744
rect 344284 59706 344336 59712
rect 328734 59664 328790 59673
rect 322110 59599 322166 59608
rect 322204 59628 322256 59634
rect 318430 59392 318486 59401
rect 318430 59327 318486 59336
rect 319442 59256 319498 59265
rect 319442 59191 319498 59200
rect 319456 14686 319484 59191
rect 320468 58410 320496 59599
rect 321006 59528 321062 59537
rect 321006 59463 321062 59472
rect 320822 59392 320878 59401
rect 320822 59327 320878 59336
rect 320456 58404 320508 58410
rect 320456 58346 320508 58352
rect 320836 14754 320864 59327
rect 321020 50590 321048 59463
rect 322124 58546 322152 59599
rect 322204 59570 322256 59576
rect 325148 59628 325200 59634
rect 328734 59599 328736 59608
rect 325148 59570 325200 59576
rect 328788 59599 328790 59608
rect 328736 59570 328788 59576
rect 324962 59392 325018 59401
rect 324962 59327 325018 59336
rect 322112 58540 322164 58546
rect 322112 58482 322164 58488
rect 323584 58540 323636 58546
rect 323584 58482 323636 58488
rect 322204 58404 322256 58410
rect 322204 58346 322256 58352
rect 321008 50584 321060 50590
rect 321008 50526 321060 50532
rect 322216 38078 322244 58346
rect 323596 47734 323624 58482
rect 323584 47728 323636 47734
rect 323584 47670 323636 47676
rect 324976 43586 325004 59327
rect 325160 49230 325188 59570
rect 325698 59528 325754 59537
rect 325698 59463 325754 59472
rect 328734 59528 328790 59537
rect 328734 59463 328790 59472
rect 325148 49224 325200 49230
rect 325148 49166 325200 49172
rect 325712 46442 325740 59463
rect 327722 59392 327778 59401
rect 327722 59327 327778 59336
rect 325700 46436 325752 46442
rect 325700 46378 325752 46384
rect 325700 45144 325752 45150
rect 325700 45086 325752 45092
rect 324964 43580 325016 43586
rect 324964 43522 325016 43528
rect 324320 38140 324372 38146
rect 324320 38082 324372 38088
rect 322204 38072 322256 38078
rect 322204 38014 322256 38020
rect 320824 14748 320876 14754
rect 320824 14690 320876 14696
rect 319444 14680 319496 14686
rect 319444 14622 319496 14628
rect 318064 14612 318116 14618
rect 318064 14554 318116 14560
rect 319720 13388 319772 13394
rect 319720 13330 319772 13336
rect 322112 13388 322164 13394
rect 322112 13330 322164 13336
rect 317432 6886 318104 6914
rect 317328 3256 317380 3262
rect 317328 3198 317380 3204
rect 317340 480 317368 3198
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 6886
rect 319732 480 319760 13330
rect 320456 13116 320508 13122
rect 320456 13058 320508 13064
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 13058
rect 322124 480 322152 13330
rect 322940 13252 322992 13258
rect 322940 13194 322992 13200
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 322952 354 322980 13194
rect 324332 3074 324360 38082
rect 325712 16574 325740 45086
rect 327736 39574 327764 59327
rect 328460 59016 328512 59022
rect 328460 58958 328512 58964
rect 327724 39568 327776 39574
rect 327724 39510 327776 39516
rect 327080 39500 327132 39506
rect 327080 39442 327132 39448
rect 327092 16574 327120 39442
rect 328472 16574 328500 58958
rect 328748 51074 328776 59463
rect 328748 51046 329144 51074
rect 329116 28490 329144 51046
rect 329300 40866 329328 59706
rect 333886 59664 333942 59673
rect 330484 59628 330536 59634
rect 333886 59599 333942 59608
rect 330484 59570 330536 59576
rect 329288 40860 329340 40866
rect 329288 40802 329340 40808
rect 330496 29850 330524 59570
rect 330850 59528 330906 59537
rect 331862 59528 331918 59537
rect 330906 59486 331076 59514
rect 330850 59463 330906 59472
rect 331048 59265 331076 59486
rect 331918 59486 332640 59514
rect 331862 59463 331918 59472
rect 331862 59392 331918 59401
rect 331862 59327 331918 59336
rect 331034 59256 331090 59265
rect 331034 59191 331090 59200
rect 331220 43648 331272 43654
rect 331220 43590 331272 43596
rect 330484 29844 330536 29850
rect 330484 29786 330536 29792
rect 329104 28484 329156 28490
rect 329104 28426 329156 28432
rect 325712 16546 326384 16574
rect 327092 16546 328040 16574
rect 328472 16546 328776 16574
rect 324412 11960 324464 11966
rect 324412 11902 324464 11908
rect 324424 3262 324452 11902
rect 324412 3256 324464 3262
rect 324412 3198 324464 3204
rect 325608 3256 325660 3262
rect 325608 3198 325660 3204
rect 324332 3046 324452 3074
rect 324424 480 324452 3046
rect 325620 480 325648 3198
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 16546
rect 328012 480 328040 16546
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 328748 354 328776 16546
rect 330392 13184 330444 13190
rect 330392 13126 330444 13132
rect 330404 480 330432 13126
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331232 354 331260 43590
rect 331876 42294 331904 59327
rect 332612 52018 332640 59486
rect 333900 59401 333928 59599
rect 334622 59528 334678 59537
rect 334622 59463 334678 59472
rect 337566 59528 337622 59537
rect 337566 59463 337622 59472
rect 333242 59392 333298 59401
rect 333242 59327 333298 59336
rect 333886 59392 333942 59401
rect 333886 59327 333942 59336
rect 332600 52012 332652 52018
rect 332600 51954 332652 51960
rect 331864 42288 331916 42294
rect 331864 42230 331916 42236
rect 332600 35556 332652 35562
rect 332600 35498 332652 35504
rect 332612 3074 332640 35498
rect 333256 24342 333284 59327
rect 334636 45150 334664 59463
rect 337382 59392 337438 59401
rect 337382 59327 337438 59336
rect 335358 59256 335414 59265
rect 335358 59191 335414 59200
rect 335372 56098 335400 59191
rect 335360 56092 335412 56098
rect 335360 56034 335412 56040
rect 334624 45144 334676 45150
rect 334624 45086 334676 45092
rect 337396 41002 337424 59327
rect 337580 45218 337608 59463
rect 338762 59256 338818 59265
rect 338762 59191 338818 59200
rect 338120 46572 338172 46578
rect 338120 46514 338172 46520
rect 337568 45212 337620 45218
rect 337568 45154 337620 45160
rect 336740 40996 336792 41002
rect 336740 40938 336792 40944
rect 337384 40996 337436 41002
rect 337384 40938 337436 40944
rect 333980 40928 334032 40934
rect 333980 40870 334032 40876
rect 333244 24336 333296 24342
rect 333244 24278 333296 24284
rect 332692 17400 332744 17406
rect 332692 17342 332744 17348
rect 332704 3262 332732 17342
rect 333992 16574 334020 40870
rect 336752 16574 336780 40938
rect 338132 16574 338160 46514
rect 338776 43790 338804 59191
rect 339512 57458 339540 59706
rect 341522 59528 341578 59537
rect 341522 59463 341578 59472
rect 340880 57520 340932 57526
rect 340880 57462 340932 57468
rect 339500 57452 339552 57458
rect 339500 57394 339552 57400
rect 338764 43784 338816 43790
rect 338764 43726 338816 43732
rect 333992 16546 334664 16574
rect 336752 16546 337056 16574
rect 338132 16546 338712 16574
rect 332692 3256 332744 3262
rect 332692 3198 332744 3204
rect 333888 3256 333940 3262
rect 333888 3198 333940 3204
rect 332612 3046 332732 3074
rect 332704 480 332732 3046
rect 333900 480 333928 3198
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 336280 13252 336332 13258
rect 336280 13194 336332 13200
rect 336292 480 336320 13194
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 338684 480 338712 16546
rect 339500 12028 339552 12034
rect 339500 11970 339552 11976
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339512 354 339540 11970
rect 340892 3074 340920 57462
rect 341536 13190 341564 59463
rect 341706 59392 341762 59401
rect 341706 59327 341762 59336
rect 341720 47870 341748 59327
rect 342902 59256 342958 59265
rect 342902 59191 342958 59200
rect 342260 57588 342312 57594
rect 342260 57530 342312 57536
rect 341708 47864 341760 47870
rect 341708 47806 341760 47812
rect 342272 16574 342300 57530
rect 342916 17338 342944 59191
rect 344296 17406 344324 59706
rect 345294 59664 345350 59673
rect 351182 59664 351238 59673
rect 345294 59599 345296 59608
rect 345348 59599 345350 59608
rect 347044 59628 347096 59634
rect 345296 59570 345348 59576
rect 351182 59599 351238 59608
rect 347044 59570 347096 59576
rect 345294 59528 345350 59537
rect 345294 59463 345350 59472
rect 345308 55214 345336 59463
rect 345846 59256 345902 59265
rect 345846 59191 345902 59200
rect 345308 55186 345704 55214
rect 345020 42356 345072 42362
rect 345020 42298 345072 42304
rect 344284 17400 344336 17406
rect 344284 17342 344336 17348
rect 342904 17332 342956 17338
rect 342904 17274 342956 17280
rect 345032 16574 345060 42298
rect 345676 17542 345704 55186
rect 345664 17536 345716 17542
rect 345664 17478 345716 17484
rect 345860 17474 345888 59191
rect 347056 17610 347084 59570
rect 347410 59528 347466 59537
rect 347410 59463 347466 59472
rect 349802 59528 349858 59537
rect 349802 59463 349858 59472
rect 347424 59265 347452 59463
rect 348422 59392 348478 59401
rect 348422 59327 348478 59336
rect 347410 59256 347466 59265
rect 347410 59191 347466 59200
rect 348436 17678 348464 59327
rect 349160 45076 349212 45082
rect 349160 45018 349212 45024
rect 348424 17672 348476 17678
rect 348424 17614 348476 17620
rect 347044 17604 347096 17610
rect 347044 17546 347096 17552
rect 345848 17468 345900 17474
rect 345848 17410 345900 17416
rect 342272 16546 342944 16574
rect 345032 16546 345336 16574
rect 341524 13184 341576 13190
rect 341524 13126 341576 13132
rect 340972 10328 341024 10334
rect 340972 10270 341024 10276
rect 340984 3262 341012 10270
rect 340972 3256 341024 3262
rect 340972 3198 341024 3204
rect 342168 3256 342220 3262
rect 342168 3198 342220 3204
rect 340892 3046 341012 3074
rect 340984 480 341012 3046
rect 342180 480 342208 3198
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 16546
rect 344560 16244 344612 16250
rect 344560 16186 344612 16192
rect 344572 480 344600 16186
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 16546
rect 348056 16176 348108 16182
rect 348056 16118 348108 16124
rect 346952 12096 347004 12102
rect 346952 12038 347004 12044
rect 346964 480 346992 12038
rect 348068 480 348096 16118
rect 349172 3074 349200 45018
rect 349252 21752 349304 21758
rect 349252 21694 349304 21700
rect 349264 3262 349292 21694
rect 349816 17814 349844 59463
rect 349986 59392 350042 59401
rect 349986 59327 350042 59336
rect 349804 17808 349856 17814
rect 349804 17750 349856 17756
rect 350000 17746 350028 59327
rect 351196 17882 351224 59599
rect 351472 59401 351500 59758
rect 359462 59800 359518 59809
rect 354678 59735 354680 59744
rect 354732 59735 354734 59744
rect 356704 59764 356756 59770
rect 354680 59706 354732 59712
rect 360934 59800 360990 59809
rect 359518 59758 359780 59786
rect 359462 59735 359518 59744
rect 356704 59706 356756 59712
rect 353942 59528 353998 59537
rect 353942 59463 353998 59472
rect 351458 59392 351514 59401
rect 351458 59327 351514 59336
rect 352562 59392 352618 59401
rect 352562 59327 352618 59336
rect 352576 35494 352604 59327
rect 353298 59256 353354 59265
rect 353298 59191 353354 59200
rect 353312 56234 353340 59191
rect 353300 56228 353352 56234
rect 353300 56170 353352 56176
rect 352564 35488 352616 35494
rect 352564 35430 352616 35436
rect 353956 27266 353984 59463
rect 355322 59256 355378 59265
rect 355322 59191 355378 59200
rect 355336 50726 355364 59191
rect 355324 50720 355376 50726
rect 355324 50662 355376 50668
rect 356716 32706 356744 59706
rect 359462 59664 359518 59673
rect 359462 59599 359518 59608
rect 358266 59528 358322 59537
rect 358266 59463 358322 59472
rect 358082 59392 358138 59401
rect 358082 59327 358138 59336
rect 356704 32700 356756 32706
rect 356704 32642 356756 32648
rect 353944 27260 353996 27266
rect 353944 27202 353996 27208
rect 357440 23112 357492 23118
rect 357440 23054 357492 23060
rect 351184 17876 351236 17882
rect 351184 17818 351236 17824
rect 349988 17740 350040 17746
rect 349988 17682 350040 17688
rect 351184 16108 351236 16114
rect 351184 16050 351236 16056
rect 349252 3256 349304 3262
rect 349252 3198 349304 3204
rect 350448 3256 350500 3262
rect 350448 3198 350500 3204
rect 349172 3046 349292 3074
rect 349264 480 349292 3046
rect 350460 480 350488 3198
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16050
rect 353576 13524 353628 13530
rect 353576 13466 353628 13472
rect 352840 10396 352892 10402
rect 352840 10338 352892 10344
rect 352852 480 352880 10338
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 353588 354 353616 13466
rect 355232 10464 355284 10470
rect 355232 10406 355284 10412
rect 356336 10464 356388 10470
rect 356336 10406 356388 10412
rect 355244 480 355272 10406
rect 356348 480 356376 10406
rect 357452 3074 357480 23054
rect 358096 16046 358124 59327
rect 358280 34134 358308 59463
rect 358268 34128 358320 34134
rect 358268 34070 358320 34076
rect 357532 16040 357584 16046
rect 357532 15982 357584 15988
rect 358084 16040 358136 16046
rect 358084 15982 358136 15988
rect 357544 3262 357572 15982
rect 359476 13462 359504 59599
rect 359752 59537 359780 59758
rect 360934 59735 360990 59744
rect 364246 59800 364302 59809
rect 364246 59735 364302 59744
rect 371146 59800 371202 59809
rect 371146 59735 371202 59744
rect 372158 59800 372160 59809
rect 373724 59832 373776 59838
rect 372212 59800 372214 59809
rect 372158 59735 372214 59744
rect 373722 59800 373724 59809
rect 430120 59832 430172 59838
rect 373776 59800 373778 59809
rect 373722 59735 373778 59744
rect 374182 59800 374238 59809
rect 374182 59735 374238 59744
rect 376482 59800 376538 59809
rect 376482 59735 376538 59744
rect 376758 59800 376814 59809
rect 376758 59735 376814 59744
rect 384118 59800 384174 59809
rect 384118 59735 384174 59744
rect 384486 59800 384542 59809
rect 384486 59735 384542 59744
rect 388718 59800 388774 59809
rect 389086 59800 389142 59809
rect 388774 59758 389086 59786
rect 388718 59735 388774 59744
rect 389086 59735 389142 59744
rect 392858 59800 392914 59809
rect 400126 59800 400182 59809
rect 392858 59735 392860 59744
rect 359738 59528 359794 59537
rect 359738 59463 359794 59472
rect 360842 59528 360898 59537
rect 360842 59463 360898 59472
rect 360856 16114 360884 59463
rect 360948 59401 360976 59735
rect 362866 59664 362922 59673
rect 362866 59599 362922 59608
rect 362880 59401 362908 59599
rect 364260 59537 364288 59735
rect 365902 59664 365958 59673
rect 365902 59599 365958 59608
rect 363602 59528 363658 59537
rect 363602 59463 363658 59472
rect 364246 59528 364302 59537
rect 364246 59463 364302 59472
rect 365810 59528 365866 59537
rect 365810 59463 365866 59472
rect 360934 59392 360990 59401
rect 360934 59327 360990 59336
rect 362222 59392 362278 59401
rect 362222 59327 362278 59336
rect 362866 59392 362922 59401
rect 362866 59327 362922 59336
rect 362130 59256 362186 59265
rect 362130 59191 362186 59200
rect 362144 54806 362172 59191
rect 362236 59090 362264 59327
rect 362224 59084 362276 59090
rect 362224 59026 362276 59032
rect 361580 54800 361632 54806
rect 361580 54742 361632 54748
rect 362132 54800 362184 54806
rect 362132 54742 362184 54748
rect 361592 16574 361620 54742
rect 361592 16546 361896 16574
rect 360844 16108 360896 16114
rect 360844 16050 360896 16056
rect 359464 13456 359516 13462
rect 359464 13398 359516 13404
rect 361120 10872 361172 10878
rect 361120 10814 361172 10820
rect 359464 10532 359516 10538
rect 359464 10474 359516 10480
rect 357532 3256 357584 3262
rect 357532 3198 357584 3204
rect 358728 3256 358780 3262
rect 358728 3198 358780 3204
rect 357452 3046 357572 3074
rect 357544 480 357572 3046
rect 358740 480 358768 3198
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 10474
rect 361132 480 361160 10814
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 361868 354 361896 16546
rect 363616 16182 363644 59463
rect 365824 59430 365852 59463
rect 365812 59424 365864 59430
rect 364982 59392 365038 59401
rect 365812 59366 365864 59372
rect 364982 59327 365038 59336
rect 364340 47116 364392 47122
rect 364340 47058 364392 47064
rect 364352 16574 364380 47058
rect 364996 35630 365024 59327
rect 365916 55214 365944 59599
rect 367098 59528 367154 59537
rect 367098 59463 367154 59472
rect 370134 59528 370190 59537
rect 370134 59463 370190 59472
rect 366548 59424 366600 59430
rect 366548 59366 366600 59372
rect 365916 55186 366404 55214
rect 364984 35624 365036 35630
rect 364984 35566 365036 35572
rect 364352 16546 364656 16574
rect 363604 16176 363656 16182
rect 363604 16118 363656 16124
rect 363512 10600 363564 10606
rect 363512 10542 363564 10548
rect 363524 480 363552 10542
rect 364628 480 364656 16546
rect 366376 15978 366404 55186
rect 366560 16250 366588 59366
rect 366548 16244 366600 16250
rect 366548 16186 366600 16192
rect 365720 15972 365772 15978
rect 365720 15914 365772 15920
rect 366364 15972 366416 15978
rect 366364 15914 366416 15920
rect 365732 3074 365760 15914
rect 365812 10668 365864 10674
rect 365812 10610 365864 10616
rect 365824 3262 365852 10610
rect 367112 6914 367140 59463
rect 367742 59392 367798 59401
rect 367742 59327 367798 59336
rect 369950 59392 370006 59401
rect 369950 59327 370006 59336
rect 367756 15366 367784 59327
rect 369964 47122 369992 59327
rect 369952 47116 370004 47122
rect 369952 47058 370004 47064
rect 368480 35420 368532 35426
rect 368480 35362 368532 35368
rect 368492 16574 368520 35362
rect 368492 16546 369440 16574
rect 367744 15360 367796 15366
rect 367744 15302 367796 15308
rect 367112 6886 367784 6914
rect 365812 3256 365864 3262
rect 365812 3198 365864 3204
rect 367008 3256 367060 3262
rect 367008 3198 367060 3204
rect 365732 3046 365852 3074
rect 365824 480 365852 3046
rect 367020 480 367048 3198
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 6886
rect 369412 480 369440 16546
rect 370148 10878 370176 59463
rect 371160 59401 371188 59735
rect 371238 59664 371294 59673
rect 371238 59599 371294 59608
rect 371146 59392 371202 59401
rect 371146 59327 371202 59336
rect 371252 23118 371280 59599
rect 373998 59392 374054 59401
rect 373998 59327 374054 59336
rect 372710 59256 372766 59265
rect 372710 59191 372766 59200
rect 372620 36848 372672 36854
rect 372620 36790 372672 36796
rect 371240 23112 371292 23118
rect 371240 23054 371292 23060
rect 371240 15360 371292 15366
rect 371240 15302 371292 15308
rect 370136 10872 370188 10878
rect 370136 10814 370188 10820
rect 370136 10736 370188 10742
rect 370136 10678 370188 10684
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370148 354 370176 10678
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 371252 354 371280 15302
rect 372632 6914 372660 36790
rect 372724 13530 372752 59191
rect 374012 57594 374040 59327
rect 374000 57588 374052 57594
rect 374000 57530 374052 57536
rect 374092 57520 374144 57526
rect 374092 57462 374144 57468
rect 374104 56386 374132 57462
rect 374012 56358 374132 56386
rect 372712 13524 372764 13530
rect 372712 13466 372764 13472
rect 372632 6886 372936 6914
rect 372908 480 372936 6886
rect 374012 3074 374040 56358
rect 374196 45554 374224 59735
rect 376496 59537 376524 59735
rect 376482 59528 376538 59537
rect 376482 59463 376538 59472
rect 374274 59392 374330 59401
rect 374274 59327 374330 59336
rect 374104 45526 374224 45554
rect 374104 21758 374132 45526
rect 374092 21752 374144 21758
rect 374092 21694 374144 21700
rect 374092 16244 374144 16250
rect 374092 16186 374144 16192
rect 374104 3262 374132 16186
rect 374288 12102 374316 59327
rect 376772 59022 376800 59735
rect 378414 59664 378470 59673
rect 378414 59599 378470 59608
rect 383750 59664 383806 59673
rect 383750 59599 383806 59608
rect 378230 59528 378286 59537
rect 378230 59463 378286 59472
rect 376850 59392 376906 59401
rect 376850 59327 376906 59336
rect 376760 59016 376812 59022
rect 376760 58958 376812 58964
rect 376760 24404 376812 24410
rect 376760 24346 376812 24352
rect 375380 20460 375432 20466
rect 375380 20402 375432 20408
rect 375392 16574 375420 20402
rect 375392 16546 376064 16574
rect 374276 12096 374328 12102
rect 374276 12038 374328 12044
rect 374092 3256 374144 3262
rect 374092 3198 374144 3204
rect 375288 3256 375340 3262
rect 375288 3198 375340 3204
rect 374012 3046 374132 3074
rect 374104 480 374132 3046
rect 375300 480 375328 3198
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 376772 6914 376800 24346
rect 376864 12034 376892 59327
rect 378244 35562 378272 59463
rect 378232 35556 378284 35562
rect 378232 35498 378284 35504
rect 378324 15972 378376 15978
rect 378324 15914 378376 15920
rect 376852 12028 376904 12034
rect 376852 11970 376904 11976
rect 378336 6914 378364 15914
rect 378428 13258 378456 59599
rect 382278 59528 382334 59537
rect 382278 59463 382334 59472
rect 380990 59256 381046 59265
rect 380990 59191 381046 59200
rect 379520 56024 379572 56030
rect 379520 55966 379572 55972
rect 378416 13252 378468 13258
rect 378416 13194 378468 13200
rect 376772 6886 377720 6914
rect 378336 6886 378456 6914
rect 377692 480 377720 6886
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 6886
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 379532 354 379560 55966
rect 381004 11966 381032 59191
rect 382292 34066 382320 59463
rect 382462 59392 382518 59401
rect 382462 59327 382518 59336
rect 382280 34060 382332 34066
rect 382280 34002 382332 34008
rect 382372 20392 382424 20398
rect 382372 20334 382424 20340
rect 382384 16574 382412 20334
rect 382292 16546 382412 16574
rect 381176 15972 381228 15978
rect 381176 15914 381228 15920
rect 380992 11960 381044 11966
rect 380992 11902 381044 11908
rect 381188 480 381216 15914
rect 382292 3262 382320 16546
rect 382476 13394 382504 59327
rect 382556 35624 382608 35630
rect 382556 35566 382608 35572
rect 382464 13388 382516 13394
rect 382464 13330 382516 13336
rect 382568 6914 382596 35566
rect 383660 25832 383712 25838
rect 383660 25774 383712 25780
rect 382384 6886 382596 6914
rect 383672 6914 383700 25774
rect 383764 11898 383792 59599
rect 384132 58410 384160 59735
rect 384500 59430 384528 59735
rect 392912 59735 392914 59744
rect 394884 59764 394936 59770
rect 392860 59706 392912 59712
rect 404174 59800 404230 59809
rect 400126 59735 400128 59744
rect 394884 59706 394936 59712
rect 400180 59735 400182 59744
rect 401600 59764 401652 59770
rect 400128 59706 400180 59712
rect 404174 59735 404230 59744
rect 409510 59800 409566 59809
rect 412638 59800 412694 59809
rect 409510 59735 409512 59744
rect 401600 59706 401652 59712
rect 390650 59664 390706 59673
rect 390650 59599 390706 59608
rect 387890 59528 387946 59537
rect 387890 59463 387946 59472
rect 384488 59424 384540 59430
rect 385224 59424 385276 59430
rect 384488 59366 384540 59372
rect 385222 59392 385224 59401
rect 385276 59392 385278 59401
rect 385222 59327 385278 59336
rect 386602 59392 386658 59401
rect 386602 59327 386658 59336
rect 386418 59256 386474 59265
rect 386418 59191 386474 59200
rect 384120 58404 384172 58410
rect 384120 58346 384172 58352
rect 385040 58404 385092 58410
rect 385040 58346 385092 58352
rect 385052 13326 385080 58346
rect 386432 54874 386460 59191
rect 386420 54868 386472 54874
rect 386420 54810 386472 54816
rect 386420 42424 386472 42430
rect 386420 42366 386472 42372
rect 386432 16574 386460 42366
rect 386616 25906 386644 59327
rect 387800 28620 387852 28626
rect 387800 28562 387852 28568
rect 386604 25900 386656 25906
rect 386604 25842 386656 25848
rect 386432 16546 386736 16574
rect 385960 16176 386012 16182
rect 385960 16118 386012 16124
rect 385040 13320 385092 13326
rect 385040 13262 385092 13268
rect 383752 11892 383804 11898
rect 383752 11834 383804 11840
rect 383672 6886 384344 6914
rect 382280 3256 382332 3262
rect 382280 3198 382332 3204
rect 382384 480 382412 6886
rect 383568 3256 383620 3262
rect 383568 3198 383620 3204
rect 383580 480 383608 3198
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 378846 -960 378958 326
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 6886
rect 385972 480 386000 16118
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 386708 354 386736 16546
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 28562
rect 387904 11762 387932 59463
rect 389270 59256 389326 59265
rect 389270 59191 389326 59200
rect 389180 59084 389232 59090
rect 389180 59026 389232 59032
rect 389192 16574 389220 59026
rect 389284 31346 389312 59191
rect 390664 50658 390692 59599
rect 392030 59528 392086 59537
rect 392030 59463 392086 59472
rect 394698 59528 394754 59537
rect 394698 59463 394754 59472
rect 390834 59392 390890 59401
rect 390834 59327 390890 59336
rect 390652 50652 390704 50658
rect 390652 50594 390704 50600
rect 390848 32774 390876 59327
rect 391940 54800 391992 54806
rect 391940 54742 391992 54748
rect 390836 32768 390888 32774
rect 390836 32710 390888 32716
rect 390560 32632 390612 32638
rect 390560 32574 390612 32580
rect 389272 31340 389324 31346
rect 389272 31282 389324 31288
rect 389192 16546 389496 16574
rect 387892 11756 387944 11762
rect 387892 11698 387944 11704
rect 389468 480 389496 16546
rect 390572 3074 390600 32574
rect 390652 11756 390704 11762
rect 390652 11698 390704 11704
rect 390664 3262 390692 11698
rect 391952 6914 391980 54742
rect 392044 11830 392072 59463
rect 393410 59392 393466 59401
rect 393410 59327 393466 59336
rect 393320 39636 393372 39642
rect 393320 39578 393372 39584
rect 393332 16574 393360 39578
rect 393424 27198 393452 59327
rect 394712 56166 394740 59463
rect 394790 59256 394846 59265
rect 394790 59191 394846 59200
rect 394700 56160 394752 56166
rect 394700 56102 394752 56108
rect 394804 47938 394832 59191
rect 394792 47932 394844 47938
rect 394792 47874 394844 47880
rect 394700 29980 394752 29986
rect 394700 29922 394752 29928
rect 393412 27192 393464 27198
rect 393412 27134 393464 27140
rect 394712 16574 394740 29922
rect 394896 24478 394924 59706
rect 399114 59528 399170 59537
rect 399114 59463 399170 59472
rect 400218 59528 400274 59537
rect 400218 59463 400274 59472
rect 398930 59392 398986 59401
rect 398930 59327 398986 59336
rect 396078 59256 396134 59265
rect 396078 59191 396134 59200
rect 396092 28558 396120 59191
rect 398840 31340 398892 31346
rect 398840 31282 398892 31288
rect 396080 28552 396132 28558
rect 396080 28494 396132 28500
rect 394884 24472 394936 24478
rect 394884 24414 394936 24420
rect 397460 22976 397512 22982
rect 397460 22918 397512 22924
rect 397472 16574 397500 22918
rect 393332 16546 394280 16574
rect 394712 16546 395384 16574
rect 397472 16546 397776 16574
rect 392032 11824 392084 11830
rect 392032 11766 392084 11772
rect 391952 6886 392624 6914
rect 390652 3256 390704 3262
rect 390652 3198 390704 3204
rect 391848 3256 391900 3262
rect 391848 3198 391900 3204
rect 390572 3046 390692 3074
rect 390664 480 390692 3046
rect 391860 480 391888 3198
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 6886
rect 394252 480 394280 16546
rect 395356 480 395384 16546
rect 396080 16108 396132 16114
rect 396080 16050 396132 16056
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 16050
rect 397748 480 397776 16546
rect 398852 3074 398880 31282
rect 398944 23050 398972 59327
rect 399128 29918 399156 59463
rect 400232 49298 400260 59463
rect 400220 49292 400272 49298
rect 400220 49234 400272 49240
rect 400220 46504 400272 46510
rect 400220 46446 400272 46452
rect 399116 29912 399168 29918
rect 399116 29854 399168 29860
rect 398932 23044 398984 23050
rect 398932 22986 398984 22992
rect 400232 16574 400260 46446
rect 401612 38282 401640 59706
rect 403162 59528 403218 59537
rect 403162 59463 403218 59472
rect 402978 59392 403034 59401
rect 402978 59327 403034 59336
rect 402992 39710 403020 59327
rect 402980 39704 403032 39710
rect 402980 39646 403032 39652
rect 401600 38276 401652 38282
rect 401600 38218 401652 38224
rect 402980 34128 403032 34134
rect 402980 34070 403032 34076
rect 402992 16574 403020 34070
rect 400232 16546 400904 16574
rect 402992 16546 403112 16574
rect 398932 13456 398984 13462
rect 398932 13398 398984 13404
rect 398944 3262 398972 13398
rect 398932 3256 398984 3262
rect 398932 3198 398984 3204
rect 400128 3256 400180 3262
rect 400128 3198 400180 3204
rect 398852 3046 398972 3074
rect 398944 480 398972 3046
rect 400140 480 400168 3198
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 16546
rect 402520 13252 402572 13258
rect 402520 13194 402572 13200
rect 402532 480 402560 13194
rect 403084 3482 403112 16546
rect 403176 6594 403204 59463
rect 404188 59401 404216 59735
rect 409564 59735 409566 59744
rect 411628 59764 411680 59770
rect 409512 59706 409564 59712
rect 418710 59800 418766 59809
rect 412638 59735 412640 59744
rect 411628 59706 411680 59712
rect 412692 59735 412694 59744
rect 414112 59764 414164 59770
rect 412640 59706 412692 59712
rect 423678 59800 423734 59809
rect 418710 59735 418712 59744
rect 414112 59706 414164 59712
rect 418764 59735 418766 59744
rect 419816 59764 419868 59770
rect 418712 59706 418764 59712
rect 423678 59735 423734 59744
rect 430118 59800 430120 59809
rect 431500 59832 431552 59838
rect 430172 59800 430174 59809
rect 430118 59735 430174 59744
rect 431498 59800 431500 59809
rect 488080 59832 488132 59838
rect 431552 59800 431554 59809
rect 431498 59735 431554 59744
rect 431958 59800 432014 59809
rect 431958 59735 432014 59744
rect 433154 59800 433210 59809
rect 433154 59735 433210 59744
rect 437478 59800 437534 59809
rect 437754 59800 437810 59809
rect 437534 59758 437754 59786
rect 437478 59735 437534 59744
rect 437754 59735 437810 59744
rect 438858 59800 438914 59809
rect 438858 59735 438914 59744
rect 444470 59800 444526 59809
rect 444470 59735 444526 59744
rect 446678 59800 446734 59809
rect 454958 59800 455014 59809
rect 446678 59735 446680 59744
rect 419816 59706 419868 59712
rect 404266 59664 404322 59673
rect 408590 59664 408646 59673
rect 404322 59622 404400 59650
rect 404266 59599 404322 59608
rect 404174 59392 404230 59401
rect 404174 59327 404230 59336
rect 404372 55214 404400 59622
rect 408590 59599 408646 59608
rect 405278 59528 405334 59537
rect 405278 59463 405280 59472
rect 405332 59463 405334 59472
rect 407118 59528 407174 59537
rect 407118 59463 407174 59472
rect 407304 59492 407356 59498
rect 405280 59434 405332 59440
rect 405830 59392 405886 59401
rect 405830 59327 405886 59336
rect 404372 55186 404492 55214
rect 404360 21684 404412 21690
rect 404360 21626 404412 21632
rect 403164 6588 403216 6594
rect 403164 6530 403216 6536
rect 403084 3454 403664 3482
rect 403636 480 403664 3454
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 21626
rect 404464 6526 404492 55186
rect 405740 11824 405792 11830
rect 405740 11766 405792 11772
rect 404452 6520 404504 6526
rect 404452 6462 404504 6468
rect 405752 3482 405780 11766
rect 405844 6458 405872 59327
rect 407132 43722 407160 59463
rect 407304 59434 407356 59440
rect 407120 43716 407172 43722
rect 407120 43658 407172 43664
rect 407120 38208 407172 38214
rect 407120 38150 407172 38156
rect 405832 6452 405884 6458
rect 405832 6394 405884 6400
rect 405752 3454 406056 3482
rect 406028 480 406056 3454
rect 407132 3262 407160 38150
rect 407316 25770 407344 59434
rect 407304 25764 407356 25770
rect 407304 25706 407356 25712
rect 408500 21684 408552 21690
rect 408500 21626 408552 21632
rect 407212 16040 407264 16046
rect 407212 15982 407264 15988
rect 407120 3256 407172 3262
rect 407120 3198 407172 3204
rect 407224 480 407252 15982
rect 408408 3256 408460 3262
rect 408408 3198 408460 3204
rect 408420 480 408448 3198
rect 408512 626 408540 21626
rect 408604 6390 408632 59599
rect 409970 59256 410026 59265
rect 409970 59191 410026 59200
rect 411442 59256 411498 59265
rect 411442 59191 411498 59200
rect 409880 32700 409932 32706
rect 409880 32642 409932 32648
rect 408592 6384 408644 6390
rect 408592 6326 408644 6332
rect 409892 3482 409920 32642
rect 409984 6322 410012 59191
rect 411260 47796 411312 47802
rect 411260 47738 411312 47744
rect 411272 16574 411300 47738
rect 411272 16546 411392 16574
rect 409972 6316 410024 6322
rect 409972 6258 410024 6264
rect 411364 3482 411392 16546
rect 411456 6186 411484 59191
rect 411640 6254 411668 59706
rect 413190 59528 413246 59537
rect 413190 59463 413246 59472
rect 412638 59256 412694 59265
rect 412638 59191 412694 59200
rect 412652 40798 412680 59191
rect 413204 57390 413232 59463
rect 413192 57384 413244 57390
rect 413192 57326 413244 57332
rect 414020 50720 414072 50726
rect 414020 50662 414072 50668
rect 412640 40792 412692 40798
rect 412640 40734 412692 40740
rect 412640 11892 412692 11898
rect 412640 11834 412692 11840
rect 411628 6248 411680 6254
rect 411628 6190 411680 6196
rect 411444 6180 411496 6186
rect 411444 6122 411496 6128
rect 409892 3454 410840 3482
rect 411364 3454 411944 3482
rect 408512 598 409184 626
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 598
rect 410812 480 410840 3454
rect 411916 480 411944 3454
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 11834
rect 414032 3482 414060 50662
rect 414124 5098 414152 59706
rect 416870 59528 416926 59537
rect 416870 59463 416926 59472
rect 419630 59528 419686 59537
rect 419630 59463 419686 59472
rect 415582 59392 415638 59401
rect 415582 59327 415638 59336
rect 415596 46374 415624 59327
rect 415584 46368 415636 46374
rect 415584 46310 415636 46316
rect 416780 27260 416832 27266
rect 416780 27202 416832 27208
rect 415400 27124 415452 27130
rect 415400 27066 415452 27072
rect 415412 16574 415440 27066
rect 415412 16546 415532 16574
rect 414112 5092 414164 5098
rect 414112 5034 414164 5040
rect 414032 3454 414336 3482
rect 414308 480 414336 3454
rect 415504 480 415532 16546
rect 416688 6384 416740 6390
rect 416688 6326 416740 6332
rect 416700 480 416728 6326
rect 416792 626 416820 27202
rect 416884 5030 416912 59463
rect 418250 59392 418306 59401
rect 418250 59327 418306 59336
rect 418160 54732 418212 54738
rect 418160 54674 418212 54680
rect 416872 5024 416924 5030
rect 416872 4966 416924 4972
rect 416792 598 417464 626
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 598
rect 418172 490 418200 54674
rect 418264 4962 418292 59327
rect 419644 45014 419672 59463
rect 419632 45008 419684 45014
rect 419632 44950 419684 44956
rect 419828 33998 419856 59706
rect 420826 59528 420882 59537
rect 420826 59463 420828 59472
rect 420880 59463 420882 59472
rect 422392 59492 422444 59498
rect 420828 59434 420880 59440
rect 422392 59434 422444 59440
rect 421010 59256 421066 59265
rect 421010 59191 421066 59200
rect 420920 56228 420972 56234
rect 420920 56170 420972 56176
rect 419816 33992 419868 33998
rect 419816 33934 419868 33940
rect 420184 16040 420236 16046
rect 420184 15982 420236 15988
rect 418252 4956 418304 4962
rect 418252 4898 418304 4904
rect 417854 354 417966 480
rect 418172 462 418568 490
rect 420196 480 420224 15982
rect 417436 326 417966 354
rect 418540 354 418568 462
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 56170
rect 421024 4894 421052 59191
rect 422300 21616 422352 21622
rect 422300 21558 422352 21564
rect 421012 4888 421064 4894
rect 421012 4830 421064 4836
rect 422312 3482 422340 21558
rect 422404 4826 422432 59434
rect 423692 55962 423720 59735
rect 424966 59664 425022 59673
rect 425022 59622 425192 59650
rect 424966 59599 425022 59608
rect 423862 59528 423918 59537
rect 423862 59463 423918 59472
rect 423770 59392 423826 59401
rect 423770 59327 423826 59336
rect 423680 55956 423732 55962
rect 423680 55898 423732 55904
rect 423784 45554 423812 59327
rect 423692 45526 423812 45554
rect 423692 35358 423720 45526
rect 423772 35420 423824 35426
rect 423772 35362 423824 35368
rect 423680 35352 423732 35358
rect 423680 35294 423732 35300
rect 422392 4820 422444 4826
rect 422392 4762 422444 4768
rect 422312 3454 422616 3482
rect 422588 480 422616 3454
rect 423784 480 423812 35362
rect 423876 24274 423904 59463
rect 425060 58948 425112 58954
rect 425060 58890 425112 58896
rect 423956 35488 424008 35494
rect 423956 35430 424008 35436
rect 423864 24268 423916 24274
rect 423864 24210 423916 24216
rect 423968 16574 423996 35430
rect 425072 16574 425100 58890
rect 425164 28422 425192 59622
rect 425334 59528 425390 59537
rect 425334 59463 425390 59472
rect 429198 59528 429254 59537
rect 429198 59463 429254 59472
rect 425348 57322 425376 59463
rect 428002 59392 428058 59401
rect 428002 59327 428058 59336
rect 425336 57316 425388 57322
rect 425336 57258 425388 57264
rect 428016 29782 428044 59327
rect 429212 38010 429240 59463
rect 430670 59392 430726 59401
rect 430670 59327 430726 59336
rect 430580 56228 430632 56234
rect 430580 56170 430632 56176
rect 429200 38004 429252 38010
rect 429200 37946 429252 37952
rect 428004 29776 428056 29782
rect 428004 29718 428056 29724
rect 425152 28416 425204 28422
rect 425152 28358 425204 28364
rect 426440 22976 426492 22982
rect 426440 22918 426492 22924
rect 426452 16574 426480 22918
rect 429200 21548 429252 21554
rect 429200 21490 429252 21496
rect 427820 17876 427872 17882
rect 427820 17818 427872 17824
rect 427832 16574 427860 17818
rect 423968 16546 425008 16574
rect 425072 16546 425744 16574
rect 426452 16546 426848 16574
rect 427832 16546 428504 16574
rect 424980 480 425008 16546
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 16546
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 16546
rect 428476 480 428504 16546
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429212 354 429240 21490
rect 430592 16574 430620 56170
rect 430684 17270 430712 59327
rect 431972 39438 432000 59735
rect 432142 59528 432198 59537
rect 432142 59463 432198 59472
rect 431960 39432 432012 39438
rect 431960 39374 432012 39380
rect 431960 21480 432012 21486
rect 431960 21422 432012 21428
rect 430672 17264 430724 17270
rect 430672 17206 430724 17212
rect 430592 16546 430896 16574
rect 430868 480 430896 16546
rect 431972 3262 432000 21422
rect 432052 17808 432104 17814
rect 432052 17750 432104 17756
rect 431960 3256 432012 3262
rect 431960 3198 432012 3204
rect 432064 480 432092 17750
rect 432156 15910 432184 59463
rect 433168 59401 433196 59735
rect 433246 59664 433302 59673
rect 437386 59664 437442 59673
rect 433302 59622 433380 59650
rect 433246 59599 433302 59608
rect 433154 59392 433210 59401
rect 433154 59327 433210 59336
rect 433352 49094 433380 59622
rect 437442 59622 437520 59650
rect 437386 59599 437442 59608
rect 434258 59528 434314 59537
rect 434258 59463 434314 59472
rect 436190 59528 436246 59537
rect 436190 59463 436246 59472
rect 434272 59265 434300 59463
rect 434718 59392 434774 59401
rect 434718 59327 434774 59336
rect 434258 59256 434314 59265
rect 434258 59191 434314 59200
rect 434732 53242 434760 59327
rect 434720 53236 434772 53242
rect 434720 53178 434772 53184
rect 436204 51882 436232 59463
rect 436374 59392 436430 59401
rect 436374 59327 436430 59336
rect 436192 51876 436244 51882
rect 436192 51818 436244 51824
rect 433340 49088 433392 49094
rect 433340 49030 433392 49036
rect 436388 36650 436416 59327
rect 437492 42158 437520 59622
rect 437480 42152 437532 42158
rect 437480 42094 437532 42100
rect 436376 36644 436428 36650
rect 436376 36586 436428 36592
rect 437480 32632 437532 32638
rect 437480 32574 437532 32580
rect 433340 27124 433392 27130
rect 433340 27066 433392 27072
rect 433352 16574 433380 27066
rect 436100 21412 436152 21418
rect 436100 21354 436152 21360
rect 434720 17740 434772 17746
rect 434720 17682 434772 17688
rect 434732 16574 434760 17682
rect 436112 16574 436140 21354
rect 433352 16546 434024 16574
rect 434732 16546 435128 16574
rect 436112 16546 436784 16574
rect 432144 15904 432196 15910
rect 432144 15846 432196 15852
rect 433248 3256 433300 3262
rect 433248 3198 433300 3204
rect 433260 480 433288 3198
rect 429630 354 429742 480
rect 429212 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 16546
rect 436756 480 436784 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 32574
rect 438872 31142 438900 59735
rect 441066 59664 441122 59673
rect 441066 59599 441122 59608
rect 441080 59401 441108 59599
rect 444484 59537 444512 59735
rect 446732 59735 446734 59744
rect 449348 59764 449400 59770
rect 446680 59706 446732 59712
rect 457994 59800 458050 59809
rect 454958 59735 454960 59744
rect 449348 59706 449400 59712
rect 455012 59735 455014 59744
rect 457628 59764 457680 59770
rect 454960 59706 455012 59712
rect 458362 59800 458418 59809
rect 458050 59758 458362 59786
rect 457994 59735 458050 59744
rect 458362 59735 458418 59744
rect 459926 59800 459982 59809
rect 459926 59735 459982 59744
rect 467286 59800 467342 59809
rect 476026 59800 476082 59809
rect 467286 59735 467288 59744
rect 457628 59706 457680 59712
rect 444562 59664 444618 59673
rect 444562 59599 444618 59608
rect 448702 59664 448758 59673
rect 448702 59599 448758 59608
rect 443550 59528 443606 59537
rect 444470 59528 444526 59537
rect 443550 59463 443552 59472
rect 443604 59463 443606 59472
rect 444380 59492 444432 59498
rect 443552 59434 443604 59440
rect 444470 59463 444526 59472
rect 444380 59434 444432 59440
rect 441066 59392 441122 59401
rect 441066 59327 441122 59336
rect 442262 59392 442318 59401
rect 442262 59327 442318 59336
rect 443642 59392 443698 59401
rect 443642 59327 443698 59336
rect 441066 59256 441122 59265
rect 441066 59191 441122 59200
rect 440882 59120 440938 59129
rect 440882 59055 440938 59064
rect 440240 44940 440292 44946
rect 440240 44882 440292 44888
rect 438860 31136 438912 31142
rect 438860 31078 438912 31084
rect 438860 17672 438912 17678
rect 438860 17614 438912 17620
rect 438872 16574 438900 17614
rect 438872 16546 439176 16574
rect 439148 480 439176 16546
rect 440252 3074 440280 44882
rect 440332 17672 440384 17678
rect 440332 17614 440384 17620
rect 440344 3262 440372 17614
rect 440896 6186 440924 59055
rect 441080 6254 441108 59191
rect 441620 17604 441672 17610
rect 441620 17546 441672 17552
rect 441632 16574 441660 17546
rect 441632 16546 442212 16574
rect 441068 6248 441120 6254
rect 441068 6190 441120 6196
rect 440884 6180 440936 6186
rect 440884 6122 440936 6128
rect 442184 3482 442212 16546
rect 442276 6322 442304 59327
rect 443656 21418 443684 59327
rect 444392 55962 444420 59434
rect 444576 57322 444604 59599
rect 446402 59528 446458 59537
rect 446402 59463 446458 59472
rect 444564 57316 444616 57322
rect 444564 57258 444616 57264
rect 444380 55956 444432 55962
rect 444380 55898 444432 55904
rect 444380 36644 444432 36650
rect 444380 36586 444432 36592
rect 443644 21412 443696 21418
rect 443644 21354 443696 21360
rect 444392 16574 444420 36586
rect 446416 35358 446444 59463
rect 448716 59401 448744 59599
rect 449162 59528 449218 59537
rect 449162 59463 449218 59472
rect 447782 59392 447838 59401
rect 447782 59327 447838 59336
rect 448702 59392 448758 59401
rect 448702 59327 448758 59336
rect 446404 35352 446456 35358
rect 446404 35294 446456 35300
rect 447796 33998 447824 59327
rect 448520 38004 448572 38010
rect 448520 37946 448572 37952
rect 447784 33992 447836 33998
rect 447784 33934 447836 33940
rect 445760 17536 445812 17542
rect 445760 17478 445812 17484
rect 444392 16546 445064 16574
rect 442264 6316 442316 6322
rect 442264 6258 442316 6264
rect 442184 3454 442672 3482
rect 440332 3256 440384 3262
rect 440332 3198 440384 3204
rect 441528 3256 441580 3262
rect 441528 3198 441580 3204
rect 440252 3046 440372 3074
rect 440344 480 440372 3046
rect 441540 480 441568 3198
rect 442644 480 442672 3454
rect 443828 3324 443880 3330
rect 443828 3266 443880 3272
rect 443840 480 443868 3266
rect 445036 480 445064 16546
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 354 445800 17478
rect 447416 3392 447468 3398
rect 447416 3334 447468 3340
rect 447428 480 447456 3334
rect 448532 3210 448560 37946
rect 449176 29782 449204 59463
rect 449360 31142 449388 59706
rect 449714 59664 449770 59673
rect 449714 59599 449770 59608
rect 449728 58954 449756 59599
rect 454682 59528 454738 59537
rect 454682 59463 454738 59472
rect 457442 59528 457498 59537
rect 457442 59463 457498 59472
rect 453302 59392 453358 59401
rect 453302 59327 453358 59336
rect 450542 59256 450598 59265
rect 450542 59191 450598 59200
rect 449716 58948 449768 58954
rect 449716 58890 449768 58896
rect 449348 31136 449400 31142
rect 449348 31078 449400 31084
rect 449164 29776 449216 29782
rect 449164 29718 449216 29724
rect 450556 28422 450584 59191
rect 450544 28416 450596 28422
rect 450544 28358 450596 28364
rect 448612 17468 448664 17474
rect 448612 17410 448664 17416
rect 451280 17468 451332 17474
rect 451280 17410 451332 17416
rect 448624 3398 448652 17410
rect 451292 16574 451320 17410
rect 452660 17400 452712 17406
rect 452660 17342 452712 17348
rect 451292 16546 451688 16574
rect 450912 4140 450964 4146
rect 450912 4082 450964 4088
rect 448612 3392 448664 3398
rect 448612 3334 448664 3340
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 448532 3182 448652 3210
rect 448624 480 448652 3182
rect 449820 480 449848 3334
rect 450924 480 450952 4082
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 452672 6914 452700 17342
rect 453316 16574 453344 59327
rect 453486 59120 453542 59129
rect 453486 59055 453542 59064
rect 453316 16546 453436 16574
rect 452672 6886 453344 6914
rect 453316 480 453344 6886
rect 453408 4894 453436 16546
rect 453396 4888 453448 4894
rect 453396 4830 453448 4836
rect 453500 4826 453528 59055
rect 454696 4962 454724 59463
rect 456062 59392 456118 59401
rect 456062 59327 456118 59336
rect 456076 17270 456104 59327
rect 456892 17332 456944 17338
rect 456892 17274 456944 17280
rect 456064 17264 456116 17270
rect 456064 17206 456116 17212
rect 455696 11960 455748 11966
rect 455696 11902 455748 11908
rect 454684 4956 454736 4962
rect 454684 4898 454736 4904
rect 453488 4820 453540 4826
rect 453488 4762 453540 4768
rect 454500 4072 454552 4078
rect 454500 4014 454552 4020
rect 454512 480 454540 4014
rect 455708 480 455736 11902
rect 456904 480 456932 17274
rect 457456 5098 457484 59463
rect 457444 5092 457496 5098
rect 457444 5034 457496 5040
rect 457640 5030 457668 59706
rect 458822 59256 458878 59265
rect 458822 59191 458878 59200
rect 458180 54732 458232 54738
rect 458180 54674 458232 54680
rect 458192 16574 458220 54674
rect 458192 16546 458772 16574
rect 457628 5024 457680 5030
rect 457628 4966 457680 4972
rect 458088 4004 458140 4010
rect 458088 3946 458140 3952
rect 458100 480 458128 3946
rect 458744 3482 458772 16546
rect 458836 5166 458864 59191
rect 459940 55214 459968 59735
rect 467340 59735 467342 59744
rect 468484 59764 468536 59770
rect 467288 59706 467340 59712
rect 476026 59735 476082 59744
rect 484858 59800 484914 59809
rect 484858 59735 484914 59744
rect 485778 59800 485834 59809
rect 485778 59735 485834 59744
rect 488078 59800 488080 59809
rect 489368 59832 489420 59838
rect 488132 59800 488134 59809
rect 488078 59735 488134 59744
rect 489366 59800 489368 59809
rect 498476 59832 498528 59838
rect 489420 59800 489422 59809
rect 489366 59735 489422 59744
rect 490102 59800 490158 59809
rect 490102 59735 490158 59744
rect 491022 59800 491078 59809
rect 491022 59735 491078 59744
rect 495622 59800 495678 59809
rect 495622 59735 495678 59744
rect 498474 59800 498476 59809
rect 499488 59832 499540 59838
rect 498528 59800 498530 59809
rect 516968 59832 517020 59838
rect 508686 59800 508742 59809
rect 499540 59780 499712 59786
rect 499488 59774 499712 59780
rect 499500 59758 499712 59774
rect 498474 59735 498530 59744
rect 468484 59706 468536 59712
rect 461122 59664 461178 59673
rect 467102 59664 467158 59673
rect 461122 59599 461124 59608
rect 461176 59599 461178 59608
rect 462964 59628 463016 59634
rect 461124 59570 461176 59576
rect 467102 59599 467158 59608
rect 462964 59570 463016 59576
rect 461122 59528 461178 59537
rect 461178 59486 461256 59514
rect 461122 59463 461178 59472
rect 461122 59392 461178 59401
rect 461122 59327 461178 59336
rect 461136 55214 461164 59327
rect 461228 58970 461256 59486
rect 461228 58942 461716 58970
rect 461688 55214 461716 58942
rect 459940 55186 460244 55214
rect 461136 55186 461624 55214
rect 461688 55186 461808 55214
rect 459928 13184 459980 13190
rect 459928 13126 459980 13132
rect 458824 5160 458876 5166
rect 458824 5102 458876 5108
rect 458744 3454 459232 3482
rect 459204 480 459232 3454
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 13126
rect 460216 5234 460244 55186
rect 461596 15910 461624 55186
rect 461780 25770 461808 55186
rect 461768 25764 461820 25770
rect 461768 25706 461820 25712
rect 462320 21548 462372 21554
rect 462320 21490 462372 21496
rect 461584 15904 461636 15910
rect 461584 15846 461636 15852
rect 460204 5228 460256 5234
rect 460204 5170 460256 5176
rect 461584 3936 461636 3942
rect 461584 3878 461636 3884
rect 461596 480 461624 3878
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 21490
rect 462976 13190 463004 59570
rect 463238 59528 463294 59537
rect 463238 59463 463294 59472
rect 465722 59528 465778 59537
rect 465722 59463 465778 59472
rect 463252 59265 463280 59463
rect 464342 59392 464398 59401
rect 464342 59327 464398 59336
rect 463238 59256 463294 59265
rect 463238 59191 463294 59200
rect 463700 47864 463752 47870
rect 463700 47806 463752 47812
rect 463712 16574 463740 47806
rect 464356 24274 464384 59327
rect 464344 24268 464396 24274
rect 464344 24210 464396 24216
rect 465736 17338 465764 59463
rect 465906 59392 465962 59401
rect 465906 59327 465962 59336
rect 465920 21486 465948 59327
rect 466460 57452 466512 57458
rect 466460 57394 466512 57400
rect 465908 21480 465960 21486
rect 465908 21422 465960 21428
rect 465724 17332 465776 17338
rect 465724 17274 465776 17280
rect 463712 16546 464016 16574
rect 462964 13184 463016 13190
rect 462964 13126 463016 13132
rect 463988 480 464016 16546
rect 465816 12980 465868 12986
rect 465816 12922 465868 12928
rect 465172 3868 465224 3874
rect 465172 3810 465224 3816
rect 465184 480 465212 3810
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 354 465856 12922
rect 466472 6914 466500 57394
rect 467116 16114 467144 59599
rect 467104 16108 467156 16114
rect 467104 16050 467156 16056
rect 468496 13326 468524 59706
rect 471978 59664 472034 59673
rect 471978 59599 472034 59608
rect 473358 59664 473414 59673
rect 473358 59599 473414 59608
rect 474554 59664 474610 59673
rect 474554 59599 474610 59608
rect 470690 59528 470746 59537
rect 470690 59463 470746 59472
rect 469862 59392 469918 59401
rect 469862 59327 469918 59336
rect 469218 59256 469274 59265
rect 469218 59191 469274 59200
rect 469232 53242 469260 59191
rect 469220 53236 469272 53242
rect 469220 53178 469272 53184
rect 469876 46374 469904 59327
rect 469864 46368 469916 46374
rect 469864 46310 469916 46316
rect 470600 43784 470652 43790
rect 470600 43726 470652 43732
rect 469864 13796 469916 13802
rect 469864 13738 469916 13744
rect 468484 13320 468536 13326
rect 468484 13262 468536 13268
rect 466472 6886 467512 6914
rect 467484 480 467512 6886
rect 468668 3800 468720 3806
rect 468668 3742 468720 3748
rect 468680 480 468708 3742
rect 469876 480 469904 13738
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 354 470640 43726
rect 470704 13802 470732 59463
rect 470692 13796 470744 13802
rect 470692 13738 470744 13744
rect 471992 12986 472020 59599
rect 473372 54738 473400 59599
rect 474568 59401 474596 59599
rect 476040 59537 476068 59735
rect 477590 59664 477646 59673
rect 480258 59664 480314 59673
rect 477646 59622 477724 59650
rect 477590 59599 477646 59608
rect 474738 59528 474794 59537
rect 474738 59463 474794 59472
rect 476026 59528 476082 59537
rect 476026 59463 476082 59472
rect 473542 59392 473598 59401
rect 473542 59327 473598 59336
rect 474554 59392 474610 59401
rect 474554 59327 474610 59336
rect 473360 54732 473412 54738
rect 473360 54674 473412 54680
rect 473360 46368 473412 46374
rect 473360 46310 473412 46316
rect 471980 12980 472032 12986
rect 471980 12922 472032 12928
rect 473372 6914 473400 46310
rect 473452 45212 473504 45218
rect 473452 45154 473504 45160
rect 473464 16574 473492 45154
rect 473556 21554 473584 59327
rect 473544 21548 473596 21554
rect 473544 21490 473596 21496
rect 473464 16546 474136 16574
rect 473372 6886 473492 6914
rect 472256 3732 472308 3738
rect 472256 3674 472308 3680
rect 472268 480 472296 3674
rect 473464 480 473492 6886
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 16546
rect 474752 11966 474780 59463
rect 476210 59392 476266 59401
rect 476210 59327 476266 59336
rect 477590 59392 477646 59401
rect 477590 59327 477646 59336
rect 476120 53236 476172 53242
rect 476120 53178 476172 53184
rect 476132 16574 476160 53178
rect 476224 17474 476252 59327
rect 477500 40996 477552 41002
rect 477500 40938 477552 40944
rect 476212 17468 476264 17474
rect 476212 17410 476264 17416
rect 477512 16574 477540 40938
rect 477604 36650 477632 59327
rect 477696 51074 477724 59622
rect 480258 59599 480314 59608
rect 481638 59664 481694 59673
rect 481638 59599 481694 59608
rect 482834 59664 482890 59673
rect 482834 59599 482890 59608
rect 478878 59528 478934 59537
rect 478878 59463 478934 59472
rect 477696 51046 477816 51074
rect 477788 38010 477816 51046
rect 477776 38004 477828 38010
rect 477776 37946 477828 37952
rect 477592 36644 477644 36650
rect 477592 36586 477644 36592
rect 478892 17678 478920 59463
rect 480272 32638 480300 59599
rect 481652 56234 481680 59599
rect 482848 59401 482876 59599
rect 484872 59537 484900 59735
rect 483018 59528 483074 59537
rect 483018 59463 483074 59472
rect 484858 59528 484914 59537
rect 484858 59463 484914 59472
rect 481822 59392 481878 59401
rect 481822 59327 481878 59336
rect 482834 59392 482890 59401
rect 482834 59327 482890 59336
rect 481640 56228 481692 56234
rect 481640 56170 481692 56176
rect 481640 56092 481692 56098
rect 481640 56034 481692 56040
rect 480260 32632 480312 32638
rect 480260 32574 480312 32580
rect 478880 17672 478932 17678
rect 478880 17614 478932 17620
rect 476132 16546 476528 16574
rect 477512 16546 478184 16574
rect 474740 11960 474792 11966
rect 474740 11902 474792 11908
rect 475752 3664 475804 3670
rect 475752 3606 475804 3612
rect 475764 480 475792 3606
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 478156 480 478184 16546
rect 480536 13320 480588 13326
rect 480536 13262 480588 13268
rect 479340 3528 479392 3534
rect 479340 3470 479392 3476
rect 479352 480 479380 3470
rect 480548 480 480576 13262
rect 481652 6914 481680 56034
rect 481732 46300 481784 46306
rect 481732 46242 481784 46248
rect 481744 16574 481772 46242
rect 481836 27130 481864 59327
rect 481824 27124 481876 27130
rect 481824 27066 481876 27072
rect 483032 22982 483060 59463
rect 485792 59401 485820 59735
rect 485962 59664 486018 59673
rect 485962 59599 486018 59608
rect 484490 59392 484546 59401
rect 484490 59327 484546 59336
rect 485778 59392 485834 59401
rect 485778 59327 485834 59336
rect 484400 45144 484452 45150
rect 484400 45086 484452 45092
rect 483020 22976 483072 22982
rect 483020 22918 483072 22924
rect 484412 16574 484440 45086
rect 484504 35426 484532 59327
rect 485780 42220 485832 42226
rect 485780 42162 485832 42168
rect 484492 35420 484544 35426
rect 484492 35362 484544 35368
rect 481744 16546 482416 16574
rect 484412 16546 484808 16574
rect 481652 6886 481772 6914
rect 481744 480 481772 6886
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 354 482416 16546
rect 484032 16108 484084 16114
rect 484032 16050 484084 16056
rect 484044 480 484072 16050
rect 482806 354 482918 480
rect 482388 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 485792 6914 485820 42162
rect 485976 16046 486004 59599
rect 486146 59528 486202 59537
rect 486146 59463 486202 59472
rect 489918 59528 489974 59537
rect 489918 59463 489974 59472
rect 485964 16040 486016 16046
rect 485964 15982 486016 15988
rect 485792 6886 486096 6914
rect 486068 3482 486096 6886
rect 486160 6390 486188 59463
rect 487250 59392 487306 59401
rect 487250 59327 487306 59336
rect 488630 59392 488686 59401
rect 488630 59327 488686 59336
rect 487160 17332 487212 17338
rect 487160 17274 487212 17280
rect 486148 6384 486200 6390
rect 486148 6326 486200 6332
rect 486068 3454 486464 3482
rect 486436 480 486464 3454
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487172 354 487200 17274
rect 487264 11898 487292 59327
rect 488540 52012 488592 52018
rect 488540 51954 488592 51960
rect 488552 16574 488580 51954
rect 488644 21690 488672 59327
rect 488632 21684 488684 21690
rect 488632 21626 488684 21632
rect 488552 16546 488856 16574
rect 487252 11892 487304 11898
rect 487252 11834 487304 11840
rect 488828 480 488856 16546
rect 489932 13258 489960 59463
rect 490012 19168 490064 19174
rect 490012 19110 490064 19116
rect 489920 13252 489972 13258
rect 489920 13194 489972 13200
rect 490024 6914 490052 19110
rect 490116 11830 490144 59735
rect 491036 59401 491064 59735
rect 491114 59664 491170 59673
rect 491170 59622 491340 59650
rect 491114 59599 491170 59608
rect 491022 59392 491078 59401
rect 491022 59327 491078 59336
rect 491312 31346 491340 59622
rect 492126 59528 492182 59537
rect 492126 59463 492128 59472
rect 492180 59463 492182 59472
rect 494058 59528 494114 59537
rect 494058 59463 494114 59472
rect 494244 59492 494296 59498
rect 492128 59434 492180 59440
rect 492678 59392 492734 59401
rect 492678 59327 492734 59336
rect 491300 31340 491352 31346
rect 491300 31282 491352 31288
rect 492692 29986 492720 59327
rect 492680 29980 492732 29986
rect 492680 29922 492732 29928
rect 494072 28626 494100 59463
rect 494244 59434 494296 59440
rect 494060 28620 494112 28626
rect 494060 28562 494112 28568
rect 491300 24336 491352 24342
rect 491300 24278 491352 24284
rect 490196 21480 490248 21486
rect 490196 21422 490248 21428
rect 490208 16574 490236 21422
rect 491312 16574 491340 24278
rect 494060 24268 494112 24274
rect 494060 24210 494112 24216
rect 492680 19100 492732 19106
rect 492680 19042 492732 19048
rect 492692 16574 492720 19042
rect 490208 16546 490696 16574
rect 491312 16546 492352 16574
rect 492692 16546 493088 16574
rect 490104 11824 490156 11830
rect 490104 11766 490156 11772
rect 489932 6886 490052 6914
rect 489932 480 489960 6886
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490668 354 490696 16546
rect 492324 480 492352 16546
rect 491086 354 491198 480
rect 490668 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494072 6914 494100 24210
rect 494256 11762 494284 59434
rect 495530 59392 495586 59401
rect 495530 59327 495586 59336
rect 495440 42288 495492 42294
rect 495440 42230 495492 42236
rect 494244 11756 494296 11762
rect 494244 11698 494296 11704
rect 494072 6886 494744 6914
rect 494716 480 494744 6886
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 42230
rect 495544 25838 495572 59327
rect 495636 57526 495664 59735
rect 498382 59664 498438 59673
rect 498382 59599 498438 59608
rect 496818 59528 496874 59537
rect 496818 59463 496874 59472
rect 495624 57520 495676 57526
rect 495624 57462 495676 57468
rect 495532 25832 495584 25838
rect 495532 25774 495584 25780
rect 496832 15978 496860 59463
rect 498200 29844 498252 29850
rect 498200 29786 498252 29792
rect 496912 19032 496964 19038
rect 496912 18974 496964 18980
rect 496924 16574 496952 18974
rect 496924 16546 497136 16574
rect 496820 15972 496872 15978
rect 496820 15914 496872 15920
rect 497108 480 497136 16546
rect 498212 3534 498240 29786
rect 498396 24410 498424 59599
rect 498384 24404 498436 24410
rect 498384 24346 498436 24352
rect 499580 18964 499632 18970
rect 499580 18906 499632 18912
rect 498292 13184 498344 13190
rect 498292 13126 498344 13132
rect 498200 3528 498252 3534
rect 498200 3470 498252 3476
rect 498304 3346 498332 13126
rect 499592 6914 499620 18906
rect 499684 10742 499712 59758
rect 509054 59800 509110 59809
rect 508742 59758 509054 59786
rect 508686 59735 508742 59744
rect 509054 59735 509110 59744
rect 512826 59800 512882 59809
rect 515954 59800 516010 59809
rect 512826 59735 512828 59744
rect 512880 59735 512882 59744
rect 514852 59764 514904 59770
rect 512828 59706 512880 59712
rect 515954 59735 516010 59744
rect 516966 59800 516968 59809
rect 518348 59832 518400 59838
rect 517020 59800 517022 59809
rect 516966 59735 517022 59744
rect 518346 59800 518348 59809
rect 518400 59800 518402 59809
rect 518346 59735 518402 59744
rect 518990 59800 519046 59809
rect 518990 59735 519046 59744
rect 520094 59800 520150 59809
rect 520094 59735 520150 59744
rect 522026 59800 522082 59809
rect 522026 59735 522082 59744
rect 524234 59800 524290 59809
rect 524234 59735 524290 59744
rect 525246 59800 525302 59809
rect 528650 59800 528706 59809
rect 525246 59735 525248 59744
rect 514852 59706 514904 59712
rect 507858 59664 507914 59673
rect 507858 59599 507914 59608
rect 510710 59664 510766 59673
rect 510766 59622 510844 59650
rect 510710 59599 510766 59608
rect 502706 59528 502762 59537
rect 502706 59463 502762 59472
rect 504546 59528 504602 59537
rect 504546 59463 504548 59472
rect 502522 59392 502578 59401
rect 502522 59327 502578 59336
rect 501050 59256 501106 59265
rect 501050 59191 501106 59200
rect 500960 25764 501012 25770
rect 500960 25706 501012 25712
rect 499672 10736 499724 10742
rect 499672 10678 499724 10684
rect 500972 6914 501000 25706
rect 501064 10674 501092 59191
rect 502340 28484 502392 28490
rect 502340 28426 502392 28432
rect 501052 10668 501104 10674
rect 501052 10610 501104 10616
rect 502352 6914 502380 28426
rect 502536 10606 502564 59327
rect 502524 10600 502576 10606
rect 502524 10542 502576 10548
rect 502720 10538 502748 59463
rect 504600 59463 504602 59472
rect 506478 59528 506534 59537
rect 506478 59463 506534 59472
rect 506664 59492 506716 59498
rect 504548 59434 504600 59440
rect 505190 59392 505246 59401
rect 505190 59327 505246 59336
rect 503810 59256 503866 59265
rect 503810 59191 503866 59200
rect 503720 18896 503772 18902
rect 503720 18838 503772 18844
rect 502708 10532 502760 10538
rect 502708 10474 502760 10480
rect 499592 6886 500632 6914
rect 500972 6886 501368 6914
rect 502352 6886 503024 6914
rect 499028 3528 499080 3534
rect 499028 3470 499080 3476
rect 498212 3318 498332 3346
rect 498212 480 498240 3318
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499040 354 499068 3470
rect 500604 480 500632 6886
rect 499366 354 499478 480
rect 499040 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501340 354 501368 6886
rect 502996 480 503024 6886
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503732 354 503760 18838
rect 503824 10470 503852 59191
rect 503812 10464 503864 10470
rect 503812 10406 503864 10412
rect 505204 10402 505232 59327
rect 506492 42362 506520 59463
rect 506664 59434 506716 59440
rect 506676 45082 506704 59434
rect 506664 45076 506716 45082
rect 506664 45018 506716 45024
rect 506480 42356 506532 42362
rect 506480 42298 506532 42304
rect 506480 40860 506532 40866
rect 506480 40802 506532 40808
rect 505376 15904 505428 15910
rect 505376 15846 505428 15852
rect 505192 10396 505244 10402
rect 505192 10338 505244 10344
rect 505388 480 505416 15846
rect 506492 480 506520 40802
rect 506572 18828 506624 18834
rect 506572 18770 506624 18776
rect 506584 16574 506612 18770
rect 506584 16546 507256 16574
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 354 507256 16546
rect 507872 10334 507900 59599
rect 509238 59392 509294 59401
rect 509238 59327 509294 59336
rect 510710 59392 510766 59401
rect 510710 59327 510766 59336
rect 509252 46578 509280 59327
rect 509240 46572 509292 46578
rect 509240 46514 509292 46520
rect 510724 43654 510752 59327
rect 510816 55214 510844 59622
rect 511998 59528 512054 59537
rect 511998 59463 512054 59472
rect 510816 55186 510936 55214
rect 510712 43648 510764 43654
rect 510712 43590 510764 43596
rect 510908 40934 510936 55186
rect 510896 40928 510948 40934
rect 510896 40870 510948 40876
rect 509240 39568 509292 39574
rect 509240 39510 509292 39516
rect 509252 16574 509280 39510
rect 512012 39506 512040 59463
rect 513470 59392 513526 59401
rect 513470 59327 513526 59336
rect 513380 46436 513432 46442
rect 513380 46378 513432 46384
rect 512000 39500 512052 39506
rect 512000 39442 512052 39448
rect 510620 18760 510672 18766
rect 510620 18702 510672 18708
rect 510632 16574 510660 18702
rect 509252 16546 509648 16574
rect 510632 16546 511304 16574
rect 507860 10328 507912 10334
rect 507860 10270 507912 10276
rect 508872 5228 508924 5234
rect 508872 5170 508924 5176
rect 508884 480 508912 5170
rect 507646 354 507758 480
rect 507228 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 511276 480 511304 16546
rect 512460 5160 512512 5166
rect 512460 5102 512512 5108
rect 512472 480 512500 5102
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513392 354 513420 46378
rect 513484 38146 513512 59327
rect 514760 51808 514812 51814
rect 514760 51750 514812 51756
rect 513472 38140 513524 38146
rect 513472 38082 513524 38088
rect 514772 480 514800 51750
rect 514864 13122 514892 59706
rect 515034 59528 515090 59537
rect 515034 59463 515090 59472
rect 515048 49162 515076 59463
rect 515968 59401 515996 59735
rect 516138 59664 516194 59673
rect 516138 59599 516194 59608
rect 515954 59392 516010 59401
rect 515954 59327 516010 59336
rect 516152 51950 516180 59599
rect 517610 59392 517666 59401
rect 517610 59327 517666 59336
rect 516140 51944 516192 51950
rect 516140 51886 516192 51892
rect 515036 49156 515088 49162
rect 515036 49098 515088 49104
rect 516140 43580 516192 43586
rect 516140 43522 516192 43528
rect 516152 16574 516180 43522
rect 517520 18692 517572 18698
rect 517520 18634 517572 18640
rect 516152 16546 517192 16574
rect 514852 13116 514904 13122
rect 514852 13058 514904 13064
rect 515956 5092 516008 5098
rect 515956 5034 516008 5040
rect 515968 480 515996 5034
rect 516784 4888 516836 4894
rect 516784 4830 516836 4836
rect 516796 4758 516824 4830
rect 516784 4752 516836 4758
rect 516784 4694 516836 4700
rect 517164 480 517192 16546
rect 517532 2774 517560 18634
rect 517624 9382 517652 59327
rect 517612 9376 517664 9382
rect 517612 9318 517664 9324
rect 519004 9314 519032 59735
rect 519082 59528 519138 59537
rect 519138 59486 519216 59514
rect 519082 59463 519138 59472
rect 518992 9308 519044 9314
rect 518992 9250 519044 9256
rect 519188 9246 519216 59486
rect 520108 59401 520136 59735
rect 522040 59537 522068 59735
rect 522118 59664 522174 59673
rect 522118 59599 522174 59608
rect 520370 59528 520426 59537
rect 520370 59463 520426 59472
rect 522026 59528 522082 59537
rect 522026 59463 522082 59472
rect 520094 59392 520150 59401
rect 520094 59327 520150 59336
rect 520280 49224 520332 49230
rect 520280 49166 520332 49172
rect 519176 9240 519228 9246
rect 519176 9182 519228 9188
rect 519544 5024 519596 5030
rect 519544 4966 519596 4972
rect 517532 2746 517928 2774
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 354 517928 2746
rect 519556 480 519584 4966
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 49166
rect 520384 9178 520412 59463
rect 522132 59401 522160 59599
rect 523038 59528 523094 59537
rect 523038 59463 523094 59472
rect 521750 59392 521806 59401
rect 521750 59327 521806 59336
rect 522118 59392 522174 59401
rect 522118 59327 522174 59336
rect 521660 18624 521712 18630
rect 521660 18566 521712 18572
rect 520372 9172 520424 9178
rect 520372 9114 520424 9120
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 18566
rect 521764 9110 521792 59327
rect 523052 53310 523080 59463
rect 524248 59401 524276 59735
rect 525300 59735 525302 59744
rect 527364 59764 527416 59770
rect 525248 59706 525300 59712
rect 528650 59735 528706 59744
rect 533710 59800 533766 59809
rect 537666 59800 537722 59809
rect 533710 59735 533712 59744
rect 527364 59706 527416 59712
rect 524510 59664 524566 59673
rect 524510 59599 524566 59608
rect 523222 59392 523278 59401
rect 523222 59327 523278 59336
rect 524234 59392 524290 59401
rect 524234 59327 524290 59336
rect 523040 53304 523092 53310
rect 523040 53246 523092 53252
rect 523040 47728 523092 47734
rect 523040 47670 523092 47676
rect 521752 9104 521804 9110
rect 521752 9046 521804 9052
rect 523052 7546 523080 47670
rect 523236 36786 523264 59327
rect 524420 58744 524472 58750
rect 524420 58686 524472 58692
rect 523224 36780 523276 36786
rect 523224 36722 523276 36728
rect 523132 17264 523184 17270
rect 523132 17206 523184 17212
rect 523040 7540 523092 7546
rect 523040 7482 523092 7488
rect 523144 2774 523172 17206
rect 523868 7540 523920 7546
rect 523868 7482 523920 7488
rect 523052 2746 523172 2774
rect 523052 480 523080 2746
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523880 354 523908 7482
rect 524432 6914 524460 58686
rect 524524 9042 524552 59599
rect 525798 59256 525854 59265
rect 525798 59191 525854 59200
rect 527178 59256 527234 59265
rect 527178 59191 527234 59200
rect 524512 9036 524564 9042
rect 524512 8978 524564 8984
rect 525812 8974 525840 59191
rect 527192 54602 527220 59191
rect 527180 54596 527232 54602
rect 527180 54538 527232 54544
rect 527180 38072 527232 38078
rect 527180 38014 527232 38020
rect 527192 16574 527220 38014
rect 527376 32570 527404 59706
rect 528558 59392 528614 59401
rect 528558 59327 528614 59336
rect 527364 32564 527416 32570
rect 527364 32506 527416 32512
rect 528572 27062 528600 59327
rect 528664 57254 528692 59735
rect 533764 59735 533766 59744
rect 535644 59764 535696 59770
rect 533712 59706 533764 59712
rect 544934 59800 544990 59809
rect 537666 59735 537668 59744
rect 535644 59706 535696 59712
rect 537720 59735 537722 59744
rect 539784 59764 539836 59770
rect 537668 59706 537720 59712
rect 544934 59735 544990 59744
rect 546958 59800 547014 59809
rect 546958 59735 547014 59744
rect 547694 59800 547750 59809
rect 547694 59735 547750 59744
rect 554318 59800 554374 59809
rect 556618 59800 556674 59809
rect 554318 59735 554320 59744
rect 539784 59706 539836 59712
rect 535550 59664 535606 59673
rect 535550 59599 535606 59608
rect 529018 59528 529074 59537
rect 529018 59463 529074 59472
rect 532698 59528 532754 59537
rect 532698 59463 532754 59472
rect 529032 58818 529060 59463
rect 529938 59392 529994 59401
rect 529938 59327 529994 59336
rect 529020 58812 529072 58818
rect 529020 58754 529072 58760
rect 528652 57248 528704 57254
rect 528652 57190 528704 57196
rect 528560 27056 528612 27062
rect 528560 26998 528612 27004
rect 528560 24200 528612 24206
rect 528560 24142 528612 24148
rect 527192 16546 527864 16574
rect 525800 8968 525852 8974
rect 525800 8910 525852 8916
rect 524432 6886 525472 6914
rect 525444 480 525472 6886
rect 526628 4956 526680 4962
rect 526628 4898 526680 4904
rect 526640 480 526668 4898
rect 527836 480 527864 16546
rect 524206 354 524318 480
rect 523880 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528572 354 528600 24142
rect 529952 22914 529980 59327
rect 530584 53168 530636 53174
rect 530584 53110 530636 53116
rect 529940 22908 529992 22914
rect 529940 22850 529992 22856
rect 530124 4752 530176 4758
rect 530124 4694 530176 4700
rect 530136 480 530164 4694
rect 530596 3058 530624 53110
rect 531412 50584 531464 50590
rect 531412 50526 531464 50532
rect 531424 6914 531452 50526
rect 532712 35290 532740 59463
rect 535564 59401 535592 59599
rect 534078 59392 534134 59401
rect 534078 59327 534134 59336
rect 535550 59392 535606 59401
rect 535550 59327 535606 59336
rect 532700 35284 532752 35290
rect 532700 35226 532752 35232
rect 534092 33930 534120 59327
rect 534080 33924 534132 33930
rect 534080 33866 534132 33872
rect 535460 29640 535512 29646
rect 535460 29582 535512 29588
rect 534448 14748 534500 14754
rect 534448 14690 534500 14696
rect 531332 6886 531452 6914
rect 530584 3052 530636 3058
rect 530584 2994 530636 3000
rect 531332 480 531360 6886
rect 533712 4820 533764 4826
rect 533712 4762 533764 4768
rect 532516 3052 532568 3058
rect 532516 2994 532568 3000
rect 532528 480 532556 2994
rect 533724 480 533752 4762
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 528990 -960 529102 326
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534460 354 534488 14690
rect 535472 6914 535500 29582
rect 535656 8022 535684 59706
rect 535826 59528 535882 59537
rect 535826 59463 535882 59472
rect 535644 8016 535696 8022
rect 535644 7958 535696 7964
rect 535840 7954 535868 59463
rect 536838 59392 536894 59401
rect 538310 59392 538366 59401
rect 536894 59350 536972 59378
rect 536838 59327 536894 59336
rect 536840 58948 536892 58954
rect 536840 58890 536892 58896
rect 536852 16574 536880 58890
rect 536944 31210 536972 59350
rect 538310 59327 538366 59336
rect 539598 59392 539654 59401
rect 539598 59327 539654 59336
rect 536932 31204 536984 31210
rect 536932 31146 536984 31152
rect 536852 16546 537248 16574
rect 535828 7948 535880 7954
rect 535828 7890 535880 7896
rect 535472 6886 536144 6914
rect 536116 480 536144 6886
rect 537220 480 537248 16546
rect 538220 14680 538272 14686
rect 538220 14622 538272 14628
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 14622
rect 538324 7886 538352 59327
rect 538864 28280 538916 28286
rect 538864 28222 538916 28228
rect 538312 7880 538364 7886
rect 538312 7822 538364 7828
rect 538876 3534 538904 28222
rect 539612 7750 539640 59327
rect 539796 7818 539824 59706
rect 540794 59664 540850 59673
rect 540794 59599 540850 59608
rect 541806 59664 541862 59673
rect 541806 59599 541808 59608
rect 540808 59401 540836 59599
rect 541860 59599 541862 59608
rect 544016 59628 544068 59634
rect 541808 59570 541860 59576
rect 544016 59570 544068 59576
rect 541070 59528 541126 59537
rect 541070 59463 541126 59472
rect 543830 59528 543886 59537
rect 543830 59463 543886 59472
rect 540794 59392 540850 59401
rect 540794 59327 540850 59336
rect 539876 28416 539928 28422
rect 539876 28358 539928 28364
rect 539888 16574 539916 28358
rect 539888 16546 540376 16574
rect 539784 7812 539836 7818
rect 539784 7754 539836 7760
rect 539600 7744 539652 7750
rect 539600 7686 539652 7692
rect 538864 3528 538916 3534
rect 538864 3470 538916 3476
rect 539600 3528 539652 3534
rect 539600 3470 539652 3476
rect 539612 480 539640 3470
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540348 354 540376 16546
rect 541084 7682 541112 59463
rect 542450 59392 542506 59401
rect 542450 59327 542506 59336
rect 542360 33856 542412 33862
rect 542360 33798 542412 33804
rect 542372 16574 542400 33798
rect 542464 29714 542492 59327
rect 543844 50522 543872 59463
rect 543832 50516 543884 50522
rect 543832 50458 543884 50464
rect 543740 29776 543792 29782
rect 543740 29718 543792 29724
rect 542452 29708 542504 29714
rect 542452 29650 542504 29656
rect 543752 16574 543780 29718
rect 544028 28354 544056 59570
rect 544948 59401 544976 59735
rect 546972 59537 547000 59735
rect 545118 59528 545174 59537
rect 545118 59463 545174 59472
rect 546958 59528 547014 59537
rect 546958 59463 547014 59472
rect 544934 59392 544990 59401
rect 544934 59327 544990 59336
rect 545132 51746 545160 59463
rect 547708 59401 547736 59735
rect 554372 59735 554374 59744
rect 556344 59764 556396 59770
rect 554320 59706 554372 59712
rect 556618 59735 556674 59744
rect 560390 59800 560446 59809
rect 566646 59800 566702 59809
rect 560390 59735 560392 59744
rect 556344 59706 556396 59712
rect 547878 59664 547934 59673
rect 547878 59599 547934 59608
rect 550086 59664 550142 59673
rect 550086 59599 550142 59608
rect 553398 59664 553454 59673
rect 553398 59599 553454 59608
rect 546498 59392 546554 59401
rect 546498 59327 546554 59336
rect 547694 59392 547750 59401
rect 547694 59327 547750 59336
rect 545212 53372 545264 53378
rect 545212 53314 545264 53320
rect 545120 51740 545172 51746
rect 545120 51682 545172 51688
rect 544016 28348 544068 28354
rect 544016 28290 544068 28296
rect 545224 16574 545252 53314
rect 546512 49026 546540 59327
rect 546592 50448 546644 50454
rect 546592 50390 546644 50396
rect 546500 49020 546552 49026
rect 546500 48962 546552 48968
rect 546604 16574 546632 50390
rect 547892 47666 547920 59599
rect 547970 59528 548026 59537
rect 547970 59463 548026 59472
rect 547984 51074 548012 59463
rect 550100 59401 550128 59599
rect 550638 59528 550694 59537
rect 550638 59463 550694 59472
rect 552294 59528 552350 59537
rect 552294 59463 552350 59472
rect 549258 59392 549314 59401
rect 549258 59327 549314 59336
rect 550086 59392 550142 59401
rect 550086 59327 550142 59336
rect 549272 53106 549300 59327
rect 549260 53100 549312 53106
rect 549260 53042 549312 53048
rect 547984 51046 548104 51074
rect 547880 47660 547932 47666
rect 547880 47602 547932 47608
rect 547880 31136 547932 31142
rect 547880 31078 547932 31084
rect 547144 31068 547196 31074
rect 547144 31010 547196 31016
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 545224 16546 545528 16574
rect 546604 16546 546724 16574
rect 541992 14612 542044 14618
rect 541992 14554 542044 14560
rect 541072 7676 541124 7682
rect 541072 7618 541124 7624
rect 542004 480 542032 14554
rect 540766 354 540878 480
rect 540348 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545500 480 545528 16546
rect 546696 480 546724 16546
rect 547156 4010 547184 31010
rect 547144 4004 547196 4010
rect 547144 3946 547196 3952
rect 547892 480 547920 31078
rect 548076 25702 548104 51046
rect 550652 46238 550680 59463
rect 552110 59392 552166 59401
rect 552110 59327 552166 59336
rect 550640 46232 550692 46238
rect 550640 46174 550692 46180
rect 552124 43518 552152 59327
rect 552112 43512 552164 43518
rect 552112 43454 552164 43460
rect 552308 42090 552336 59463
rect 552296 42084 552348 42090
rect 552296 42026 552348 42032
rect 552020 36712 552072 36718
rect 552020 36654 552072 36660
rect 550640 33992 550692 33998
rect 550640 33934 550692 33940
rect 548064 25696 548116 25702
rect 548064 25638 548116 25644
rect 550652 16574 550680 33934
rect 552032 16574 552060 36654
rect 553412 24138 553440 59599
rect 554778 59392 554834 59401
rect 554778 59327 554834 59336
rect 554792 40730 554820 59327
rect 556160 54664 556212 54670
rect 556160 54606 556212 54612
rect 554780 40724 554832 40730
rect 554780 40666 554832 40672
rect 554780 35352 554832 35358
rect 554780 35294 554832 35300
rect 553492 25628 553544 25634
rect 553492 25570 553544 25576
rect 553400 24132 553452 24138
rect 553400 24074 553452 24080
rect 553504 16574 553532 25570
rect 550652 16546 551048 16574
rect 552032 16546 552704 16574
rect 553504 16546 553808 16574
rect 548616 14544 548668 14550
rect 548616 14486 548668 14492
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 548628 354 548656 14486
rect 550272 4004 550324 4010
rect 550272 3946 550324 3952
rect 550284 480 550312 3946
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 552676 480 552704 16546
rect 553780 480 553808 16546
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 35294
rect 556172 480 556200 54606
rect 556356 39370 556384 59706
rect 556526 59528 556582 59537
rect 556526 59463 556582 59472
rect 556344 39364 556396 39370
rect 556344 39306 556396 39312
rect 556540 37942 556568 59463
rect 556632 54534 556660 59735
rect 560444 59735 560446 59744
rect 561772 59764 561824 59770
rect 560392 59706 560444 59712
rect 567014 59800 567070 59809
rect 566702 59758 567014 59786
rect 566646 59735 566702 59744
rect 567014 59735 567070 59744
rect 567290 59800 567346 59809
rect 567290 59735 567346 59744
rect 561772 59706 561824 59712
rect 561494 59664 561550 59673
rect 561494 59599 561496 59608
rect 561548 59599 561550 59608
rect 561496 59570 561548 59576
rect 560574 59528 560630 59537
rect 560574 59463 560630 59472
rect 560390 59392 560446 59401
rect 560390 59327 560446 59336
rect 557630 59256 557686 59265
rect 557630 59191 557686 59200
rect 557540 57316 557592 57322
rect 557540 57258 557592 57264
rect 556620 54528 556672 54534
rect 556620 54470 556672 54476
rect 556528 37936 556580 37942
rect 556528 37878 556580 37884
rect 556252 20324 556304 20330
rect 556252 20266 556304 20272
rect 556264 16574 556292 20266
rect 557552 16574 557580 57258
rect 557644 36582 557672 59191
rect 557632 36576 557684 36582
rect 557632 36518 557684 36524
rect 560404 32434 560432 59327
rect 560392 32428 560444 32434
rect 560392 32370 560444 32376
rect 560588 26926 560616 59463
rect 561680 55956 561732 55962
rect 561680 55898 561732 55904
rect 560576 26920 560628 26926
rect 560576 26862 560628 26868
rect 560300 20256 560352 20262
rect 560300 20198 560352 20204
rect 560312 16574 560340 20198
rect 561692 16574 561720 55898
rect 561784 25566 561812 59706
rect 563060 59628 563112 59634
rect 563060 59570 563112 59576
rect 561862 59528 561918 59537
rect 561862 59463 561918 59472
rect 561876 58682 561904 59463
rect 561864 58676 561916 58682
rect 561864 58618 561916 58624
rect 563072 35222 563100 59570
rect 565818 59528 565874 59537
rect 565818 59463 565874 59472
rect 564622 59392 564678 59401
rect 564622 59327 564678 59336
rect 563060 35216 563112 35222
rect 563060 35158 563112 35164
rect 564636 33794 564664 59327
rect 565832 47598 565860 59463
rect 567198 59392 567254 59401
rect 567198 59327 567254 59336
rect 567212 50386 567240 59327
rect 567304 55894 567332 59735
rect 571338 59528 571394 59537
rect 571338 59463 571394 59472
rect 569958 59392 570014 59401
rect 569958 59327 570014 59336
rect 568854 59256 568910 59265
rect 568854 59191 568910 59200
rect 567292 55888 567344 55894
rect 567292 55830 567344 55836
rect 567200 50380 567252 50386
rect 567200 50322 567252 50328
rect 565820 47592 565872 47598
rect 565820 47534 565872 47540
rect 566464 43444 566516 43450
rect 566464 43386 566516 43392
rect 564624 33788 564676 33794
rect 564624 33730 564676 33736
rect 563060 32496 563112 32502
rect 563060 32438 563112 32444
rect 561772 25560 561824 25566
rect 561772 25502 561824 25508
rect 556264 16546 556936 16574
rect 557552 16546 558592 16574
rect 560312 16546 560432 16574
rect 561692 16546 562088 16574
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558564 480 558592 16546
rect 559288 14476 559340 14482
rect 559288 14418 559340 14424
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 14418
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 562060 480 562088 16546
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 32438
rect 565820 26988 565872 26994
rect 565820 26930 565872 26936
rect 564440 21412 564492 21418
rect 564440 21354 564492 21360
rect 564452 3534 564480 21354
rect 564532 20188 564584 20194
rect 564532 20130 564584 20136
rect 564440 3528 564492 3534
rect 564440 3470 564492 3476
rect 564544 3346 564572 20130
rect 565832 16574 565860 26930
rect 565832 16546 566412 16574
rect 565268 3528 565320 3534
rect 565268 3470 565320 3476
rect 566384 3482 566412 16546
rect 566476 4146 566504 43386
rect 568868 7614 568896 59191
rect 569972 44878 570000 59327
rect 569960 44872 570012 44878
rect 569960 44814 570012 44820
rect 569960 22840 570012 22846
rect 569960 22782 570012 22788
rect 569972 16574 570000 22782
rect 571352 22778 571380 59463
rect 572720 58880 572772 58886
rect 572720 58822 572772 58828
rect 571340 22772 571392 22778
rect 571340 22714 571392 22720
rect 571340 20120 571392 20126
rect 571340 20062 571392 20068
rect 569972 16546 570368 16574
rect 568856 7608 568908 7614
rect 568856 7550 568908 7556
rect 569132 6316 569184 6322
rect 569132 6258 569184 6264
rect 566464 4140 566516 4146
rect 566464 4082 566516 4088
rect 568028 4140 568080 4146
rect 568028 4082 568080 4088
rect 564452 3318 564572 3346
rect 564452 480 564480 3318
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565280 354 565308 3470
rect 566384 3454 566872 3482
rect 566844 480 566872 3454
rect 568040 480 568068 4082
rect 569144 480 569172 6258
rect 570340 480 570368 16546
rect 565606 354 565718 480
rect 565280 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571352 354 571380 20062
rect 572732 16574 572760 58822
rect 576124 31272 576176 31278
rect 576124 31214 576176 31220
rect 574100 20052 574152 20058
rect 574100 19994 574152 20000
rect 574112 16574 574140 19994
rect 572732 16546 573496 16574
rect 574112 16546 575152 16574
rect 572720 6248 572772 6254
rect 572720 6190 572772 6196
rect 572732 480 572760 6190
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573468 354 573496 16546
rect 575124 480 575152 16546
rect 576136 4146 576164 31214
rect 578240 19984 578292 19990
rect 578240 19926 578292 19932
rect 578252 16574 578280 19926
rect 578252 16546 578648 16574
rect 576308 6180 576360 6186
rect 576308 6122 576360 6128
rect 576124 4140 576176 4146
rect 576124 4082 576176 4088
rect 576320 480 576348 6122
rect 577412 4140 577464 4146
rect 577412 4082 577464 4088
rect 577424 480 577452 4082
rect 578620 480 578648 16546
rect 581000 3596 581052 3602
rect 581000 3538 581052 3544
rect 581012 480 581040 3538
rect 582196 3460 582248 3466
rect 582196 3402 582248 3408
rect 582208 480 582236 3402
rect 583390 3360 583446 3369
rect 583390 3295 583446 3304
rect 583404 480 583432 3295
rect 573886 354 573998 480
rect 573468 326 573998 354
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 57610 387640 57666 387696
rect 60646 59744 60702 59800
rect 60554 59628 60610 59664
rect 60554 59608 60556 59628
rect 60556 59608 60608 59628
rect 60608 59608 60610 59628
rect 57794 59492 57850 59528
rect 57794 59472 57796 59492
rect 57796 59472 57848 59492
rect 57848 59472 57850 59492
rect 62302 59608 62358 59664
rect 61382 59472 61438 59528
rect 64510 59472 64566 59528
rect 58162 59372 58164 59392
rect 58164 59372 58216 59392
rect 58216 59372 58218 59392
rect 58162 59336 58218 59372
rect 60646 59336 60702 59392
rect 19430 3304 19486 3360
rect 62762 59336 62818 59392
rect 66442 59744 66498 59800
rect 67546 59608 67602 59664
rect 64694 59336 64750 59392
rect 65982 59336 66038 59392
rect 66166 59336 66222 59392
rect 68650 59472 68706 59528
rect 70582 59744 70638 59800
rect 71594 59744 71650 59800
rect 74722 59764 74778 59800
rect 74722 59744 74724 59764
rect 74724 59744 74776 59764
rect 74776 59744 74778 59764
rect 79874 59764 79930 59800
rect 79874 59744 79876 59764
rect 79876 59744 79928 59764
rect 79928 59744 79930 59764
rect 83002 59764 83058 59800
rect 83002 59744 83004 59764
rect 83004 59744 83056 59764
rect 83056 59744 83058 59764
rect 87418 59764 87474 59800
rect 87418 59744 87420 59764
rect 87420 59744 87472 59764
rect 87472 59744 87474 59764
rect 94502 59744 94558 59800
rect 97170 59744 97226 59800
rect 97538 59744 97594 59800
rect 98458 59744 98514 59800
rect 104806 59744 104862 59800
rect 71686 59608 71742 59664
rect 68834 59336 68890 59392
rect 70122 59336 70178 59392
rect 70306 59336 70362 59392
rect 71594 59336 71650 59392
rect 72882 59472 72938 59528
rect 75826 59608 75882 59664
rect 74446 59336 74502 59392
rect 77206 59472 77262 59528
rect 77022 59336 77078 59392
rect 79874 59608 79930 59664
rect 80886 59472 80942 59528
rect 83462 59472 83518 59528
rect 82082 59336 82138 59392
rect 84842 59336 84898 59392
rect 85486 59200 85542 59256
rect 87602 59608 87658 59664
rect 91282 59628 91338 59664
rect 91282 59608 91284 59628
rect 91284 59608 91336 59628
rect 91336 59608 91338 59628
rect 88982 59472 89038 59528
rect 93306 59608 93362 59664
rect 94318 59608 94374 59664
rect 93306 59472 93362 59528
rect 90362 59336 90418 59392
rect 91742 59336 91798 59392
rect 92938 59336 92994 59392
rect 93122 59336 93178 59392
rect 97814 59608 97870 59664
rect 94502 59472 94558 59528
rect 95882 59472 95938 59528
rect 97630 59472 97686 59528
rect 94318 59336 94374 59392
rect 94502 59336 94558 59392
rect 93122 3304 93178 3360
rect 104714 59608 104770 59664
rect 98458 59472 98514 59528
rect 99286 59336 99342 59392
rect 100666 59200 100722 59256
rect 102598 59472 102654 59528
rect 102230 59336 102286 59392
rect 103426 59356 103482 59392
rect 103426 59336 103428 59356
rect 103428 59336 103480 59356
rect 103480 59336 103482 59356
rect 105726 59472 105782 59528
rect 104806 59336 104862 59392
rect 105542 59336 105598 59392
rect 108210 59744 108266 59800
rect 112534 59744 112590 59800
rect 108302 59608 108358 59664
rect 110878 59608 110934 59664
rect 112442 59608 112498 59664
rect 106922 59336 106978 59392
rect 107934 59336 107990 59392
rect 109682 59472 109738 59528
rect 111062 59336 111118 59392
rect 120262 59764 120318 59800
rect 120262 59744 120264 59764
rect 120264 59744 120316 59764
rect 120316 59744 120318 59764
rect 121274 59744 121330 59800
rect 118146 59628 118202 59664
rect 118146 59608 118148 59628
rect 118148 59608 118200 59628
rect 118200 59608 118202 59628
rect 113822 59472 113878 59528
rect 112534 59336 112590 59392
rect 116122 59492 116178 59528
rect 116122 59472 116124 59492
rect 116124 59472 116176 59492
rect 116176 59472 116178 59492
rect 115202 59336 115258 59392
rect 118146 59472 118202 59528
rect 120906 59608 120962 59664
rect 119342 59336 119398 59392
rect 120722 59336 120778 59392
rect 125414 59628 125470 59664
rect 125414 59608 125416 59628
rect 125416 59608 125468 59628
rect 125468 59608 125470 59628
rect 121274 59472 121330 59528
rect 122102 59336 122158 59392
rect 122838 59336 122894 59392
rect 123114 59200 123170 59256
rect 128450 59744 128506 59800
rect 131578 59764 131634 59800
rect 131578 59744 131580 59764
rect 131580 59744 131632 59764
rect 131632 59744 131634 59764
rect 137834 59764 137890 59800
rect 137834 59744 137836 59764
rect 137836 59744 137888 59764
rect 137888 59744 137890 59764
rect 138938 59744 138994 59800
rect 125414 59472 125470 59528
rect 128082 59472 128138 59528
rect 124862 59200 124918 59256
rect 126242 59336 126298 59392
rect 127714 59200 127770 59256
rect 129186 59472 129242 59528
rect 130382 59336 130438 59392
rect 132590 59608 132646 59664
rect 133142 59472 133198 59528
rect 133326 59336 133382 59392
rect 134522 59200 134578 59256
rect 137834 59608 137890 59664
rect 137466 59472 137522 59528
rect 137282 59336 137338 59392
rect 141974 59764 142030 59800
rect 141974 59744 141976 59764
rect 141976 59744 142028 59764
rect 142028 59744 142030 59764
rect 145010 59764 145066 59800
rect 145010 59744 145012 59764
rect 145012 59744 145064 59764
rect 145064 59744 145066 59764
rect 148138 59764 148194 59800
rect 148138 59744 148140 59764
rect 148140 59744 148192 59764
rect 148192 59744 148194 59764
rect 150254 59744 150310 59800
rect 138938 59472 138994 59528
rect 137834 59336 137890 59392
rect 138662 59336 138718 59392
rect 141422 59472 141478 59528
rect 141606 59336 141662 59392
rect 145562 59472 145618 59528
rect 144182 59200 144238 59256
rect 149702 59608 149758 59664
rect 148322 59472 148378 59528
rect 146942 59336 146998 59392
rect 152278 59764 152334 59800
rect 152278 59744 152280 59764
rect 152280 59744 152332 59764
rect 152332 59744 152334 59764
rect 156602 59764 156658 59800
rect 156602 59744 156604 59764
rect 156604 59744 156656 59764
rect 156656 59744 156658 59764
rect 157430 59744 157486 59800
rect 159546 59744 159602 59800
rect 150254 59472 150310 59528
rect 151082 59336 151138 59392
rect 152462 59200 152518 59256
rect 154302 59608 154358 59664
rect 156602 59608 156658 59664
rect 154026 59472 154082 59528
rect 154302 59336 154358 59392
rect 155222 59336 155278 59392
rect 158626 59608 158682 59664
rect 157982 59472 158038 59528
rect 157430 59336 157486 59392
rect 162582 59764 162638 59800
rect 162582 59744 162584 59764
rect 162584 59744 162636 59764
rect 162636 59744 162638 59764
rect 165710 59744 165766 59800
rect 170954 59744 171010 59800
rect 178222 59744 178278 59800
rect 159546 59472 159602 59528
rect 159362 59336 159418 59392
rect 164882 59608 164938 59664
rect 162582 59472 162638 59528
rect 162582 59336 162638 59392
rect 164146 59200 164202 59256
rect 170862 59608 170918 59664
rect 166814 59472 166870 59528
rect 165710 59336 165766 59392
rect 166630 59336 166686 59392
rect 168286 59200 168342 59256
rect 166814 3304 166870 3360
rect 177118 59492 177174 59528
rect 177118 59472 177120 59492
rect 177120 59472 177172 59492
rect 177172 59472 177174 59492
rect 172426 59336 172482 59392
rect 173806 59200 173862 59256
rect 174910 59064 174966 59120
rect 176566 59336 176622 59392
rect 178130 59608 178186 59664
rect 181258 59764 181314 59800
rect 181258 59744 181260 59764
rect 181260 59744 181312 59764
rect 181312 59744 181314 59764
rect 190550 59764 190606 59800
rect 190550 59744 190552 59764
rect 190552 59744 190604 59764
rect 190604 59744 190606 59764
rect 195794 59764 195850 59800
rect 195794 59744 195796 59764
rect 195796 59744 195848 59764
rect 195848 59744 195850 59764
rect 196806 59744 196862 59800
rect 198830 59744 198886 59800
rect 179142 59472 179198 59528
rect 178222 59336 178278 59392
rect 182086 59608 182142 59664
rect 180706 59336 180762 59392
rect 183190 59472 183246 59528
rect 187422 59472 187478 59528
rect 183466 59336 183522 59392
rect 184846 59200 184902 59256
rect 187514 59336 187570 59392
rect 188986 59608 189042 59664
rect 190550 59608 190606 59664
rect 191470 59472 191526 59528
rect 193678 59492 193734 59528
rect 193678 59472 193680 59492
rect 193680 59472 193732 59492
rect 193732 59472 193734 59492
rect 193126 59336 193182 59392
rect 195794 59608 195850 59664
rect 195702 59472 195758 59528
rect 196806 59472 196862 59528
rect 198646 59472 198702 59528
rect 197266 59336 197322 59392
rect 208122 59764 208178 59800
rect 208122 59744 208124 59764
rect 208124 59744 208176 59764
rect 208176 59744 208178 59764
rect 209962 59744 210018 59800
rect 210330 59744 210386 59800
rect 211250 59744 211306 59800
rect 200026 59608 200082 59664
rect 199842 59472 199898 59528
rect 198830 59336 198886 59392
rect 206098 59492 206154 59528
rect 206098 59472 206100 59492
rect 206100 59472 206152 59492
rect 206152 59472 206154 59492
rect 201406 59336 201462 59392
rect 202786 59200 202842 59256
rect 205546 59336 205602 59392
rect 204074 59200 204130 59256
rect 208214 59608 208270 59664
rect 211066 59608 211122 59664
rect 208122 59472 208178 59528
rect 209686 59336 209742 59392
rect 222566 59764 222622 59800
rect 222566 59744 222568 59764
rect 222568 59744 222620 59764
rect 222620 59744 222622 59764
rect 223670 59744 223726 59800
rect 227902 59744 227958 59800
rect 238758 59744 238814 59800
rect 217966 59608 218022 59664
rect 219898 59608 219954 59664
rect 212262 59472 212318 59528
rect 216402 59472 216458 59528
rect 211250 59336 211306 59392
rect 212354 59336 212410 59392
rect 213826 59200 213882 59256
rect 216494 59336 216550 59392
rect 217874 59200 217930 59256
rect 219346 59472 219402 59528
rect 219898 59336 219954 59392
rect 223486 59608 223542 59664
rect 220634 59336 220690 59392
rect 222106 59200 222162 59256
rect 224682 59472 224738 59528
rect 223670 59336 223726 59392
rect 226706 59492 226762 59528
rect 226706 59472 226708 59492
rect 226708 59472 226760 59492
rect 226760 59472 226762 59492
rect 226246 59336 226302 59392
rect 227810 59608 227866 59664
rect 232962 59608 233018 59664
rect 229006 59472 229062 59528
rect 232870 59472 232926 59528
rect 227902 59336 227958 59392
rect 228822 59336 228878 59392
rect 230386 59336 230442 59392
rect 231766 59336 231822 59392
rect 244278 59764 244334 59800
rect 244278 59744 244280 59764
rect 244280 59744 244332 59764
rect 244332 59744 244334 59764
rect 246762 59744 246818 59800
rect 248418 59744 248474 59800
rect 252650 59744 252706 59800
rect 242714 59608 242770 59664
rect 234986 59492 235042 59528
rect 234986 59472 234988 59492
rect 234988 59472 235040 59492
rect 235040 59472 235042 59492
rect 238758 59472 238814 59528
rect 241334 59472 241390 59528
rect 232962 59336 233018 59392
rect 234526 59336 234582 59392
rect 238666 59336 238722 59392
rect 241242 59336 241298 59392
rect 235906 59200 235962 59256
rect 237194 59200 237250 59256
rect 237010 59064 237066 59120
rect 245474 59608 245530 59664
rect 244186 59472 244242 59528
rect 248326 59472 248382 59528
rect 249430 59472 249486 59528
rect 251546 59492 251602 59528
rect 251546 59472 251548 59492
rect 251548 59472 251600 59492
rect 251600 59472 251602 59492
rect 251086 59336 251142 59392
rect 252558 59608 252614 59664
rect 259826 59764 259882 59800
rect 259826 59744 259828 59764
rect 259828 59744 259880 59764
rect 259880 59744 259882 59764
rect 263966 59744 264022 59800
rect 266174 59744 266230 59800
rect 253662 59472 253718 59528
rect 252650 59336 252706 59392
rect 255686 59492 255742 59528
rect 255686 59472 255688 59492
rect 255688 59472 255740 59492
rect 255740 59472 255742 59492
rect 257802 59492 257858 59528
rect 257802 59472 257804 59492
rect 257804 59472 257856 59492
rect 257856 59472 257858 59492
rect 255226 59336 255282 59392
rect 257802 59336 257858 59392
rect 260746 59472 260802 59528
rect 259366 59200 259422 59256
rect 261942 59336 261998 59392
rect 266082 59608 266138 59664
rect 264242 59472 264298 59528
rect 262862 59200 262918 59256
rect 268106 59764 268162 59800
rect 268106 59744 268108 59764
rect 268108 59744 268160 59764
rect 268160 59744 268162 59764
rect 266174 59472 266230 59528
rect 270222 59608 270278 59664
rect 269946 59472 270002 59528
rect 267002 59336 267058 59392
rect 268382 59200 268438 59256
rect 269762 59200 269818 59256
rect 272522 59744 272578 59800
rect 275466 59744 275522 59800
rect 276386 59744 276442 59800
rect 272522 59608 272578 59664
rect 275374 59608 275430 59664
rect 270222 59336 270278 59392
rect 271142 59336 271198 59392
rect 272246 59336 272302 59392
rect 274086 59472 274142 59528
rect 273902 59336 273958 59392
rect 275466 59472 275522 59528
rect 280618 59764 280674 59800
rect 280618 59744 280620 59764
rect 280620 59744 280672 59764
rect 280672 59744 280674 59764
rect 289818 59764 289874 59800
rect 289818 59744 289820 59764
rect 289820 59744 289872 59764
rect 289872 59744 289874 59764
rect 292946 59764 293002 59800
rect 292946 59744 292948 59764
rect 292948 59744 293000 59764
rect 293000 59744 293002 59764
rect 297086 59764 297142 59800
rect 297086 59744 297088 59764
rect 297088 59744 297140 59764
rect 297140 59744 297142 59764
rect 302238 59764 302294 59800
rect 302238 59744 302240 59764
rect 302240 59744 302292 59764
rect 302292 59744 302294 59764
rect 306194 59744 306250 59800
rect 276386 59336 276442 59392
rect 276662 59200 276718 59256
rect 278226 59200 278282 59256
rect 278042 59064 278098 59120
rect 280802 59608 280858 59664
rect 286690 59628 286746 59664
rect 286690 59608 286692 59628
rect 286692 59608 286744 59628
rect 286744 59608 286746 59628
rect 282366 59472 282422 59528
rect 284666 59492 284722 59528
rect 284666 59472 284668 59492
rect 284668 59472 284720 59492
rect 284720 59472 284722 59492
rect 283562 59336 283618 59392
rect 286690 59472 286746 59528
rect 286322 59200 286378 59256
rect 290462 59472 290518 59528
rect 289082 59200 289138 59256
rect 293222 59472 293278 59528
rect 291842 59336 291898 59392
rect 299110 59608 299166 59664
rect 296074 59472 296130 59528
rect 298926 59472 298982 59528
rect 294786 59336 294842 59392
rect 295798 59336 295854 59392
rect 295982 59336 296038 59392
rect 297362 59200 297418 59256
rect 298742 59200 298798 59256
rect 299110 59336 299166 59392
rect 303342 59472 303398 59528
rect 301594 59200 301650 59256
rect 304906 59336 304962 59392
rect 310518 59764 310574 59800
rect 310518 59744 310520 59764
rect 310520 59744 310572 59764
rect 310572 59744 310574 59764
rect 318430 59744 318486 59800
rect 322202 59744 322258 59800
rect 326710 59764 326766 59800
rect 326710 59744 326712 59764
rect 326712 59744 326764 59764
rect 326764 59744 326766 59764
rect 306286 59336 306342 59392
rect 307574 59336 307630 59392
rect 307390 59064 307446 59120
rect 310426 59472 310482 59528
rect 311806 59472 311862 59528
rect 318062 59472 318118 59528
rect 311622 59336 311678 59392
rect 320454 59608 320510 59664
rect 322110 59608 322166 59664
rect 338026 59764 338082 59800
rect 338026 59744 338028 59764
rect 338028 59744 338080 59764
rect 338080 59744 338082 59764
rect 342166 59764 342222 59800
rect 342166 59744 342168 59764
rect 342168 59744 342220 59764
rect 342220 59744 342222 59764
rect 351182 59744 351238 59800
rect 318430 59336 318486 59392
rect 319442 59200 319498 59256
rect 321006 59472 321062 59528
rect 320822 59336 320878 59392
rect 328734 59628 328790 59664
rect 328734 59608 328736 59628
rect 328736 59608 328788 59628
rect 328788 59608 328790 59628
rect 324962 59336 325018 59392
rect 325698 59472 325754 59528
rect 328734 59472 328790 59528
rect 327722 59336 327778 59392
rect 333886 59608 333942 59664
rect 330850 59472 330906 59528
rect 331862 59472 331918 59528
rect 331862 59336 331918 59392
rect 331034 59200 331090 59256
rect 334622 59472 334678 59528
rect 337566 59472 337622 59528
rect 333242 59336 333298 59392
rect 333886 59336 333942 59392
rect 337382 59336 337438 59392
rect 335358 59200 335414 59256
rect 338762 59200 338818 59256
rect 341522 59472 341578 59528
rect 341706 59336 341762 59392
rect 342902 59200 342958 59256
rect 345294 59628 345350 59664
rect 345294 59608 345296 59628
rect 345296 59608 345348 59628
rect 345348 59608 345350 59628
rect 351182 59608 351238 59664
rect 345294 59472 345350 59528
rect 345846 59200 345902 59256
rect 347410 59472 347466 59528
rect 349802 59472 349858 59528
rect 348422 59336 348478 59392
rect 347410 59200 347466 59256
rect 349986 59336 350042 59392
rect 354678 59764 354734 59800
rect 354678 59744 354680 59764
rect 354680 59744 354732 59764
rect 354732 59744 354734 59764
rect 359462 59744 359518 59800
rect 353942 59472 353998 59528
rect 351458 59336 351514 59392
rect 352562 59336 352618 59392
rect 353298 59200 353354 59256
rect 355322 59200 355378 59256
rect 359462 59608 359518 59664
rect 358266 59472 358322 59528
rect 358082 59336 358138 59392
rect 360934 59744 360990 59800
rect 364246 59744 364302 59800
rect 371146 59744 371202 59800
rect 372158 59780 372160 59800
rect 372160 59780 372212 59800
rect 372212 59780 372214 59800
rect 372158 59744 372214 59780
rect 373722 59780 373724 59800
rect 373724 59780 373776 59800
rect 373776 59780 373778 59800
rect 373722 59744 373778 59780
rect 374182 59744 374238 59800
rect 376482 59744 376538 59800
rect 376758 59744 376814 59800
rect 384118 59744 384174 59800
rect 384486 59744 384542 59800
rect 388718 59744 388774 59800
rect 389086 59744 389142 59800
rect 392858 59764 392914 59800
rect 392858 59744 392860 59764
rect 392860 59744 392912 59764
rect 392912 59744 392914 59764
rect 359738 59472 359794 59528
rect 360842 59472 360898 59528
rect 362866 59608 362922 59664
rect 365902 59608 365958 59664
rect 363602 59472 363658 59528
rect 364246 59472 364302 59528
rect 365810 59472 365866 59528
rect 360934 59336 360990 59392
rect 362222 59336 362278 59392
rect 362866 59336 362922 59392
rect 362130 59200 362186 59256
rect 364982 59336 365038 59392
rect 367098 59472 367154 59528
rect 370134 59472 370190 59528
rect 367742 59336 367798 59392
rect 369950 59336 370006 59392
rect 371238 59608 371294 59664
rect 371146 59336 371202 59392
rect 373998 59336 374054 59392
rect 372710 59200 372766 59256
rect 376482 59472 376538 59528
rect 374274 59336 374330 59392
rect 378414 59608 378470 59664
rect 383750 59608 383806 59664
rect 378230 59472 378286 59528
rect 376850 59336 376906 59392
rect 382278 59472 382334 59528
rect 380990 59200 381046 59256
rect 382462 59336 382518 59392
rect 400126 59764 400182 59800
rect 400126 59744 400128 59764
rect 400128 59744 400180 59764
rect 400180 59744 400182 59764
rect 404174 59744 404230 59800
rect 409510 59764 409566 59800
rect 409510 59744 409512 59764
rect 409512 59744 409564 59764
rect 409564 59744 409566 59764
rect 390650 59608 390706 59664
rect 387890 59472 387946 59528
rect 385222 59372 385224 59392
rect 385224 59372 385276 59392
rect 385276 59372 385278 59392
rect 385222 59336 385278 59372
rect 386602 59336 386658 59392
rect 386418 59200 386474 59256
rect 389270 59200 389326 59256
rect 392030 59472 392086 59528
rect 394698 59472 394754 59528
rect 390834 59336 390890 59392
rect 393410 59336 393466 59392
rect 394790 59200 394846 59256
rect 399114 59472 399170 59528
rect 400218 59472 400274 59528
rect 398930 59336 398986 59392
rect 396078 59200 396134 59256
rect 403162 59472 403218 59528
rect 402978 59336 403034 59392
rect 412638 59764 412694 59800
rect 412638 59744 412640 59764
rect 412640 59744 412692 59764
rect 412692 59744 412694 59764
rect 418710 59764 418766 59800
rect 418710 59744 418712 59764
rect 418712 59744 418764 59764
rect 418764 59744 418766 59764
rect 423678 59744 423734 59800
rect 430118 59780 430120 59800
rect 430120 59780 430172 59800
rect 430172 59780 430174 59800
rect 430118 59744 430174 59780
rect 431498 59780 431500 59800
rect 431500 59780 431552 59800
rect 431552 59780 431554 59800
rect 431498 59744 431554 59780
rect 431958 59744 432014 59800
rect 433154 59744 433210 59800
rect 437478 59744 437534 59800
rect 437754 59744 437810 59800
rect 438858 59744 438914 59800
rect 444470 59744 444526 59800
rect 446678 59764 446734 59800
rect 446678 59744 446680 59764
rect 446680 59744 446732 59764
rect 446732 59744 446734 59764
rect 404266 59608 404322 59664
rect 404174 59336 404230 59392
rect 408590 59608 408646 59664
rect 405278 59492 405334 59528
rect 405278 59472 405280 59492
rect 405280 59472 405332 59492
rect 405332 59472 405334 59492
rect 407118 59472 407174 59528
rect 405830 59336 405886 59392
rect 409970 59200 410026 59256
rect 411442 59200 411498 59256
rect 413190 59472 413246 59528
rect 412638 59200 412694 59256
rect 416870 59472 416926 59528
rect 419630 59472 419686 59528
rect 415582 59336 415638 59392
rect 418250 59336 418306 59392
rect 420826 59492 420882 59528
rect 420826 59472 420828 59492
rect 420828 59472 420880 59492
rect 420880 59472 420882 59492
rect 421010 59200 421066 59256
rect 424966 59608 425022 59664
rect 423862 59472 423918 59528
rect 423770 59336 423826 59392
rect 425334 59472 425390 59528
rect 429198 59472 429254 59528
rect 428002 59336 428058 59392
rect 430670 59336 430726 59392
rect 432142 59472 432198 59528
rect 433246 59608 433302 59664
rect 433154 59336 433210 59392
rect 437386 59608 437442 59664
rect 434258 59472 434314 59528
rect 436190 59472 436246 59528
rect 434718 59336 434774 59392
rect 434258 59200 434314 59256
rect 436374 59336 436430 59392
rect 441066 59608 441122 59664
rect 454958 59764 455014 59800
rect 454958 59744 454960 59764
rect 454960 59744 455012 59764
rect 455012 59744 455014 59764
rect 457994 59744 458050 59800
rect 458362 59744 458418 59800
rect 459926 59744 459982 59800
rect 467286 59764 467342 59800
rect 467286 59744 467288 59764
rect 467288 59744 467340 59764
rect 467340 59744 467342 59764
rect 444562 59608 444618 59664
rect 448702 59608 448758 59664
rect 443550 59492 443606 59528
rect 443550 59472 443552 59492
rect 443552 59472 443604 59492
rect 443604 59472 443606 59492
rect 444470 59472 444526 59528
rect 441066 59336 441122 59392
rect 442262 59336 442318 59392
rect 443642 59336 443698 59392
rect 441066 59200 441122 59256
rect 440882 59064 440938 59120
rect 446402 59472 446458 59528
rect 449162 59472 449218 59528
rect 447782 59336 447838 59392
rect 448702 59336 448758 59392
rect 449714 59608 449770 59664
rect 454682 59472 454738 59528
rect 457442 59472 457498 59528
rect 453302 59336 453358 59392
rect 450542 59200 450598 59256
rect 453486 59064 453542 59120
rect 456062 59336 456118 59392
rect 458822 59200 458878 59256
rect 476026 59744 476082 59800
rect 484858 59744 484914 59800
rect 485778 59744 485834 59800
rect 488078 59780 488080 59800
rect 488080 59780 488132 59800
rect 488132 59780 488134 59800
rect 488078 59744 488134 59780
rect 489366 59780 489368 59800
rect 489368 59780 489420 59800
rect 489420 59780 489422 59800
rect 489366 59744 489422 59780
rect 490102 59744 490158 59800
rect 491022 59744 491078 59800
rect 495622 59744 495678 59800
rect 498474 59780 498476 59800
rect 498476 59780 498528 59800
rect 498528 59780 498530 59800
rect 498474 59744 498530 59780
rect 461122 59628 461178 59664
rect 461122 59608 461124 59628
rect 461124 59608 461176 59628
rect 461176 59608 461178 59628
rect 467102 59608 467158 59664
rect 461122 59472 461178 59528
rect 461122 59336 461178 59392
rect 463238 59472 463294 59528
rect 465722 59472 465778 59528
rect 464342 59336 464398 59392
rect 463238 59200 463294 59256
rect 465906 59336 465962 59392
rect 471978 59608 472034 59664
rect 473358 59608 473414 59664
rect 474554 59608 474610 59664
rect 470690 59472 470746 59528
rect 469862 59336 469918 59392
rect 469218 59200 469274 59256
rect 477590 59608 477646 59664
rect 474738 59472 474794 59528
rect 476026 59472 476082 59528
rect 473542 59336 473598 59392
rect 474554 59336 474610 59392
rect 476210 59336 476266 59392
rect 477590 59336 477646 59392
rect 480258 59608 480314 59664
rect 481638 59608 481694 59664
rect 482834 59608 482890 59664
rect 478878 59472 478934 59528
rect 483018 59472 483074 59528
rect 484858 59472 484914 59528
rect 481822 59336 481878 59392
rect 482834 59336 482890 59392
rect 485962 59608 486018 59664
rect 484490 59336 484546 59392
rect 485778 59336 485834 59392
rect 486146 59472 486202 59528
rect 489918 59472 489974 59528
rect 487250 59336 487306 59392
rect 488630 59336 488686 59392
rect 491114 59608 491170 59664
rect 491022 59336 491078 59392
rect 492126 59492 492182 59528
rect 492126 59472 492128 59492
rect 492128 59472 492180 59492
rect 492180 59472 492182 59492
rect 494058 59472 494114 59528
rect 492678 59336 492734 59392
rect 495530 59336 495586 59392
rect 498382 59608 498438 59664
rect 496818 59472 496874 59528
rect 508686 59744 508742 59800
rect 509054 59744 509110 59800
rect 512826 59764 512882 59800
rect 512826 59744 512828 59764
rect 512828 59744 512880 59764
rect 512880 59744 512882 59764
rect 515954 59744 516010 59800
rect 516966 59780 516968 59800
rect 516968 59780 517020 59800
rect 517020 59780 517022 59800
rect 516966 59744 517022 59780
rect 518346 59780 518348 59800
rect 518348 59780 518400 59800
rect 518400 59780 518402 59800
rect 518346 59744 518402 59780
rect 518990 59744 519046 59800
rect 520094 59744 520150 59800
rect 522026 59744 522082 59800
rect 524234 59744 524290 59800
rect 525246 59764 525302 59800
rect 525246 59744 525248 59764
rect 525248 59744 525300 59764
rect 525300 59744 525302 59764
rect 507858 59608 507914 59664
rect 510710 59608 510766 59664
rect 502706 59472 502762 59528
rect 504546 59492 504602 59528
rect 504546 59472 504548 59492
rect 504548 59472 504600 59492
rect 504600 59472 504602 59492
rect 502522 59336 502578 59392
rect 501050 59200 501106 59256
rect 506478 59472 506534 59528
rect 505190 59336 505246 59392
rect 503810 59200 503866 59256
rect 509238 59336 509294 59392
rect 510710 59336 510766 59392
rect 511998 59472 512054 59528
rect 513470 59336 513526 59392
rect 515034 59472 515090 59528
rect 516138 59608 516194 59664
rect 515954 59336 516010 59392
rect 517610 59336 517666 59392
rect 519082 59472 519138 59528
rect 522118 59608 522174 59664
rect 520370 59472 520426 59528
rect 522026 59472 522082 59528
rect 520094 59336 520150 59392
rect 523038 59472 523094 59528
rect 521750 59336 521806 59392
rect 522118 59336 522174 59392
rect 528650 59744 528706 59800
rect 533710 59764 533766 59800
rect 533710 59744 533712 59764
rect 533712 59744 533764 59764
rect 533764 59744 533766 59764
rect 524510 59608 524566 59664
rect 523222 59336 523278 59392
rect 524234 59336 524290 59392
rect 525798 59200 525854 59256
rect 527178 59200 527234 59256
rect 528558 59336 528614 59392
rect 537666 59764 537722 59800
rect 537666 59744 537668 59764
rect 537668 59744 537720 59764
rect 537720 59744 537722 59764
rect 544934 59744 544990 59800
rect 546958 59744 547014 59800
rect 547694 59744 547750 59800
rect 554318 59764 554374 59800
rect 554318 59744 554320 59764
rect 554320 59744 554372 59764
rect 554372 59744 554374 59764
rect 535550 59608 535606 59664
rect 529018 59472 529074 59528
rect 532698 59472 532754 59528
rect 529938 59336 529994 59392
rect 534078 59336 534134 59392
rect 535550 59336 535606 59392
rect 535826 59472 535882 59528
rect 536838 59336 536894 59392
rect 538310 59336 538366 59392
rect 539598 59336 539654 59392
rect 540794 59608 540850 59664
rect 541806 59628 541862 59664
rect 541806 59608 541808 59628
rect 541808 59608 541860 59628
rect 541860 59608 541862 59628
rect 541070 59472 541126 59528
rect 543830 59472 543886 59528
rect 540794 59336 540850 59392
rect 542450 59336 542506 59392
rect 545118 59472 545174 59528
rect 546958 59472 547014 59528
rect 544934 59336 544990 59392
rect 556618 59744 556674 59800
rect 560390 59764 560446 59800
rect 560390 59744 560392 59764
rect 560392 59744 560444 59764
rect 560444 59744 560446 59764
rect 547878 59608 547934 59664
rect 550086 59608 550142 59664
rect 553398 59608 553454 59664
rect 546498 59336 546554 59392
rect 547694 59336 547750 59392
rect 547970 59472 548026 59528
rect 550638 59472 550694 59528
rect 552294 59472 552350 59528
rect 549258 59336 549314 59392
rect 550086 59336 550142 59392
rect 552110 59336 552166 59392
rect 554778 59336 554834 59392
rect 556526 59472 556582 59528
rect 566646 59744 566702 59800
rect 567014 59744 567070 59800
rect 567290 59744 567346 59800
rect 561494 59628 561550 59664
rect 561494 59608 561496 59628
rect 561496 59608 561548 59628
rect 561548 59608 561550 59628
rect 560574 59472 560630 59528
rect 560390 59336 560446 59392
rect 557630 59200 557686 59256
rect 561862 59472 561918 59528
rect 565818 59472 565874 59528
rect 564622 59336 564678 59392
rect 567198 59336 567254 59392
rect 571338 59472 571394 59528
rect 569958 59336 570014 59392
rect 568854 59200 568910 59256
rect 583390 3304 583446 3360
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect 57605 387698 57671 387701
rect 57605 387696 59554 387698
rect 57605 387640 57610 387696
rect 57666 387654 59554 387696
rect 57666 387640 60076 387654
rect 57605 387638 60076 387640
rect 57605 387635 57671 387638
rect 59494 387594 60076 387638
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 57789 59530 57855 59533
rect 60384 59530 60444 60044
rect 60641 59802 60707 59805
rect 61120 59802 61180 60044
rect 60641 59800 61180 59802
rect 60641 59744 60646 59800
rect 60702 59744 61180 59800
rect 60641 59742 61180 59744
rect 60641 59739 60707 59742
rect 60549 59666 60615 59669
rect 62132 59666 62192 60044
rect 60549 59664 62192 59666
rect 60549 59608 60554 59664
rect 60610 59608 62192 59664
rect 60549 59606 62192 59608
rect 62297 59666 62363 59669
rect 63144 59666 63204 60044
rect 62297 59664 63204 59666
rect 62297 59608 62302 59664
rect 62358 59608 63204 59664
rect 62297 59606 63204 59608
rect 60549 59603 60615 59606
rect 62297 59603 62363 59606
rect 57789 59528 60444 59530
rect 57789 59472 57794 59528
rect 57850 59472 60444 59528
rect 57789 59470 60444 59472
rect 61377 59530 61443 59533
rect 64156 59530 64216 60044
rect 65260 59666 65320 60044
rect 61377 59528 64216 59530
rect 61377 59472 61382 59528
rect 61438 59472 64216 59528
rect 61377 59470 64216 59472
rect 64278 59606 65320 59666
rect 57789 59467 57855 59470
rect 61377 59467 61443 59470
rect 58157 59394 58223 59397
rect 60641 59394 60707 59397
rect 58157 59392 60707 59394
rect 58157 59336 58162 59392
rect 58218 59336 60646 59392
rect 60702 59336 60707 59392
rect 58157 59334 60707 59336
rect 58157 59331 58223 59334
rect 60641 59331 60707 59334
rect 62757 59394 62823 59397
rect 64278 59394 64338 59606
rect 64505 59530 64571 59533
rect 66272 59530 66332 60044
rect 67284 59938 67344 60044
rect 66486 59878 67344 59938
rect 66486 59805 66546 59878
rect 66437 59800 66546 59805
rect 68296 59802 68356 60044
rect 66437 59744 66442 59800
rect 66498 59744 66546 59800
rect 66437 59742 66546 59744
rect 67406 59742 68356 59802
rect 66437 59739 66503 59742
rect 64505 59528 66332 59530
rect 64505 59472 64510 59528
rect 64566 59472 66332 59528
rect 64505 59470 66332 59472
rect 64505 59467 64571 59470
rect 62757 59392 64338 59394
rect 62757 59336 62762 59392
rect 62818 59336 64338 59392
rect 62757 59334 64338 59336
rect 64689 59394 64755 59397
rect 65977 59394 66043 59397
rect 64689 59392 66043 59394
rect 64689 59336 64694 59392
rect 64750 59336 65982 59392
rect 66038 59336 66043 59392
rect 64689 59334 66043 59336
rect 62757 59331 62823 59334
rect 64689 59331 64755 59334
rect 65977 59331 66043 59334
rect 66161 59394 66227 59397
rect 67406 59394 67466 59742
rect 67541 59666 67607 59669
rect 69400 59666 69460 60044
rect 67541 59664 69460 59666
rect 67541 59608 67546 59664
rect 67602 59608 69460 59664
rect 67541 59606 69460 59608
rect 67541 59603 67607 59606
rect 68645 59530 68711 59533
rect 70412 59530 70472 60044
rect 70577 59802 70643 59805
rect 71424 59802 71484 60044
rect 70577 59800 71484 59802
rect 70577 59744 70582 59800
rect 70638 59744 71484 59800
rect 70577 59742 71484 59744
rect 71589 59802 71655 59805
rect 72436 59802 72496 60044
rect 71589 59800 72496 59802
rect 71589 59744 71594 59800
rect 71650 59744 72496 59800
rect 71589 59742 72496 59744
rect 70577 59739 70643 59742
rect 71589 59739 71655 59742
rect 71681 59666 71747 59669
rect 73540 59666 73600 60044
rect 71681 59664 73600 59666
rect 71681 59608 71686 59664
rect 71742 59608 73600 59664
rect 71681 59606 73600 59608
rect 71681 59603 71747 59606
rect 68645 59528 70472 59530
rect 68645 59472 68650 59528
rect 68706 59472 70472 59528
rect 68645 59470 70472 59472
rect 72877 59530 72943 59533
rect 74552 59530 74612 60044
rect 75564 59938 75624 60044
rect 74766 59878 75624 59938
rect 74766 59805 74826 59878
rect 74717 59800 74826 59805
rect 76576 59802 76636 60044
rect 74717 59744 74722 59800
rect 74778 59744 74826 59800
rect 74717 59742 74826 59744
rect 75686 59742 76636 59802
rect 74717 59739 74783 59742
rect 72877 59528 74612 59530
rect 72877 59472 72882 59528
rect 72938 59472 74612 59528
rect 72877 59470 74612 59472
rect 68645 59467 68711 59470
rect 72877 59467 72943 59470
rect 66161 59392 67466 59394
rect 66161 59336 66166 59392
rect 66222 59336 67466 59392
rect 66161 59334 67466 59336
rect 68829 59394 68895 59397
rect 70117 59394 70183 59397
rect 68829 59392 70183 59394
rect 68829 59336 68834 59392
rect 68890 59336 70122 59392
rect 70178 59336 70183 59392
rect 68829 59334 70183 59336
rect 66161 59331 66227 59334
rect 68829 59331 68895 59334
rect 70117 59331 70183 59334
rect 70301 59394 70367 59397
rect 71589 59394 71655 59397
rect 70301 59392 71655 59394
rect 70301 59336 70306 59392
rect 70362 59336 71594 59392
rect 71650 59336 71655 59392
rect 70301 59334 71655 59336
rect 70301 59331 70367 59334
rect 71589 59331 71655 59334
rect 74441 59394 74507 59397
rect 75686 59394 75746 59742
rect 75821 59666 75887 59669
rect 77680 59666 77740 60044
rect 75821 59664 77740 59666
rect 75821 59608 75826 59664
rect 75882 59608 77740 59664
rect 75821 59606 77740 59608
rect 75821 59603 75887 59606
rect 77201 59530 77267 59533
rect 78692 59530 78752 60044
rect 77201 59528 78752 59530
rect 77201 59472 77206 59528
rect 77262 59472 78752 59528
rect 77201 59470 78752 59472
rect 77201 59467 77267 59470
rect 74441 59392 75746 59394
rect 74441 59336 74446 59392
rect 74502 59336 75746 59392
rect 74441 59334 75746 59336
rect 77017 59394 77083 59397
rect 79704 59394 79764 60044
rect 79869 59802 79935 59805
rect 80716 59802 80776 60044
rect 79869 59800 80776 59802
rect 79869 59744 79874 59800
rect 79930 59744 80776 59800
rect 79869 59742 80776 59744
rect 79869 59739 79935 59742
rect 79869 59666 79935 59669
rect 81820 59666 81880 60044
rect 79869 59664 81880 59666
rect 79869 59608 79874 59664
rect 79930 59608 81880 59664
rect 79869 59606 81880 59608
rect 79869 59603 79935 59606
rect 80881 59530 80947 59533
rect 82832 59530 82892 60044
rect 82997 59802 83063 59805
rect 83844 59802 83904 60044
rect 82997 59800 83904 59802
rect 82997 59744 83002 59800
rect 83058 59744 83904 59800
rect 82997 59742 83904 59744
rect 82997 59739 83063 59742
rect 84856 59666 84916 60044
rect 80881 59528 82892 59530
rect 80881 59472 80886 59528
rect 80942 59472 82892 59528
rect 80881 59470 82892 59472
rect 83046 59606 84916 59666
rect 80881 59467 80947 59470
rect 77017 59392 79764 59394
rect 77017 59336 77022 59392
rect 77078 59336 79764 59392
rect 77017 59334 79764 59336
rect 82077 59394 82143 59397
rect 83046 59394 83106 59606
rect 83457 59530 83523 59533
rect 85960 59530 86020 60044
rect 83457 59528 86020 59530
rect 83457 59472 83462 59528
rect 83518 59472 86020 59528
rect 83457 59470 86020 59472
rect 83457 59467 83523 59470
rect 82077 59392 83106 59394
rect 82077 59336 82082 59392
rect 82138 59336 83106 59392
rect 82077 59334 83106 59336
rect 84837 59394 84903 59397
rect 86972 59394 87032 60044
rect 87984 59938 88044 60044
rect 84837 59392 87032 59394
rect 84837 59336 84842 59392
rect 84898 59336 87032 59392
rect 84837 59334 87032 59336
rect 87094 59878 88044 59938
rect 74441 59331 74507 59334
rect 77017 59331 77083 59334
rect 82077 59331 82143 59334
rect 84837 59331 84903 59334
rect 85481 59258 85547 59261
rect 87094 59258 87154 59878
rect 87413 59802 87479 59805
rect 88996 59802 89056 60044
rect 87413 59800 89056 59802
rect 87413 59744 87418 59800
rect 87474 59744 89056 59800
rect 87413 59742 89056 59744
rect 87413 59739 87479 59742
rect 87597 59666 87663 59669
rect 90008 59666 90068 60044
rect 87597 59664 90068 59666
rect 87597 59608 87602 59664
rect 87658 59608 90068 59664
rect 87597 59606 90068 59608
rect 87597 59603 87663 59606
rect 88977 59530 89043 59533
rect 91112 59530 91172 60044
rect 91277 59666 91343 59669
rect 92124 59666 92184 60044
rect 91277 59664 92184 59666
rect 91277 59608 91282 59664
rect 91338 59608 92184 59664
rect 91277 59606 92184 59608
rect 91277 59603 91343 59606
rect 93136 59530 93196 60044
rect 93301 59666 93367 59669
rect 94148 59666 94208 60044
rect 94497 59802 94563 59805
rect 95252 59802 95312 60044
rect 94497 59800 95312 59802
rect 94497 59744 94502 59800
rect 94558 59744 95312 59800
rect 94497 59742 95312 59744
rect 94497 59739 94563 59742
rect 93301 59664 94208 59666
rect 93301 59608 93306 59664
rect 93362 59608 94208 59664
rect 93301 59606 94208 59608
rect 94313 59666 94379 59669
rect 96264 59666 96324 60044
rect 97276 59938 97336 60044
rect 97276 59878 97458 59938
rect 97165 59802 97231 59805
rect 94313 59664 96324 59666
rect 94313 59608 94318 59664
rect 94374 59608 96324 59664
rect 94313 59606 96324 59608
rect 96478 59800 97231 59802
rect 96478 59744 97170 59800
rect 97226 59744 97231 59800
rect 96478 59742 97231 59744
rect 93301 59603 93367 59606
rect 94313 59603 94379 59606
rect 88977 59528 91172 59530
rect 88977 59472 88982 59528
rect 89038 59472 91172 59528
rect 88977 59470 91172 59472
rect 91326 59470 93196 59530
rect 93301 59530 93367 59533
rect 94497 59530 94563 59533
rect 93301 59528 94563 59530
rect 93301 59472 93306 59528
rect 93362 59472 94502 59528
rect 94558 59472 94563 59528
rect 93301 59470 94563 59472
rect 88977 59467 89043 59470
rect 90357 59394 90423 59397
rect 91326 59394 91386 59470
rect 93301 59467 93367 59470
rect 94497 59467 94563 59470
rect 95877 59530 95943 59533
rect 96478 59530 96538 59742
rect 97165 59739 97231 59742
rect 97398 59666 97458 59878
rect 97533 59802 97599 59805
rect 98288 59802 98348 60044
rect 97533 59800 98348 59802
rect 97533 59744 97538 59800
rect 97594 59744 98348 59800
rect 97533 59742 98348 59744
rect 98453 59802 98519 59805
rect 99392 59802 99452 60044
rect 98453 59800 99452 59802
rect 98453 59744 98458 59800
rect 98514 59744 99452 59800
rect 98453 59742 99452 59744
rect 97533 59739 97599 59742
rect 98453 59739 98519 59742
rect 95877 59528 96538 59530
rect 95877 59472 95882 59528
rect 95938 59472 96538 59528
rect 95877 59470 96538 59472
rect 97276 59606 97458 59666
rect 97809 59666 97875 59669
rect 100404 59666 100464 60044
rect 97809 59664 100464 59666
rect 97809 59608 97814 59664
rect 97870 59608 100464 59664
rect 97809 59606 100464 59608
rect 95877 59467 95943 59470
rect 90357 59392 91386 59394
rect 90357 59336 90362 59392
rect 90418 59336 91386 59392
rect 90357 59334 91386 59336
rect 91737 59394 91803 59397
rect 92933 59394 92999 59397
rect 91737 59392 92999 59394
rect 91737 59336 91742 59392
rect 91798 59336 92938 59392
rect 92994 59336 92999 59392
rect 91737 59334 92999 59336
rect 90357 59331 90423 59334
rect 91737 59331 91803 59334
rect 92933 59331 92999 59334
rect 93117 59394 93183 59397
rect 94313 59394 94379 59397
rect 93117 59392 94379 59394
rect 93117 59336 93122 59392
rect 93178 59336 94318 59392
rect 94374 59336 94379 59392
rect 93117 59334 94379 59336
rect 93117 59331 93183 59334
rect 94313 59331 94379 59334
rect 94497 59394 94563 59397
rect 97276 59394 97336 59606
rect 97809 59603 97875 59606
rect 97625 59530 97691 59533
rect 98453 59530 98519 59533
rect 97625 59528 98519 59530
rect 97625 59472 97630 59528
rect 97686 59472 98458 59528
rect 98514 59472 98519 59528
rect 97625 59470 98519 59472
rect 97625 59467 97691 59470
rect 98453 59467 98519 59470
rect 94497 59392 97336 59394
rect 94497 59336 94502 59392
rect 94558 59336 97336 59392
rect 94497 59334 97336 59336
rect 99281 59394 99347 59397
rect 101416 59394 101476 60044
rect 102428 59530 102488 60044
rect 99281 59392 101476 59394
rect 99281 59336 99286 59392
rect 99342 59336 101476 59392
rect 99281 59334 101476 59336
rect 101630 59470 102488 59530
rect 102593 59530 102659 59533
rect 103532 59530 103592 60044
rect 102593 59528 103592 59530
rect 102593 59472 102598 59528
rect 102654 59472 103592 59528
rect 102593 59470 103592 59472
rect 94497 59331 94563 59334
rect 99281 59331 99347 59334
rect 85481 59256 87154 59258
rect 85481 59200 85486 59256
rect 85542 59200 87154 59256
rect 85481 59198 87154 59200
rect 100661 59258 100727 59261
rect 101630 59258 101690 59470
rect 102593 59467 102659 59470
rect 102225 59394 102291 59397
rect 103421 59394 103487 59397
rect 104544 59394 104604 60044
rect 104801 59802 104867 59805
rect 105556 59802 105616 60044
rect 104801 59800 105616 59802
rect 104801 59744 104806 59800
rect 104862 59744 105616 59800
rect 104801 59742 105616 59744
rect 104801 59739 104867 59742
rect 104709 59666 104775 59669
rect 106568 59666 106628 60044
rect 104709 59664 106628 59666
rect 104709 59608 104714 59664
rect 104770 59608 106628 59664
rect 104709 59606 106628 59608
rect 104709 59603 104775 59606
rect 105721 59530 105787 59533
rect 107672 59530 107732 60044
rect 108684 59938 108744 60044
rect 105721 59528 107732 59530
rect 105721 59472 105726 59528
rect 105782 59472 107732 59528
rect 105721 59470 107732 59472
rect 108070 59878 108744 59938
rect 105721 59467 105787 59470
rect 104801 59394 104867 59397
rect 102225 59392 103346 59394
rect 102225 59336 102230 59392
rect 102286 59336 103346 59392
rect 102225 59334 103346 59336
rect 102225 59331 102291 59334
rect 100661 59256 101690 59258
rect 100661 59200 100666 59256
rect 100722 59200 101690 59256
rect 100661 59198 101690 59200
rect 103286 59258 103346 59334
rect 103421 59392 104604 59394
rect 103421 59336 103426 59392
rect 103482 59336 104604 59392
rect 103421 59334 104604 59336
rect 104758 59392 104867 59394
rect 104758 59336 104806 59392
rect 104862 59336 104867 59392
rect 103421 59331 103487 59334
rect 104758 59331 104867 59336
rect 105537 59394 105603 59397
rect 106917 59394 106983 59397
rect 107929 59394 107995 59397
rect 105537 59392 106842 59394
rect 105537 59336 105542 59392
rect 105598 59336 106842 59392
rect 105537 59334 106842 59336
rect 105537 59331 105603 59334
rect 104758 59258 104818 59331
rect 103286 59198 104818 59258
rect 106782 59258 106842 59334
rect 106917 59392 107995 59394
rect 106917 59336 106922 59392
rect 106978 59336 107934 59392
rect 107990 59336 107995 59392
rect 106917 59334 107995 59336
rect 106917 59331 106983 59334
rect 107929 59331 107995 59334
rect 108070 59258 108130 59878
rect 108205 59802 108271 59805
rect 109696 59802 109756 60044
rect 108205 59800 109756 59802
rect 108205 59744 108210 59800
rect 108266 59744 109756 59800
rect 108205 59742 109756 59744
rect 108205 59739 108271 59742
rect 108297 59666 108363 59669
rect 110708 59666 110768 60044
rect 108297 59664 110768 59666
rect 108297 59608 108302 59664
rect 108358 59608 110768 59664
rect 108297 59606 110768 59608
rect 110873 59666 110939 59669
rect 111812 59666 111872 60044
rect 112824 59938 112884 60044
rect 110873 59664 111872 59666
rect 110873 59608 110878 59664
rect 110934 59608 111872 59664
rect 110873 59606 111872 59608
rect 112302 59878 112884 59938
rect 108297 59603 108363 59606
rect 110873 59603 110939 59606
rect 109677 59530 109743 59533
rect 112302 59530 112362 59878
rect 112529 59802 112595 59805
rect 113836 59802 113896 60044
rect 112529 59800 113896 59802
rect 112529 59744 112534 59800
rect 112590 59744 113896 59800
rect 112529 59742 113896 59744
rect 112529 59739 112595 59742
rect 112437 59666 112503 59669
rect 114848 59666 114908 60044
rect 112437 59664 114908 59666
rect 112437 59608 112442 59664
rect 112498 59608 114908 59664
rect 112437 59606 114908 59608
rect 112437 59603 112503 59606
rect 109677 59528 112362 59530
rect 109677 59472 109682 59528
rect 109738 59472 112362 59528
rect 109677 59470 112362 59472
rect 113817 59530 113883 59533
rect 115952 59530 116012 60044
rect 113817 59528 116012 59530
rect 113817 59472 113822 59528
rect 113878 59472 116012 59528
rect 113817 59470 116012 59472
rect 116117 59530 116183 59533
rect 116964 59530 117024 60044
rect 116117 59528 117024 59530
rect 116117 59472 116122 59528
rect 116178 59472 117024 59528
rect 116117 59470 117024 59472
rect 109677 59467 109743 59470
rect 113817 59467 113883 59470
rect 116117 59467 116183 59470
rect 111057 59394 111123 59397
rect 112529 59394 112595 59397
rect 111057 59392 112595 59394
rect 111057 59336 111062 59392
rect 111118 59336 112534 59392
rect 112590 59336 112595 59392
rect 111057 59334 112595 59336
rect 111057 59331 111123 59334
rect 112529 59331 112595 59334
rect 115197 59394 115263 59397
rect 117976 59394 118036 60044
rect 118141 59666 118207 59669
rect 118988 59666 119048 60044
rect 118141 59664 119048 59666
rect 118141 59608 118146 59664
rect 118202 59608 119048 59664
rect 118141 59606 119048 59608
rect 118141 59603 118207 59606
rect 118141 59530 118207 59533
rect 120092 59530 120152 60044
rect 120257 59802 120323 59805
rect 121104 59802 121164 60044
rect 120257 59800 121164 59802
rect 120257 59744 120262 59800
rect 120318 59744 121164 59800
rect 120257 59742 121164 59744
rect 121269 59802 121335 59805
rect 122116 59802 122176 60044
rect 121269 59800 122176 59802
rect 121269 59744 121274 59800
rect 121330 59744 122176 59800
rect 121269 59742 122176 59744
rect 120257 59739 120323 59742
rect 121269 59739 121335 59742
rect 120901 59666 120967 59669
rect 120901 59664 122298 59666
rect 120901 59608 120906 59664
rect 120962 59608 122298 59664
rect 120901 59606 122298 59608
rect 120901 59603 120967 59606
rect 121269 59530 121335 59533
rect 118141 59528 120152 59530
rect 118141 59472 118146 59528
rect 118202 59472 120152 59528
rect 118141 59470 120152 59472
rect 120214 59528 121335 59530
rect 120214 59472 121274 59528
rect 121330 59472 121335 59528
rect 120214 59470 121335 59472
rect 122238 59530 122298 59606
rect 123128 59530 123188 60044
rect 122238 59470 123188 59530
rect 118141 59467 118207 59470
rect 115197 59392 118036 59394
rect 115197 59336 115202 59392
rect 115258 59336 118036 59392
rect 115197 59334 118036 59336
rect 119337 59394 119403 59397
rect 120214 59394 120274 59470
rect 121269 59467 121335 59470
rect 119337 59392 120274 59394
rect 119337 59336 119342 59392
rect 119398 59336 120274 59392
rect 119337 59334 120274 59336
rect 120717 59394 120783 59397
rect 122097 59394 122163 59397
rect 122833 59394 122899 59397
rect 124140 59394 124200 60044
rect 125244 59394 125304 60044
rect 125409 59666 125475 59669
rect 126256 59666 126316 60044
rect 125409 59664 126316 59666
rect 125409 59608 125414 59664
rect 125470 59608 126316 59664
rect 125409 59606 126316 59608
rect 125409 59603 125475 59606
rect 125409 59530 125475 59533
rect 127268 59530 127328 60044
rect 128077 59530 128143 59533
rect 125409 59528 127328 59530
rect 125409 59472 125414 59528
rect 125470 59472 127328 59528
rect 125409 59470 127328 59472
rect 127390 59528 128143 59530
rect 127390 59472 128082 59528
rect 128138 59472 128143 59528
rect 127390 59470 128143 59472
rect 125409 59467 125475 59470
rect 120717 59392 121930 59394
rect 120717 59336 120722 59392
rect 120778 59336 121930 59392
rect 120717 59334 121930 59336
rect 115197 59331 115263 59334
rect 119337 59331 119403 59334
rect 120717 59331 120783 59334
rect 106782 59198 108130 59258
rect 121870 59258 121930 59334
rect 122097 59392 122899 59394
rect 122097 59336 122102 59392
rect 122158 59336 122838 59392
rect 122894 59336 122899 59392
rect 122097 59334 122899 59336
rect 122097 59331 122163 59334
rect 122833 59331 122899 59334
rect 122974 59334 124200 59394
rect 124262 59334 125304 59394
rect 126237 59394 126303 59397
rect 127390 59394 127450 59470
rect 128077 59467 128143 59470
rect 128280 59394 128340 60044
rect 128445 59802 128511 59805
rect 129384 59802 129444 60044
rect 128445 59800 129444 59802
rect 128445 59744 128450 59800
rect 128506 59744 129444 59800
rect 128445 59742 129444 59744
rect 128445 59739 128511 59742
rect 130396 59666 130456 60044
rect 126237 59392 127450 59394
rect 126237 59336 126242 59392
rect 126298 59336 127450 59392
rect 126237 59334 127450 59336
rect 127574 59334 128340 59394
rect 128494 59606 130456 59666
rect 122974 59258 123034 59334
rect 121870 59198 123034 59258
rect 123109 59258 123175 59261
rect 124262 59258 124322 59334
rect 126237 59331 126303 59334
rect 123109 59256 124322 59258
rect 123109 59200 123114 59256
rect 123170 59200 124322 59256
rect 123109 59198 124322 59200
rect 124857 59258 124923 59261
rect 127574 59258 127634 59334
rect 124857 59256 127634 59258
rect 124857 59200 124862 59256
rect 124918 59200 127634 59256
rect 124857 59198 127634 59200
rect 127709 59258 127775 59261
rect 128494 59258 128554 59606
rect 129181 59530 129247 59533
rect 131408 59530 131468 60044
rect 132420 59938 132480 60044
rect 131622 59878 132480 59938
rect 131622 59805 131682 59878
rect 131573 59800 131682 59805
rect 133524 59802 133584 60044
rect 131573 59744 131578 59800
rect 131634 59744 131682 59800
rect 131573 59742 131682 59744
rect 132450 59742 133584 59802
rect 131573 59739 131639 59742
rect 129181 59528 131468 59530
rect 129181 59472 129186 59528
rect 129242 59472 131468 59528
rect 129181 59470 131468 59472
rect 129181 59467 129247 59470
rect 130377 59394 130443 59397
rect 132450 59394 132510 59742
rect 132585 59666 132651 59669
rect 134536 59666 134596 60044
rect 132585 59664 134596 59666
rect 132585 59608 132590 59664
rect 132646 59608 134596 59664
rect 132585 59606 134596 59608
rect 132585 59603 132651 59606
rect 133137 59530 133203 59533
rect 135548 59530 135608 60044
rect 133137 59528 135608 59530
rect 133137 59472 133142 59528
rect 133198 59472 135608 59528
rect 133137 59470 135608 59472
rect 133137 59467 133203 59470
rect 130377 59392 132510 59394
rect 130377 59336 130382 59392
rect 130438 59336 132510 59392
rect 130377 59334 132510 59336
rect 133321 59394 133387 59397
rect 136560 59394 136620 60044
rect 137664 59666 137724 60044
rect 137829 59802 137895 59805
rect 138676 59802 138736 60044
rect 139688 59938 139748 60044
rect 138982 59878 139748 59938
rect 138982 59805 139042 59878
rect 137829 59800 138736 59802
rect 137829 59744 137834 59800
rect 137890 59744 138736 59800
rect 137829 59742 138736 59744
rect 138933 59800 139042 59805
rect 140700 59802 140760 60044
rect 138933 59744 138938 59800
rect 138994 59744 139042 59800
rect 138933 59742 139042 59744
rect 139718 59742 140760 59802
rect 137829 59739 137895 59742
rect 138933 59739 138999 59742
rect 133321 59392 136620 59394
rect 133321 59336 133326 59392
rect 133382 59336 136620 59392
rect 133321 59334 136620 59336
rect 136774 59606 137724 59666
rect 137829 59666 137895 59669
rect 139718 59666 139778 59742
rect 141804 59666 141864 60044
rect 141969 59802 142035 59805
rect 142816 59802 142876 60044
rect 141969 59800 142876 59802
rect 141969 59744 141974 59800
rect 142030 59744 142876 59800
rect 141969 59742 142876 59744
rect 141969 59739 142035 59742
rect 137829 59664 139778 59666
rect 137829 59608 137834 59664
rect 137890 59608 139778 59664
rect 137829 59606 139778 59608
rect 139902 59606 141864 59666
rect 130377 59331 130443 59334
rect 133321 59331 133387 59334
rect 127709 59256 128554 59258
rect 127709 59200 127714 59256
rect 127770 59200 128554 59256
rect 127709 59198 128554 59200
rect 134517 59258 134583 59261
rect 136774 59258 136834 59606
rect 137829 59603 137895 59606
rect 137461 59530 137527 59533
rect 138933 59530 138999 59533
rect 137461 59528 138999 59530
rect 137461 59472 137466 59528
rect 137522 59472 138938 59528
rect 138994 59472 138999 59528
rect 137461 59470 138999 59472
rect 137461 59467 137527 59470
rect 138933 59467 138999 59470
rect 137277 59394 137343 59397
rect 137829 59394 137895 59397
rect 137277 59392 137895 59394
rect 137277 59336 137282 59392
rect 137338 59336 137834 59392
rect 137890 59336 137895 59392
rect 137277 59334 137895 59336
rect 137277 59331 137343 59334
rect 137829 59331 137895 59334
rect 138657 59394 138723 59397
rect 139902 59394 139962 59606
rect 141417 59530 141483 59533
rect 143828 59530 143888 60044
rect 141417 59528 143888 59530
rect 141417 59472 141422 59528
rect 141478 59472 143888 59528
rect 141417 59470 143888 59472
rect 141417 59467 141483 59470
rect 138657 59392 139962 59394
rect 138657 59336 138662 59392
rect 138718 59336 139962 59392
rect 138657 59334 139962 59336
rect 141601 59394 141667 59397
rect 144840 59394 144900 60044
rect 145005 59802 145071 59805
rect 145944 59802 146004 60044
rect 145005 59800 146004 59802
rect 145005 59744 145010 59800
rect 145066 59744 146004 59800
rect 145005 59742 146004 59744
rect 145005 59739 145071 59742
rect 146956 59666 147016 60044
rect 141601 59392 144900 59394
rect 141601 59336 141606 59392
rect 141662 59336 144900 59392
rect 141601 59334 144900 59336
rect 145054 59606 147016 59666
rect 138657 59331 138723 59334
rect 141601 59331 141667 59334
rect 134517 59256 136834 59258
rect 134517 59200 134522 59256
rect 134578 59200 136834 59256
rect 134517 59198 136834 59200
rect 144177 59258 144243 59261
rect 145054 59258 145114 59606
rect 145557 59530 145623 59533
rect 147968 59530 148028 60044
rect 148980 59938 149040 60044
rect 148182 59878 149040 59938
rect 148182 59805 148242 59878
rect 148133 59800 148242 59805
rect 150084 59802 150144 60044
rect 148133 59744 148138 59800
rect 148194 59744 148242 59800
rect 148133 59742 148242 59744
rect 148550 59742 150144 59802
rect 150249 59802 150315 59805
rect 151096 59802 151156 60044
rect 150249 59800 151156 59802
rect 150249 59744 150254 59800
rect 150310 59744 151156 59800
rect 150249 59742 151156 59744
rect 148133 59739 148199 59742
rect 148550 59666 148610 59742
rect 150249 59739 150315 59742
rect 145557 59528 148028 59530
rect 145557 59472 145562 59528
rect 145618 59472 148028 59528
rect 145557 59470 148028 59472
rect 148182 59606 148610 59666
rect 149697 59666 149763 59669
rect 149697 59664 151830 59666
rect 149697 59608 149702 59664
rect 149758 59608 151830 59664
rect 149697 59606 151830 59608
rect 145557 59467 145623 59470
rect 146937 59394 147003 59397
rect 148182 59394 148242 59606
rect 149697 59603 149763 59606
rect 148317 59530 148383 59533
rect 150249 59530 150315 59533
rect 148317 59528 150315 59530
rect 148317 59472 148322 59528
rect 148378 59472 150254 59528
rect 150310 59472 150315 59528
rect 148317 59470 150315 59472
rect 151770 59530 151830 59606
rect 152108 59530 152168 60044
rect 152273 59802 152339 59805
rect 153120 59802 153180 60044
rect 152273 59800 153180 59802
rect 152273 59744 152278 59800
rect 152334 59744 153180 59800
rect 152273 59742 153180 59744
rect 152273 59739 152339 59742
rect 154132 59666 154192 60044
rect 151770 59470 152168 59530
rect 152966 59606 154192 59666
rect 154297 59666 154363 59669
rect 155236 59666 155296 60044
rect 154297 59664 155296 59666
rect 154297 59608 154302 59664
rect 154358 59608 155296 59664
rect 154297 59606 155296 59608
rect 148317 59467 148383 59470
rect 150249 59467 150315 59470
rect 146937 59392 148242 59394
rect 146937 59336 146942 59392
rect 146998 59336 148242 59392
rect 146937 59334 148242 59336
rect 151077 59394 151143 59397
rect 152966 59394 153026 59606
rect 154297 59603 154363 59606
rect 154021 59530 154087 59533
rect 156248 59530 156308 60044
rect 156597 59802 156663 59805
rect 157260 59802 157320 60044
rect 158272 59938 158332 60044
rect 159376 59938 159436 60044
rect 160388 59938 160448 60044
rect 157566 59878 158332 59938
rect 158486 59878 159436 59938
rect 159590 59878 160448 59938
rect 156597 59800 157320 59802
rect 156597 59744 156602 59800
rect 156658 59744 157320 59800
rect 156597 59742 157320 59744
rect 157425 59802 157491 59805
rect 157566 59802 157626 59878
rect 157425 59800 157626 59802
rect 157425 59744 157430 59800
rect 157486 59744 157626 59800
rect 157425 59742 157626 59744
rect 156597 59739 156663 59742
rect 157425 59739 157491 59742
rect 156597 59666 156663 59669
rect 158486 59666 158546 59878
rect 159590 59805 159650 59878
rect 159541 59800 159650 59805
rect 159541 59744 159546 59800
rect 159602 59744 159650 59800
rect 159541 59742 159650 59744
rect 159541 59739 159607 59742
rect 156597 59664 158546 59666
rect 156597 59608 156602 59664
rect 156658 59608 158546 59664
rect 156597 59606 158546 59608
rect 158621 59666 158687 59669
rect 158621 59664 159834 59666
rect 158621 59608 158626 59664
rect 158682 59608 159834 59664
rect 158621 59606 159834 59608
rect 156597 59603 156663 59606
rect 158621 59603 158687 59606
rect 154021 59528 156308 59530
rect 154021 59472 154026 59528
rect 154082 59472 156308 59528
rect 154021 59470 156308 59472
rect 157977 59530 158043 59533
rect 159541 59530 159607 59533
rect 157977 59528 159607 59530
rect 157977 59472 157982 59528
rect 158038 59472 159546 59528
rect 159602 59472 159607 59528
rect 157977 59470 159607 59472
rect 159774 59530 159834 59606
rect 161400 59530 161460 60044
rect 159774 59470 161460 59530
rect 154021 59467 154087 59470
rect 157977 59467 158043 59470
rect 159541 59467 159607 59470
rect 154297 59394 154363 59397
rect 151077 59392 153026 59394
rect 151077 59336 151082 59392
rect 151138 59336 153026 59392
rect 151077 59334 153026 59336
rect 153120 59392 154363 59394
rect 153120 59336 154302 59392
rect 154358 59336 154363 59392
rect 153120 59334 154363 59336
rect 146937 59331 147003 59334
rect 151077 59331 151143 59334
rect 144177 59256 145114 59258
rect 144177 59200 144182 59256
rect 144238 59200 145114 59256
rect 144177 59198 145114 59200
rect 152457 59258 152523 59261
rect 153120 59258 153180 59334
rect 154297 59331 154363 59334
rect 155217 59394 155283 59397
rect 157425 59394 157491 59397
rect 155217 59392 157491 59394
rect 155217 59336 155222 59392
rect 155278 59336 157430 59392
rect 157486 59336 157491 59392
rect 155217 59334 157491 59336
rect 155217 59331 155283 59334
rect 157425 59331 157491 59334
rect 159357 59394 159423 59397
rect 162412 59394 162472 60044
rect 162577 59802 162643 59805
rect 163516 59802 163576 60044
rect 162577 59800 163576 59802
rect 162577 59744 162582 59800
rect 162638 59744 163576 59800
rect 162577 59742 163576 59744
rect 162577 59739 162643 59742
rect 162577 59530 162643 59533
rect 164528 59530 164588 60044
rect 165540 59802 165600 60044
rect 162577 59528 164588 59530
rect 162577 59472 162582 59528
rect 162638 59472 164588 59528
rect 162577 59470 164588 59472
rect 164742 59742 165600 59802
rect 165705 59802 165771 59805
rect 166552 59802 166612 60044
rect 165705 59800 166612 59802
rect 165705 59744 165710 59800
rect 165766 59744 166612 59800
rect 165705 59742 166612 59744
rect 162577 59467 162643 59470
rect 159357 59392 162472 59394
rect 159357 59336 159362 59392
rect 159418 59336 162472 59392
rect 159357 59334 162472 59336
rect 162577 59394 162643 59397
rect 164742 59394 164802 59742
rect 165705 59739 165771 59742
rect 164877 59666 164943 59669
rect 167656 59666 167716 60044
rect 164877 59664 167716 59666
rect 164877 59608 164882 59664
rect 164938 59608 167716 59664
rect 164877 59606 167716 59608
rect 164877 59603 164943 59606
rect 166809 59530 166875 59533
rect 168668 59530 168728 60044
rect 166809 59528 168728 59530
rect 166809 59472 166814 59528
rect 166870 59472 168728 59528
rect 166809 59470 168728 59472
rect 166809 59467 166875 59470
rect 165705 59394 165771 59397
rect 162577 59392 164802 59394
rect 162577 59336 162582 59392
rect 162638 59336 164802 59392
rect 162577 59334 164802 59336
rect 164926 59392 165771 59394
rect 164926 59336 165710 59392
rect 165766 59336 165771 59392
rect 164926 59334 165771 59336
rect 159357 59331 159423 59334
rect 162577 59331 162643 59334
rect 152457 59256 153180 59258
rect 152457 59200 152462 59256
rect 152518 59200 153180 59256
rect 152457 59198 153180 59200
rect 164141 59258 164207 59261
rect 164926 59258 164986 59334
rect 165705 59331 165771 59334
rect 166625 59394 166691 59397
rect 169680 59394 169740 60044
rect 170692 59394 170752 60044
rect 170949 59802 171015 59805
rect 172808 59802 172868 60044
rect 170949 59800 172868 59802
rect 170949 59744 170954 59800
rect 171010 59744 172868 59800
rect 170949 59742 172868 59744
rect 170949 59739 171015 59742
rect 170857 59666 170923 59669
rect 173820 59666 173880 60044
rect 170857 59664 173880 59666
rect 170857 59608 170862 59664
rect 170918 59608 173880 59664
rect 170857 59606 173880 59608
rect 170857 59603 170923 59606
rect 166625 59392 169740 59394
rect 166625 59336 166630 59392
rect 166686 59336 169740 59392
rect 166625 59334 169740 59336
rect 169894 59334 170752 59394
rect 172421 59394 172487 59397
rect 174832 59394 174892 60044
rect 175936 59394 175996 60044
rect 176948 59530 177008 60044
rect 172421 59392 174892 59394
rect 172421 59336 172426 59392
rect 172482 59336 174892 59392
rect 172421 59334 174892 59336
rect 175046 59334 175996 59394
rect 176150 59470 177008 59530
rect 177113 59530 177179 59533
rect 177960 59530 178020 60044
rect 178217 59802 178283 59805
rect 178972 59802 179032 60044
rect 178217 59800 179032 59802
rect 178217 59744 178222 59800
rect 178278 59744 179032 59800
rect 178217 59742 179032 59744
rect 178217 59739 178283 59742
rect 178125 59666 178191 59669
rect 180076 59666 180136 60044
rect 178125 59664 180136 59666
rect 178125 59608 178130 59664
rect 178186 59608 180136 59664
rect 178125 59606 180136 59608
rect 178125 59603 178191 59606
rect 177113 59528 178020 59530
rect 177113 59472 177118 59528
rect 177174 59472 178020 59528
rect 177113 59470 178020 59472
rect 179137 59530 179203 59533
rect 181088 59530 181148 60044
rect 182100 59938 182160 60044
rect 181302 59878 182160 59938
rect 181302 59805 181362 59878
rect 181253 59800 181362 59805
rect 183112 59802 183172 60044
rect 181253 59744 181258 59800
rect 181314 59744 181362 59800
rect 181253 59742 181362 59744
rect 181670 59742 183172 59802
rect 181253 59739 181319 59742
rect 181670 59530 181730 59742
rect 182081 59666 182147 59669
rect 184124 59666 184184 60044
rect 182081 59664 184184 59666
rect 182081 59608 182086 59664
rect 182142 59608 184184 59664
rect 182081 59606 184184 59608
rect 182081 59603 182147 59606
rect 179137 59528 181148 59530
rect 179137 59472 179142 59528
rect 179198 59472 181148 59528
rect 179137 59470 181148 59472
rect 181302 59470 181730 59530
rect 183185 59530 183251 59533
rect 185228 59530 185288 60044
rect 186240 59666 186300 60044
rect 183185 59528 185288 59530
rect 183185 59472 183190 59528
rect 183246 59472 185288 59528
rect 183185 59470 185288 59472
rect 185350 59606 186300 59666
rect 166625 59331 166691 59334
rect 164141 59256 164986 59258
rect 164141 59200 164146 59256
rect 164202 59200 164986 59256
rect 164141 59198 164986 59200
rect 168281 59258 168347 59261
rect 169894 59258 169954 59334
rect 172421 59331 172487 59334
rect 168281 59256 169954 59258
rect 168281 59200 168286 59256
rect 168342 59200 169954 59256
rect 168281 59198 169954 59200
rect 173801 59258 173867 59261
rect 175046 59258 175106 59334
rect 173801 59256 175106 59258
rect 173801 59200 173806 59256
rect 173862 59200 175106 59256
rect 173801 59198 175106 59200
rect 85481 59195 85547 59198
rect 100661 59195 100727 59198
rect 123109 59195 123175 59198
rect 124857 59195 124923 59198
rect 127709 59195 127775 59198
rect 134517 59195 134583 59198
rect 144177 59195 144243 59198
rect 152457 59195 152523 59198
rect 164141 59195 164207 59198
rect 168281 59195 168347 59198
rect 173801 59195 173867 59198
rect 174905 59122 174971 59125
rect 176150 59122 176210 59470
rect 177113 59467 177179 59470
rect 179137 59467 179203 59470
rect 176561 59394 176627 59397
rect 178217 59394 178283 59397
rect 176561 59392 178283 59394
rect 176561 59336 176566 59392
rect 176622 59336 178222 59392
rect 178278 59336 178283 59392
rect 176561 59334 178283 59336
rect 176561 59331 176627 59334
rect 178217 59331 178283 59334
rect 180701 59394 180767 59397
rect 181302 59394 181362 59470
rect 183185 59467 183251 59470
rect 180701 59392 181362 59394
rect 180701 59336 180706 59392
rect 180762 59336 181362 59392
rect 180701 59334 181362 59336
rect 183461 59394 183527 59397
rect 185350 59394 185410 59606
rect 187252 59530 187312 60044
rect 188264 59666 188324 60044
rect 188981 59666 189047 59669
rect 188264 59664 189047 59666
rect 188264 59608 188986 59664
rect 189042 59608 189047 59664
rect 188264 59606 189047 59608
rect 188981 59603 189047 59606
rect 186270 59470 187312 59530
rect 187417 59530 187483 59533
rect 189368 59530 189428 60044
rect 187417 59528 189428 59530
rect 187417 59472 187422 59528
rect 187478 59472 189428 59528
rect 187417 59470 189428 59472
rect 186270 59394 186330 59470
rect 187417 59467 187483 59470
rect 183461 59392 185410 59394
rect 183461 59336 183466 59392
rect 183522 59336 185410 59392
rect 183461 59334 185410 59336
rect 185534 59334 186330 59394
rect 187509 59394 187575 59397
rect 190380 59394 190440 60044
rect 190545 59802 190611 59805
rect 191392 59802 191452 60044
rect 190545 59800 191452 59802
rect 190545 59744 190550 59800
rect 190606 59744 191452 59800
rect 190545 59742 191452 59744
rect 190545 59739 190611 59742
rect 190545 59666 190611 59669
rect 192404 59666 192464 60044
rect 190545 59664 192464 59666
rect 190545 59608 190550 59664
rect 190606 59608 192464 59664
rect 190545 59606 192464 59608
rect 190545 59603 190611 59606
rect 191465 59530 191531 59533
rect 193508 59530 193568 60044
rect 191465 59528 193568 59530
rect 191465 59472 191470 59528
rect 191526 59472 193568 59528
rect 191465 59470 193568 59472
rect 193673 59530 193739 59533
rect 194520 59530 194580 60044
rect 195532 59938 195592 60044
rect 193673 59528 194580 59530
rect 193673 59472 193678 59528
rect 193734 59472 194580 59528
rect 193673 59470 194580 59472
rect 194734 59878 195592 59938
rect 191465 59467 191531 59470
rect 193673 59467 193739 59470
rect 187509 59392 190440 59394
rect 187509 59336 187514 59392
rect 187570 59336 190440 59392
rect 187509 59334 190440 59336
rect 193121 59394 193187 59397
rect 194734 59394 194794 59878
rect 195789 59802 195855 59805
rect 196544 59802 196604 60044
rect 195789 59800 196604 59802
rect 195789 59744 195794 59800
rect 195850 59744 196604 59800
rect 195789 59742 196604 59744
rect 196801 59802 196867 59805
rect 197648 59802 197708 60044
rect 196801 59800 197708 59802
rect 196801 59744 196806 59800
rect 196862 59744 197708 59800
rect 196801 59742 197708 59744
rect 195789 59739 195855 59742
rect 196801 59739 196867 59742
rect 195789 59666 195855 59669
rect 198660 59666 198720 60044
rect 198825 59802 198891 59805
rect 199672 59802 199732 60044
rect 200684 59938 200744 60044
rect 198825 59800 199732 59802
rect 198825 59744 198830 59800
rect 198886 59744 199732 59800
rect 198825 59742 199732 59744
rect 199886 59878 200744 59938
rect 198825 59739 198891 59742
rect 199886 59666 199946 59878
rect 195789 59664 198720 59666
rect 195789 59608 195794 59664
rect 195850 59608 198720 59664
rect 195789 59606 198720 59608
rect 199702 59606 199946 59666
rect 200021 59666 200087 59669
rect 201788 59666 201848 60044
rect 200021 59664 201848 59666
rect 200021 59608 200026 59664
rect 200082 59608 201848 59664
rect 200021 59606 201848 59608
rect 195789 59603 195855 59606
rect 195697 59530 195763 59533
rect 196801 59530 196867 59533
rect 195697 59528 196867 59530
rect 195697 59472 195702 59528
rect 195758 59472 196806 59528
rect 196862 59472 196867 59528
rect 195697 59470 196867 59472
rect 195697 59467 195763 59470
rect 196801 59467 196867 59470
rect 198641 59530 198707 59533
rect 199702 59530 199762 59606
rect 200021 59603 200087 59606
rect 198641 59528 199762 59530
rect 198641 59472 198646 59528
rect 198702 59472 199762 59528
rect 198641 59470 199762 59472
rect 199837 59530 199903 59533
rect 202800 59530 202860 60044
rect 199837 59528 202860 59530
rect 199837 59472 199842 59528
rect 199898 59472 202860 59528
rect 199837 59470 202860 59472
rect 198641 59467 198707 59470
rect 199837 59467 199903 59470
rect 193121 59392 194794 59394
rect 193121 59336 193126 59392
rect 193182 59336 194794 59392
rect 193121 59334 194794 59336
rect 197261 59394 197327 59397
rect 198825 59394 198891 59397
rect 197261 59392 198891 59394
rect 197261 59336 197266 59392
rect 197322 59336 198830 59392
rect 198886 59336 198891 59392
rect 197261 59334 198891 59336
rect 180701 59331 180767 59334
rect 183461 59331 183527 59334
rect 184841 59258 184907 59261
rect 185534 59258 185594 59334
rect 187509 59331 187575 59334
rect 193121 59331 193187 59334
rect 197261 59331 197327 59334
rect 198825 59331 198891 59334
rect 201401 59394 201467 59397
rect 203812 59394 203872 60044
rect 204824 59394 204884 60044
rect 205928 59530 205988 60044
rect 201401 59392 203872 59394
rect 201401 59336 201406 59392
rect 201462 59336 203872 59392
rect 201401 59334 203872 59336
rect 203934 59334 204884 59394
rect 205038 59470 205988 59530
rect 206093 59530 206159 59533
rect 206940 59530 207000 60044
rect 206093 59528 207000 59530
rect 206093 59472 206098 59528
rect 206154 59472 207000 59528
rect 206093 59470 207000 59472
rect 201401 59331 201467 59334
rect 184841 59256 185594 59258
rect 184841 59200 184846 59256
rect 184902 59200 185594 59256
rect 184841 59198 185594 59200
rect 202781 59258 202847 59261
rect 203934 59258 203994 59334
rect 202781 59256 203994 59258
rect 202781 59200 202786 59256
rect 202842 59200 203994 59256
rect 202781 59198 203994 59200
rect 204069 59258 204135 59261
rect 205038 59258 205098 59470
rect 206093 59467 206159 59470
rect 205541 59394 205607 59397
rect 207952 59394 208012 60044
rect 208964 59938 209024 60044
rect 208166 59878 209024 59938
rect 210068 59938 210128 60044
rect 210068 59878 210250 59938
rect 208166 59805 208226 59878
rect 208117 59800 208226 59805
rect 209957 59802 210023 59805
rect 208117 59744 208122 59800
rect 208178 59744 208226 59800
rect 208117 59742 208226 59744
rect 209086 59800 210023 59802
rect 209086 59744 209962 59800
rect 210018 59744 210023 59800
rect 209086 59742 210023 59744
rect 208117 59739 208183 59742
rect 208209 59666 208275 59669
rect 209086 59666 209146 59742
rect 209957 59739 210023 59742
rect 210190 59666 210250 59878
rect 210325 59802 210391 59805
rect 211080 59802 211140 60044
rect 210325 59800 211140 59802
rect 210325 59744 210330 59800
rect 210386 59744 211140 59800
rect 210325 59742 211140 59744
rect 211245 59802 211311 59805
rect 212092 59802 212152 60044
rect 211245 59800 212152 59802
rect 211245 59744 211250 59800
rect 211306 59744 212152 59800
rect 211245 59742 212152 59744
rect 210325 59739 210391 59742
rect 211245 59739 211311 59742
rect 208209 59664 209146 59666
rect 208209 59608 208214 59664
rect 208270 59608 209146 59664
rect 208209 59606 209146 59608
rect 210068 59606 210250 59666
rect 211061 59666 211127 59669
rect 213104 59666 213164 60044
rect 211061 59664 213164 59666
rect 211061 59608 211066 59664
rect 211122 59608 213164 59664
rect 211061 59606 213164 59608
rect 208209 59603 208275 59606
rect 208117 59530 208183 59533
rect 210068 59530 210128 59606
rect 211061 59603 211127 59606
rect 208117 59528 210128 59530
rect 208117 59472 208122 59528
rect 208178 59472 210128 59528
rect 208117 59470 210128 59472
rect 212257 59530 212323 59533
rect 214116 59530 214176 60044
rect 215220 59666 215280 60044
rect 212257 59528 214176 59530
rect 212257 59472 212262 59528
rect 212318 59472 214176 59528
rect 212257 59470 214176 59472
rect 214238 59606 215280 59666
rect 208117 59467 208183 59470
rect 212257 59467 212323 59470
rect 205541 59392 208012 59394
rect 205541 59336 205546 59392
rect 205602 59336 208012 59392
rect 205541 59334 208012 59336
rect 209681 59394 209747 59397
rect 211245 59394 211311 59397
rect 209681 59392 211311 59394
rect 209681 59336 209686 59392
rect 209742 59336 211250 59392
rect 211306 59336 211311 59392
rect 209681 59334 211311 59336
rect 205541 59331 205607 59334
rect 209681 59331 209747 59334
rect 211245 59331 211311 59334
rect 212349 59394 212415 59397
rect 214238 59394 214298 59606
rect 216232 59530 216292 60044
rect 217244 59666 217304 60044
rect 217961 59666 218027 59669
rect 217244 59664 218027 59666
rect 217244 59608 217966 59664
rect 218022 59608 218027 59664
rect 217244 59606 218027 59608
rect 217961 59603 218027 59606
rect 215250 59470 216292 59530
rect 216397 59530 216463 59533
rect 218256 59530 218316 60044
rect 219360 59666 219420 60044
rect 216397 59528 218316 59530
rect 216397 59472 216402 59528
rect 216458 59472 218316 59528
rect 216397 59470 218316 59472
rect 218470 59606 219420 59666
rect 219893 59666 219959 59669
rect 220372 59666 220432 60044
rect 219893 59664 220432 59666
rect 219893 59608 219898 59664
rect 219954 59608 220432 59664
rect 219893 59606 220432 59608
rect 215250 59394 215310 59470
rect 216397 59467 216463 59470
rect 212349 59392 214298 59394
rect 212349 59336 212354 59392
rect 212410 59336 214298 59392
rect 212349 59334 214298 59336
rect 214422 59334 215310 59394
rect 216489 59394 216555 59397
rect 218470 59394 218530 59606
rect 219893 59603 219959 59606
rect 219341 59530 219407 59533
rect 221384 59530 221444 60044
rect 219341 59528 221444 59530
rect 219341 59472 219346 59528
rect 219402 59472 221444 59528
rect 219341 59470 221444 59472
rect 219341 59467 219407 59470
rect 219893 59394 219959 59397
rect 216489 59392 218530 59394
rect 216489 59336 216494 59392
rect 216550 59336 218530 59392
rect 216489 59334 218530 59336
rect 218654 59392 219959 59394
rect 218654 59336 219898 59392
rect 219954 59336 219959 59392
rect 218654 59334 219959 59336
rect 212349 59331 212415 59334
rect 204069 59256 205098 59258
rect 204069 59200 204074 59256
rect 204130 59200 205098 59256
rect 204069 59198 205098 59200
rect 213821 59258 213887 59261
rect 214422 59258 214482 59334
rect 216489 59331 216555 59334
rect 213821 59256 214482 59258
rect 213821 59200 213826 59256
rect 213882 59200 214482 59256
rect 213821 59198 214482 59200
rect 217869 59258 217935 59261
rect 218654 59258 218714 59334
rect 219893 59331 219959 59334
rect 220629 59394 220695 59397
rect 222396 59394 222456 60044
rect 222561 59802 222627 59805
rect 223500 59802 223560 60044
rect 222561 59800 223560 59802
rect 222561 59744 222566 59800
rect 222622 59744 223560 59800
rect 222561 59742 223560 59744
rect 223665 59802 223731 59805
rect 224512 59802 224572 60044
rect 223665 59800 224572 59802
rect 223665 59744 223670 59800
rect 223726 59744 224572 59800
rect 223665 59742 224572 59744
rect 222561 59739 222627 59742
rect 223665 59739 223731 59742
rect 223481 59666 223547 59669
rect 225524 59666 225584 60044
rect 223481 59664 225584 59666
rect 223481 59608 223486 59664
rect 223542 59608 225584 59664
rect 223481 59606 225584 59608
rect 223481 59603 223547 59606
rect 224677 59530 224743 59533
rect 226536 59530 226596 60044
rect 224677 59528 226596 59530
rect 224677 59472 224682 59528
rect 224738 59472 226596 59528
rect 224677 59470 226596 59472
rect 226701 59530 226767 59533
rect 227640 59530 227700 60044
rect 227897 59802 227963 59805
rect 228652 59802 228712 60044
rect 227897 59800 228712 59802
rect 227897 59744 227902 59800
rect 227958 59744 228712 59800
rect 227897 59742 228712 59744
rect 227897 59739 227963 59742
rect 227805 59666 227871 59669
rect 229664 59666 229724 60044
rect 230676 59938 230736 60044
rect 227805 59664 229724 59666
rect 227805 59608 227810 59664
rect 227866 59608 229724 59664
rect 227805 59606 229724 59608
rect 229878 59878 230736 59938
rect 227805 59603 227871 59606
rect 226701 59528 227700 59530
rect 226701 59472 226706 59528
rect 226762 59472 227700 59528
rect 226701 59470 227700 59472
rect 229001 59530 229067 59533
rect 229878 59530 229938 59878
rect 231780 59802 231840 60044
rect 230798 59742 231840 59802
rect 230798 59530 230858 59742
rect 232792 59666 232852 60044
rect 229001 59528 229938 59530
rect 229001 59472 229006 59528
rect 229062 59472 229938 59528
rect 229001 59470 229938 59472
rect 230246 59470 230858 59530
rect 231166 59606 232852 59666
rect 232957 59666 233023 59669
rect 233804 59666 233864 60044
rect 232957 59664 233864 59666
rect 232957 59608 232962 59664
rect 233018 59608 233864 59664
rect 232957 59606 233864 59608
rect 224677 59467 224743 59470
rect 226701 59467 226767 59470
rect 229001 59467 229067 59470
rect 223665 59394 223731 59397
rect 220629 59392 222456 59394
rect 220629 59336 220634 59392
rect 220690 59336 222456 59392
rect 220629 59334 222456 59336
rect 222518 59392 223731 59394
rect 222518 59336 223670 59392
rect 223726 59336 223731 59392
rect 222518 59334 223731 59336
rect 220629 59331 220695 59334
rect 217869 59256 218714 59258
rect 217869 59200 217874 59256
rect 217930 59200 218714 59256
rect 217869 59198 218714 59200
rect 222101 59258 222167 59261
rect 222518 59258 222578 59334
rect 223665 59331 223731 59334
rect 226241 59394 226307 59397
rect 227897 59394 227963 59397
rect 226241 59392 227963 59394
rect 226241 59336 226246 59392
rect 226302 59336 227902 59392
rect 227958 59336 227963 59392
rect 226241 59334 227963 59336
rect 226241 59331 226307 59334
rect 227897 59331 227963 59334
rect 228817 59394 228883 59397
rect 230246 59394 230306 59470
rect 228817 59392 230306 59394
rect 228817 59336 228822 59392
rect 228878 59336 230306 59392
rect 228817 59334 230306 59336
rect 230381 59394 230447 59397
rect 231166 59394 231226 59606
rect 232957 59603 233023 59606
rect 232865 59530 232931 59533
rect 234816 59530 234876 60044
rect 232865 59528 234876 59530
rect 232865 59472 232870 59528
rect 232926 59472 234876 59528
rect 232865 59470 234876 59472
rect 234981 59530 235047 59533
rect 235920 59530 235980 60044
rect 234981 59528 235980 59530
rect 234981 59472 234986 59528
rect 235042 59472 235980 59528
rect 234981 59470 235980 59472
rect 232865 59467 232931 59470
rect 234981 59467 235047 59470
rect 230381 59392 231226 59394
rect 230381 59336 230386 59392
rect 230442 59336 231226 59392
rect 230381 59334 231226 59336
rect 231761 59394 231827 59397
rect 232957 59394 233023 59397
rect 231761 59392 233023 59394
rect 231761 59336 231766 59392
rect 231822 59336 232962 59392
rect 233018 59336 233023 59392
rect 231761 59334 233023 59336
rect 228817 59331 228883 59334
rect 230381 59331 230447 59334
rect 231761 59331 231827 59334
rect 232957 59331 233023 59334
rect 234521 59394 234587 59397
rect 236932 59394 236992 60044
rect 237944 59394 238004 60044
rect 238753 59802 238819 59805
rect 238956 59802 239016 60044
rect 238753 59800 239016 59802
rect 238753 59744 238758 59800
rect 238814 59744 239016 59800
rect 238753 59742 239016 59744
rect 238753 59739 238819 59742
rect 240060 59666 240120 60044
rect 234521 59392 236992 59394
rect 234521 59336 234526 59392
rect 234582 59336 236992 59392
rect 234521 59334 236992 59336
rect 237054 59334 238004 59394
rect 238158 59606 240120 59666
rect 234521 59331 234587 59334
rect 222101 59256 222578 59258
rect 222101 59200 222106 59256
rect 222162 59200 222578 59256
rect 222101 59198 222578 59200
rect 235901 59258 235967 59261
rect 237054 59258 237114 59334
rect 235901 59256 237114 59258
rect 235901 59200 235906 59256
rect 235962 59200 237114 59256
rect 235901 59198 237114 59200
rect 237189 59258 237255 59261
rect 238158 59258 238218 59606
rect 238753 59530 238819 59533
rect 237189 59256 238218 59258
rect 237189 59200 237194 59256
rect 237250 59200 238218 59256
rect 237189 59198 238218 59200
rect 238342 59528 238819 59530
rect 238342 59472 238758 59528
rect 238814 59472 238819 59528
rect 238342 59470 238819 59472
rect 184841 59195 184907 59198
rect 202781 59195 202847 59198
rect 204069 59195 204135 59198
rect 213821 59195 213887 59198
rect 217869 59195 217935 59198
rect 222101 59195 222167 59198
rect 235901 59195 235967 59198
rect 237189 59195 237255 59198
rect 174905 59120 176210 59122
rect 174905 59064 174910 59120
rect 174966 59064 176210 59120
rect 174905 59062 176210 59064
rect 237005 59122 237071 59125
rect 238342 59122 238402 59470
rect 238753 59467 238819 59470
rect 238661 59394 238727 59397
rect 241072 59394 241132 60044
rect 242084 59666 242144 60044
rect 242709 59666 242775 59669
rect 242084 59664 242775 59666
rect 242084 59608 242714 59664
rect 242770 59608 242775 59664
rect 242084 59606 242775 59608
rect 242709 59603 242775 59606
rect 241329 59530 241395 59533
rect 243096 59530 243156 60044
rect 244108 59938 244168 60044
rect 241329 59528 243156 59530
rect 241329 59472 241334 59528
rect 241390 59472 243156 59528
rect 241329 59470 243156 59472
rect 244046 59878 244168 59938
rect 241329 59467 241395 59470
rect 238661 59392 241132 59394
rect 238661 59336 238666 59392
rect 238722 59336 241132 59392
rect 238661 59334 241132 59336
rect 241237 59394 241303 59397
rect 244046 59394 244106 59878
rect 244273 59802 244339 59805
rect 245212 59802 245272 60044
rect 246224 59938 246284 60044
rect 247236 59938 247296 60044
rect 248248 59938 248308 60044
rect 244273 59800 245272 59802
rect 244273 59744 244278 59800
rect 244334 59744 245272 59800
rect 244273 59742 245272 59744
rect 245334 59878 246284 59938
rect 246438 59878 247296 59938
rect 247358 59878 248308 59938
rect 244273 59739 244339 59742
rect 244181 59530 244247 59533
rect 245334 59530 245394 59878
rect 245469 59666 245535 59669
rect 246438 59666 246498 59878
rect 246757 59802 246823 59805
rect 247358 59802 247418 59878
rect 246757 59800 247418 59802
rect 246757 59744 246762 59800
rect 246818 59744 247418 59800
rect 246757 59742 247418 59744
rect 248413 59802 248479 59805
rect 249352 59802 249412 60044
rect 248413 59800 249412 59802
rect 248413 59744 248418 59800
rect 248474 59744 249412 59800
rect 248413 59742 249412 59744
rect 246757 59739 246823 59742
rect 248413 59739 248479 59742
rect 250364 59666 250424 60044
rect 245469 59664 246498 59666
rect 245469 59608 245474 59664
rect 245530 59608 246498 59664
rect 245469 59606 246498 59608
rect 248462 59606 250424 59666
rect 245469 59603 245535 59606
rect 244181 59528 245394 59530
rect 244181 59472 244186 59528
rect 244242 59472 245394 59528
rect 244181 59470 245394 59472
rect 248321 59530 248387 59533
rect 248462 59530 248522 59606
rect 248321 59528 248522 59530
rect 248321 59472 248326 59528
rect 248382 59472 248522 59528
rect 248321 59470 248522 59472
rect 249425 59530 249491 59533
rect 251376 59530 251436 60044
rect 249425 59528 251436 59530
rect 249425 59472 249430 59528
rect 249486 59472 251436 59528
rect 249425 59470 251436 59472
rect 251541 59530 251607 59533
rect 252388 59530 252448 60044
rect 252645 59802 252711 59805
rect 253492 59802 253552 60044
rect 252645 59800 253552 59802
rect 252645 59744 252650 59800
rect 252706 59744 253552 59800
rect 252645 59742 253552 59744
rect 252645 59739 252711 59742
rect 252553 59666 252619 59669
rect 254504 59666 254564 60044
rect 252553 59664 254564 59666
rect 252553 59608 252558 59664
rect 252614 59608 254564 59664
rect 252553 59606 254564 59608
rect 252553 59603 252619 59606
rect 251541 59528 252448 59530
rect 251541 59472 251546 59528
rect 251602 59472 252448 59528
rect 251541 59470 252448 59472
rect 253657 59530 253723 59533
rect 255516 59530 255576 60044
rect 253657 59528 255576 59530
rect 253657 59472 253662 59528
rect 253718 59472 255576 59528
rect 253657 59470 255576 59472
rect 255681 59530 255747 59533
rect 256528 59530 256588 60044
rect 255681 59528 256588 59530
rect 255681 59472 255686 59528
rect 255742 59472 256588 59528
rect 255681 59470 256588 59472
rect 244181 59467 244247 59470
rect 248321 59467 248387 59470
rect 249425 59467 249491 59470
rect 251541 59467 251607 59470
rect 253657 59467 253723 59470
rect 255681 59467 255747 59470
rect 241237 59392 242634 59394
rect 241237 59336 241242 59392
rect 241298 59336 242634 59392
rect 241237 59334 242634 59336
rect 238661 59331 238727 59334
rect 241237 59331 241303 59334
rect 242574 59258 242634 59334
rect 243494 59334 244106 59394
rect 251081 59394 251147 59397
rect 252645 59394 252711 59397
rect 251081 59392 252711 59394
rect 251081 59336 251086 59392
rect 251142 59336 252650 59392
rect 252706 59336 252711 59392
rect 251081 59334 252711 59336
rect 243494 59258 243554 59334
rect 251081 59331 251147 59334
rect 252645 59331 252711 59334
rect 255221 59394 255287 59397
rect 257632 59394 257692 60044
rect 257797 59530 257863 59533
rect 258644 59530 258704 60044
rect 257797 59528 258704 59530
rect 257797 59472 257802 59528
rect 257858 59472 258704 59528
rect 257797 59470 258704 59472
rect 257797 59467 257863 59470
rect 255221 59392 257692 59394
rect 255221 59336 255226 59392
rect 255282 59336 257692 59392
rect 255221 59334 257692 59336
rect 257797 59394 257863 59397
rect 259656 59394 259716 60044
rect 259821 59802 259887 59805
rect 260668 59802 260728 60044
rect 259821 59800 260728 59802
rect 259821 59744 259826 59800
rect 259882 59744 260728 59800
rect 259821 59742 260728 59744
rect 259821 59739 259887 59742
rect 261772 59666 261832 60044
rect 257797 59392 259716 59394
rect 257797 59336 257802 59392
rect 257858 59336 259716 59392
rect 257797 59334 259716 59336
rect 259870 59606 261832 59666
rect 255221 59331 255287 59334
rect 257797 59331 257863 59334
rect 242574 59198 243554 59258
rect 259361 59258 259427 59261
rect 259870 59258 259930 59606
rect 260741 59530 260807 59533
rect 262784 59530 262844 60044
rect 260741 59528 262844 59530
rect 260741 59472 260746 59528
rect 260802 59472 262844 59528
rect 260741 59470 262844 59472
rect 260741 59467 260807 59470
rect 261937 59394 262003 59397
rect 263796 59394 263856 60044
rect 263961 59802 264027 59805
rect 264808 59802 264868 60044
rect 263961 59800 264868 59802
rect 263961 59744 263966 59800
rect 264022 59744 264868 59800
rect 263961 59742 264868 59744
rect 263961 59739 264027 59742
rect 265912 59666 265972 60044
rect 266169 59802 266235 59805
rect 266924 59802 266984 60044
rect 266169 59800 266984 59802
rect 266169 59744 266174 59800
rect 266230 59744 266984 59800
rect 266169 59742 266984 59744
rect 266169 59739 266235 59742
rect 261937 59392 263856 59394
rect 261937 59336 261942 59392
rect 261998 59336 263856 59392
rect 261937 59334 263856 59336
rect 263918 59606 265972 59666
rect 266077 59666 266143 59669
rect 266077 59664 267106 59666
rect 266077 59608 266082 59664
rect 266138 59608 267106 59664
rect 266077 59606 267106 59608
rect 261937 59331 262003 59334
rect 259361 59256 259930 59258
rect 259361 59200 259366 59256
rect 259422 59200 259930 59256
rect 259361 59198 259930 59200
rect 262857 59258 262923 59261
rect 263918 59258 263978 59606
rect 266077 59603 266143 59606
rect 264237 59530 264303 59533
rect 266169 59530 266235 59533
rect 264237 59528 266235 59530
rect 264237 59472 264242 59528
rect 264298 59472 266174 59528
rect 266230 59472 266235 59528
rect 264237 59470 266235 59472
rect 267046 59530 267106 59606
rect 267936 59530 267996 60044
rect 268101 59802 268167 59805
rect 268948 59802 269008 60044
rect 268101 59800 269008 59802
rect 268101 59744 268106 59800
rect 268162 59744 269008 59800
rect 268101 59742 269008 59744
rect 268101 59739 268167 59742
rect 270052 59666 270112 60044
rect 267046 59470 267996 59530
rect 268886 59606 270112 59666
rect 270217 59666 270283 59669
rect 271064 59666 271124 60044
rect 270217 59664 271124 59666
rect 270217 59608 270222 59664
rect 270278 59608 271124 59664
rect 270217 59606 271124 59608
rect 264237 59467 264303 59470
rect 266169 59467 266235 59470
rect 266997 59394 267063 59397
rect 268886 59394 268946 59606
rect 270217 59603 270283 59606
rect 269941 59530 270007 59533
rect 272076 59530 272136 60044
rect 273088 59938 273148 60044
rect 269941 59528 272136 59530
rect 269941 59472 269946 59528
rect 270002 59472 272136 59528
rect 269941 59470 272136 59472
rect 272382 59878 273148 59938
rect 269941 59467 270007 59470
rect 270217 59394 270283 59397
rect 266997 59392 268946 59394
rect 266997 59336 267002 59392
rect 267058 59336 268946 59392
rect 266997 59334 268946 59336
rect 269070 59392 270283 59394
rect 269070 59336 270222 59392
rect 270278 59336 270283 59392
rect 269070 59334 270283 59336
rect 266997 59331 267063 59334
rect 262857 59256 263978 59258
rect 262857 59200 262862 59256
rect 262918 59200 263978 59256
rect 262857 59198 263978 59200
rect 268377 59258 268443 59261
rect 269070 59258 269130 59334
rect 270217 59331 270283 59334
rect 271137 59394 271203 59397
rect 272241 59394 272307 59397
rect 271137 59392 272307 59394
rect 271137 59336 271142 59392
rect 271198 59336 272246 59392
rect 272302 59336 272307 59392
rect 271137 59334 272307 59336
rect 271137 59331 271203 59334
rect 272241 59331 272307 59334
rect 268377 59256 269130 59258
rect 268377 59200 268382 59256
rect 268438 59200 269130 59256
rect 268377 59198 269130 59200
rect 269757 59258 269823 59261
rect 272382 59258 272442 59878
rect 272517 59802 272583 59805
rect 274100 59802 274160 60044
rect 272517 59800 274160 59802
rect 272517 59744 272522 59800
rect 272578 59744 274160 59800
rect 272517 59742 274160 59744
rect 272517 59739 272583 59742
rect 272517 59666 272583 59669
rect 275204 59666 275264 60044
rect 275461 59802 275527 59805
rect 276216 59802 276276 60044
rect 275461 59800 276276 59802
rect 275461 59744 275466 59800
rect 275522 59744 276276 59800
rect 275461 59742 276276 59744
rect 276381 59802 276447 59805
rect 277228 59802 277288 60044
rect 276381 59800 277288 59802
rect 276381 59744 276386 59800
rect 276442 59744 277288 59800
rect 276381 59742 277288 59744
rect 275461 59739 275527 59742
rect 276381 59739 276447 59742
rect 272517 59664 275264 59666
rect 272517 59608 272522 59664
rect 272578 59608 275264 59664
rect 272517 59606 275264 59608
rect 275369 59666 275435 59669
rect 278240 59666 278300 60044
rect 275369 59664 278300 59666
rect 275369 59608 275374 59664
rect 275430 59608 278300 59664
rect 275369 59606 278300 59608
rect 272517 59603 272583 59606
rect 275369 59603 275435 59606
rect 274081 59530 274147 59533
rect 275461 59530 275527 59533
rect 274081 59528 275527 59530
rect 274081 59472 274086 59528
rect 274142 59472 275466 59528
rect 275522 59472 275527 59528
rect 274081 59470 275527 59472
rect 274081 59467 274147 59470
rect 275461 59467 275527 59470
rect 273897 59394 273963 59397
rect 276381 59394 276447 59397
rect 279344 59394 279404 60044
rect 280356 59394 280416 60044
rect 281368 59938 281428 60044
rect 273897 59392 276447 59394
rect 273897 59336 273902 59392
rect 273958 59336 276386 59392
rect 276442 59336 276447 59392
rect 273897 59334 276447 59336
rect 273897 59331 273963 59334
rect 276381 59331 276447 59334
rect 277350 59334 279404 59394
rect 279558 59334 280416 59394
rect 280478 59878 281428 59938
rect 269757 59256 272442 59258
rect 269757 59200 269762 59256
rect 269818 59200 272442 59256
rect 269757 59198 272442 59200
rect 276657 59258 276723 59261
rect 277350 59258 277410 59334
rect 276657 59256 277410 59258
rect 276657 59200 276662 59256
rect 276718 59200 277410 59256
rect 276657 59198 277410 59200
rect 278221 59258 278287 59261
rect 279558 59258 279618 59334
rect 278221 59256 279618 59258
rect 278221 59200 278226 59256
rect 278282 59200 279618 59256
rect 278221 59198 279618 59200
rect 259361 59195 259427 59198
rect 262857 59195 262923 59198
rect 268377 59195 268443 59198
rect 269757 59195 269823 59198
rect 276657 59195 276723 59198
rect 278221 59195 278287 59198
rect 237005 59120 238402 59122
rect 237005 59064 237010 59120
rect 237066 59064 238402 59120
rect 237005 59062 238402 59064
rect 278037 59122 278103 59125
rect 280478 59122 280538 59878
rect 280613 59802 280679 59805
rect 282380 59802 282440 60044
rect 280613 59800 282440 59802
rect 280613 59744 280618 59800
rect 280674 59744 282440 59800
rect 280613 59742 282440 59744
rect 280613 59739 280679 59742
rect 280797 59666 280863 59669
rect 283484 59666 283544 60044
rect 280797 59664 283544 59666
rect 280797 59608 280802 59664
rect 280858 59608 283544 59664
rect 280797 59606 283544 59608
rect 280797 59603 280863 59606
rect 282361 59530 282427 59533
rect 284496 59530 284556 60044
rect 282361 59528 284556 59530
rect 282361 59472 282366 59528
rect 282422 59472 284556 59528
rect 282361 59470 284556 59472
rect 284661 59530 284727 59533
rect 285508 59530 285568 60044
rect 284661 59528 285568 59530
rect 284661 59472 284666 59528
rect 284722 59472 285568 59528
rect 284661 59470 285568 59472
rect 282361 59467 282427 59470
rect 284661 59467 284727 59470
rect 283557 59394 283623 59397
rect 286520 59394 286580 60044
rect 286685 59666 286751 59669
rect 287624 59666 287684 60044
rect 286685 59664 287684 59666
rect 286685 59608 286690 59664
rect 286746 59608 287684 59664
rect 286685 59606 287684 59608
rect 286685 59603 286751 59606
rect 286685 59530 286751 59533
rect 288636 59530 288696 60044
rect 286685 59528 288696 59530
rect 286685 59472 286690 59528
rect 286746 59472 288696 59528
rect 286685 59470 288696 59472
rect 286685 59467 286751 59470
rect 289648 59394 289708 60044
rect 289813 59802 289879 59805
rect 290660 59802 290720 60044
rect 289813 59800 290720 59802
rect 289813 59744 289818 59800
rect 289874 59744 290720 59800
rect 289813 59742 290720 59744
rect 289813 59739 289879 59742
rect 291764 59666 291824 60044
rect 283557 59392 286580 59394
rect 283557 59336 283562 59392
rect 283618 59336 286580 59392
rect 283557 59334 286580 59336
rect 286734 59334 289708 59394
rect 289862 59606 291824 59666
rect 283557 59331 283623 59334
rect 286317 59258 286383 59261
rect 286734 59258 286794 59334
rect 286317 59256 286794 59258
rect 286317 59200 286322 59256
rect 286378 59200 286794 59256
rect 286317 59198 286794 59200
rect 289077 59258 289143 59261
rect 289862 59258 289922 59606
rect 290457 59530 290523 59533
rect 292776 59530 292836 60044
rect 292941 59802 293007 59805
rect 293788 59802 293848 60044
rect 292941 59800 293848 59802
rect 292941 59744 292946 59800
rect 293002 59744 293848 59800
rect 292941 59742 293848 59744
rect 292941 59739 293007 59742
rect 294800 59666 294860 60044
rect 290457 59528 292836 59530
rect 290457 59472 290462 59528
rect 290518 59472 292836 59528
rect 290457 59470 292836 59472
rect 292990 59606 294860 59666
rect 290457 59467 290523 59470
rect 291837 59394 291903 59397
rect 292990 59394 293050 59606
rect 293217 59530 293283 59533
rect 295904 59530 295964 60044
rect 293217 59528 295964 59530
rect 293217 59472 293222 59528
rect 293278 59472 295964 59528
rect 293217 59470 295964 59472
rect 296069 59530 296135 59533
rect 296916 59530 296976 60044
rect 297081 59802 297147 59805
rect 297928 59802 297988 60044
rect 297081 59800 297988 59802
rect 297081 59744 297086 59800
rect 297142 59744 297988 59800
rect 297081 59742 297988 59744
rect 297081 59739 297147 59742
rect 298940 59666 299000 60044
rect 296069 59528 296976 59530
rect 296069 59472 296074 59528
rect 296130 59472 296976 59528
rect 296069 59470 296976 59472
rect 297774 59606 299000 59666
rect 299105 59666 299171 59669
rect 300044 59666 300104 60044
rect 299105 59664 300104 59666
rect 299105 59608 299110 59664
rect 299166 59608 300104 59664
rect 299105 59606 300104 59608
rect 293217 59467 293283 59470
rect 296069 59467 296135 59470
rect 291837 59392 293050 59394
rect 291837 59336 291842 59392
rect 291898 59336 293050 59392
rect 291837 59334 293050 59336
rect 294781 59394 294847 59397
rect 295793 59394 295859 59397
rect 294781 59392 295859 59394
rect 294781 59336 294786 59392
rect 294842 59336 295798 59392
rect 295854 59336 295859 59392
rect 294781 59334 295859 59336
rect 291837 59331 291903 59334
rect 294781 59331 294847 59334
rect 295793 59331 295859 59334
rect 295977 59394 296043 59397
rect 297774 59394 297834 59606
rect 299105 59603 299171 59606
rect 298921 59530 298987 59533
rect 301056 59530 301116 60044
rect 302068 59938 302128 60044
rect 302006 59878 302128 59938
rect 302006 59802 302066 59878
rect 298921 59528 301116 59530
rect 298921 59472 298926 59528
rect 298982 59472 301116 59528
rect 298921 59470 301116 59472
rect 301454 59742 302066 59802
rect 302233 59802 302299 59805
rect 303080 59802 303140 60044
rect 302233 59800 303140 59802
rect 302233 59744 302238 59800
rect 302294 59744 303140 59800
rect 302233 59742 303140 59744
rect 298921 59467 298987 59470
rect 299105 59394 299171 59397
rect 295977 59392 297834 59394
rect 295977 59336 295982 59392
rect 296038 59336 297834 59392
rect 295977 59334 297834 59336
rect 297928 59392 299171 59394
rect 297928 59336 299110 59392
rect 299166 59336 299171 59392
rect 297928 59334 299171 59336
rect 295977 59331 296043 59334
rect 289077 59256 289922 59258
rect 289077 59200 289082 59256
rect 289138 59200 289922 59256
rect 289077 59198 289922 59200
rect 297357 59258 297423 59261
rect 297928 59258 297988 59334
rect 299105 59331 299171 59334
rect 297357 59256 297988 59258
rect 297357 59200 297362 59256
rect 297418 59200 297988 59256
rect 297357 59198 297988 59200
rect 298737 59258 298803 59261
rect 301454 59258 301514 59742
rect 302233 59739 302299 59742
rect 304092 59666 304152 60044
rect 302190 59606 304152 59666
rect 298737 59256 301514 59258
rect 298737 59200 298742 59256
rect 298798 59200 301514 59256
rect 298737 59198 301514 59200
rect 301589 59258 301655 59261
rect 302190 59258 302250 59606
rect 303337 59530 303403 59533
rect 305196 59530 305256 60044
rect 306208 59805 306268 60044
rect 306189 59800 306268 59805
rect 306189 59744 306194 59800
rect 306250 59744 306268 59800
rect 306189 59742 306268 59744
rect 306189 59739 306255 59742
rect 307220 59666 307280 60044
rect 303337 59528 305256 59530
rect 303337 59472 303342 59528
rect 303398 59472 305256 59528
rect 303337 59470 305256 59472
rect 305318 59606 307280 59666
rect 303337 59467 303403 59470
rect 304901 59394 304967 59397
rect 305318 59394 305378 59606
rect 308232 59530 308292 60044
rect 306330 59470 308292 59530
rect 306330 59397 306390 59470
rect 304901 59392 305378 59394
rect 304901 59336 304906 59392
rect 304962 59336 305378 59392
rect 304901 59334 305378 59336
rect 306281 59392 306390 59397
rect 306281 59336 306286 59392
rect 306342 59336 306390 59392
rect 306281 59334 306390 59336
rect 307569 59394 307635 59397
rect 309336 59394 309396 60044
rect 310348 59666 310408 60044
rect 310513 59802 310579 59805
rect 311360 59802 311420 60044
rect 310513 59800 311420 59802
rect 310513 59744 310518 59800
rect 310574 59744 311420 59800
rect 310513 59742 311420 59744
rect 310513 59739 310579 59742
rect 312372 59666 312432 60044
rect 307569 59392 309396 59394
rect 307569 59336 307574 59392
rect 307630 59336 309396 59392
rect 307569 59334 309396 59336
rect 309734 59606 310408 59666
rect 310470 59606 312432 59666
rect 304901 59331 304967 59334
rect 306281 59331 306347 59334
rect 307569 59331 307635 59334
rect 301589 59256 302250 59258
rect 301589 59200 301594 59256
rect 301650 59200 302250 59256
rect 301589 59198 302250 59200
rect 286317 59195 286383 59198
rect 289077 59195 289143 59198
rect 297357 59195 297423 59198
rect 298737 59195 298803 59198
rect 301589 59195 301655 59198
rect 278037 59120 280538 59122
rect 278037 59064 278042 59120
rect 278098 59064 280538 59120
rect 278037 59062 280538 59064
rect 307385 59122 307451 59125
rect 309734 59122 309794 59606
rect 310470 59533 310530 59606
rect 310421 59528 310530 59533
rect 310421 59472 310426 59528
rect 310482 59472 310530 59528
rect 310421 59470 310530 59472
rect 311801 59530 311867 59533
rect 313476 59530 313536 60044
rect 311801 59528 313536 59530
rect 311801 59472 311806 59528
rect 311862 59472 313536 59528
rect 311801 59470 313536 59472
rect 310421 59467 310487 59470
rect 311801 59467 311867 59470
rect 311617 59394 311683 59397
rect 314488 59394 314548 60044
rect 315500 59530 315560 60044
rect 316512 59666 316572 60044
rect 317616 59802 317676 60044
rect 318425 59802 318491 59805
rect 317616 59800 318491 59802
rect 317616 59744 318430 59800
rect 318486 59744 318491 59800
rect 317616 59742 318491 59744
rect 318425 59739 318491 59742
rect 316512 59606 318258 59666
rect 318057 59530 318123 59533
rect 315500 59528 318123 59530
rect 315500 59472 318062 59528
rect 318118 59472 318123 59528
rect 315500 59470 318123 59472
rect 318057 59467 318123 59470
rect 311617 59392 314548 59394
rect 311617 59336 311622 59392
rect 311678 59336 314548 59392
rect 311617 59334 314548 59336
rect 311617 59331 311683 59334
rect 318198 59258 318258 59606
rect 318628 59530 318688 60044
rect 319640 59666 319700 60044
rect 320449 59666 320515 59669
rect 319640 59664 320515 59666
rect 319640 59608 320454 59664
rect 320510 59608 320515 59664
rect 319640 59606 320515 59608
rect 320652 59666 320712 60044
rect 321756 59938 321816 60044
rect 321756 59878 322260 59938
rect 322200 59805 322260 59878
rect 322197 59800 322263 59805
rect 322197 59744 322202 59800
rect 322258 59744 322263 59800
rect 322197 59739 322263 59744
rect 322105 59666 322171 59669
rect 320652 59664 322171 59666
rect 320652 59608 322110 59664
rect 322166 59608 322171 59664
rect 320652 59606 322171 59608
rect 320449 59603 320515 59606
rect 322105 59603 322171 59606
rect 321001 59530 321067 59533
rect 318628 59528 321067 59530
rect 318628 59472 321006 59528
rect 321062 59472 321067 59528
rect 318628 59470 321067 59472
rect 321001 59467 321067 59470
rect 318425 59394 318491 59397
rect 320817 59394 320883 59397
rect 318425 59392 320883 59394
rect 318425 59336 318430 59392
rect 318486 59336 320822 59392
rect 320878 59336 320883 59392
rect 318425 59334 320883 59336
rect 322768 59394 322828 60044
rect 323780 59530 323840 60044
rect 324792 59666 324852 60044
rect 325896 59802 325956 60044
rect 326705 59802 326771 59805
rect 325896 59800 326771 59802
rect 325896 59744 326710 59800
rect 326766 59744 326771 59800
rect 325896 59742 326771 59744
rect 326705 59739 326771 59742
rect 324792 59606 326722 59666
rect 325693 59530 325759 59533
rect 323780 59528 325759 59530
rect 323780 59472 325698 59528
rect 325754 59472 325759 59528
rect 323780 59470 325759 59472
rect 325693 59467 325759 59470
rect 324957 59394 325023 59397
rect 322768 59392 325023 59394
rect 322768 59336 324962 59392
rect 325018 59336 325023 59392
rect 322768 59334 325023 59336
rect 326662 59394 326722 59606
rect 326908 59530 326968 60044
rect 327920 59666 327980 60044
rect 328729 59666 328795 59669
rect 327920 59664 328795 59666
rect 327920 59608 328734 59664
rect 328790 59608 328795 59664
rect 327920 59606 328795 59608
rect 328729 59603 328795 59606
rect 328729 59530 328795 59533
rect 326908 59528 328795 59530
rect 326908 59472 328734 59528
rect 328790 59472 328795 59528
rect 326908 59470 328795 59472
rect 328729 59467 328795 59470
rect 327717 59394 327783 59397
rect 326662 59392 327783 59394
rect 326662 59336 327722 59392
rect 327778 59336 327783 59392
rect 326662 59334 327783 59336
rect 328932 59394 328992 60044
rect 330036 59530 330096 60044
rect 330845 59530 330911 59533
rect 330036 59528 330911 59530
rect 330036 59472 330850 59528
rect 330906 59472 330911 59528
rect 330036 59470 330911 59472
rect 331048 59530 331108 60044
rect 331857 59530 331923 59533
rect 331048 59528 331923 59530
rect 331048 59472 331862 59528
rect 331918 59472 331923 59528
rect 331048 59470 331923 59472
rect 332060 59530 332120 60044
rect 333072 59666 333132 60044
rect 333881 59666 333947 59669
rect 333072 59664 333947 59666
rect 333072 59608 333886 59664
rect 333942 59608 333947 59664
rect 333072 59606 333947 59608
rect 334084 59666 334144 60044
rect 334084 59606 335002 59666
rect 333881 59603 333947 59606
rect 334617 59530 334683 59533
rect 332060 59528 334683 59530
rect 332060 59472 334622 59528
rect 334678 59472 334683 59528
rect 332060 59470 334683 59472
rect 330845 59467 330911 59470
rect 331857 59467 331923 59470
rect 334617 59467 334683 59470
rect 331857 59394 331923 59397
rect 333237 59394 333303 59397
rect 328932 59334 329850 59394
rect 318425 59331 318491 59334
rect 320817 59331 320883 59334
rect 324957 59331 325023 59334
rect 327717 59331 327783 59334
rect 319437 59258 319503 59261
rect 318198 59256 319503 59258
rect 318198 59200 319442 59256
rect 319498 59200 319503 59256
rect 318198 59198 319503 59200
rect 329790 59258 329850 59334
rect 330894 59392 331923 59394
rect 330894 59336 331862 59392
rect 331918 59336 331923 59392
rect 330894 59334 331923 59336
rect 330894 59258 330954 59334
rect 331857 59331 331923 59334
rect 331998 59392 333303 59394
rect 331998 59336 333242 59392
rect 333298 59336 333303 59392
rect 331998 59334 333303 59336
rect 329790 59198 330954 59258
rect 331029 59258 331095 59261
rect 331998 59258 332058 59334
rect 333237 59331 333303 59334
rect 333881 59394 333947 59397
rect 334942 59394 335002 59606
rect 335188 59530 335248 60044
rect 336200 59666 336260 60044
rect 337212 59802 337272 60044
rect 338021 59802 338087 59805
rect 337212 59800 338087 59802
rect 337212 59744 338026 59800
rect 338082 59744 338087 59800
rect 337212 59742 338087 59744
rect 338021 59739 338087 59742
rect 336200 59606 338130 59666
rect 337561 59530 337627 59533
rect 335188 59528 337627 59530
rect 335188 59472 337566 59528
rect 337622 59472 337627 59528
rect 335188 59470 337627 59472
rect 337561 59467 337627 59470
rect 337377 59394 337443 59397
rect 333881 59392 334818 59394
rect 333881 59336 333886 59392
rect 333942 59336 334818 59392
rect 333881 59334 334818 59336
rect 334942 59392 337443 59394
rect 334942 59336 337382 59392
rect 337438 59336 337443 59392
rect 334942 59334 337443 59336
rect 333881 59331 333947 59334
rect 331029 59256 332058 59258
rect 331029 59200 331034 59256
rect 331090 59200 332058 59256
rect 331029 59198 332058 59200
rect 334758 59258 334818 59334
rect 337377 59331 337443 59334
rect 335353 59258 335419 59261
rect 334758 59256 335419 59258
rect 334758 59200 335358 59256
rect 335414 59200 335419 59256
rect 334758 59198 335419 59200
rect 338070 59258 338130 59606
rect 338224 59394 338284 60044
rect 339328 59530 339388 60044
rect 340340 59666 340400 60044
rect 341352 59802 341412 60044
rect 342161 59802 342227 59805
rect 341352 59800 342227 59802
rect 341352 59744 342166 59800
rect 342222 59744 342227 59800
rect 341352 59742 342227 59744
rect 342161 59739 342227 59742
rect 340340 59606 342178 59666
rect 341517 59530 341583 59533
rect 339328 59528 341583 59530
rect 339328 59472 341522 59528
rect 341578 59472 341583 59528
rect 339328 59470 341583 59472
rect 341517 59467 341583 59470
rect 341701 59394 341767 59397
rect 338224 59392 341767 59394
rect 338224 59336 341706 59392
rect 341762 59336 341767 59392
rect 338224 59334 341767 59336
rect 341701 59331 341767 59334
rect 338757 59258 338823 59261
rect 338070 59256 338823 59258
rect 338070 59200 338762 59256
rect 338818 59200 338823 59256
rect 338070 59198 338823 59200
rect 342118 59258 342178 59606
rect 342364 59394 342424 60044
rect 343468 59530 343528 60044
rect 344480 59666 344540 60044
rect 345289 59666 345355 59669
rect 344480 59664 345355 59666
rect 344480 59608 345294 59664
rect 345350 59608 345355 59664
rect 344480 59606 345355 59608
rect 345289 59603 345355 59606
rect 345289 59530 345355 59533
rect 343468 59528 345355 59530
rect 343468 59472 345294 59528
rect 345350 59472 345355 59528
rect 343468 59470 345355 59472
rect 345289 59467 345355 59470
rect 345492 59394 345552 60044
rect 346504 59530 346564 60044
rect 347405 59530 347471 59533
rect 346504 59528 347471 59530
rect 346504 59472 347410 59528
rect 347466 59472 347471 59528
rect 346504 59470 347471 59472
rect 347608 59530 347668 60044
rect 348620 59666 348680 60044
rect 349632 59802 349692 60044
rect 350644 59938 350704 60044
rect 350644 59878 351378 59938
rect 351177 59802 351243 59805
rect 349632 59800 351243 59802
rect 349632 59744 351182 59800
rect 351238 59744 351243 59800
rect 349632 59742 351243 59744
rect 351177 59739 351243 59742
rect 351177 59666 351243 59669
rect 348620 59664 351243 59666
rect 348620 59608 351182 59664
rect 351238 59608 351243 59664
rect 348620 59606 351243 59608
rect 351177 59603 351243 59606
rect 349797 59530 349863 59533
rect 347608 59528 349863 59530
rect 347608 59472 349802 59528
rect 349858 59472 349863 59528
rect 347608 59470 349863 59472
rect 347405 59467 347471 59470
rect 349797 59467 349863 59470
rect 348417 59394 348483 59397
rect 349981 59394 350047 59397
rect 342364 59334 345306 59394
rect 345492 59392 348483 59394
rect 345492 59336 348422 59392
rect 348478 59336 348483 59392
rect 345492 59334 348483 59336
rect 342897 59258 342963 59261
rect 342118 59256 342963 59258
rect 342118 59200 342902 59256
rect 342958 59200 342963 59256
rect 342118 59198 342963 59200
rect 345246 59258 345306 59334
rect 348417 59331 348483 59334
rect 348558 59392 350047 59394
rect 348558 59336 349986 59392
rect 350042 59336 350047 59392
rect 348558 59334 350047 59336
rect 345841 59258 345907 59261
rect 345246 59256 345907 59258
rect 345246 59200 345846 59256
rect 345902 59200 345907 59256
rect 345246 59198 345907 59200
rect 319437 59195 319503 59198
rect 331029 59195 331095 59198
rect 335353 59195 335419 59198
rect 338757 59195 338823 59198
rect 342897 59195 342963 59198
rect 345841 59195 345907 59198
rect 347405 59258 347471 59261
rect 348558 59258 348618 59334
rect 349981 59331 350047 59334
rect 347405 59256 348618 59258
rect 347405 59200 347410 59256
rect 347466 59200 348618 59256
rect 347405 59198 348618 59200
rect 351318 59258 351378 59878
rect 351748 59530 351808 60044
rect 352760 59666 352820 60044
rect 353772 59802 353832 60044
rect 354784 59938 354844 60044
rect 354784 59878 355794 59938
rect 354673 59802 354739 59805
rect 353772 59800 354739 59802
rect 353772 59744 354678 59800
rect 354734 59744 354739 59800
rect 353772 59742 354739 59744
rect 354673 59739 354739 59742
rect 352760 59606 354690 59666
rect 353937 59530 354003 59533
rect 351748 59528 354003 59530
rect 351748 59472 353942 59528
rect 353998 59472 354003 59528
rect 351748 59470 354003 59472
rect 353937 59467 354003 59470
rect 351453 59394 351519 59397
rect 352557 59394 352623 59397
rect 351453 59392 352623 59394
rect 351453 59336 351458 59392
rect 351514 59336 352562 59392
rect 352618 59336 352623 59392
rect 351453 59334 352623 59336
rect 351453 59331 351519 59334
rect 352557 59331 352623 59334
rect 353293 59258 353359 59261
rect 351318 59256 353359 59258
rect 351318 59200 353298 59256
rect 353354 59200 353359 59256
rect 351318 59198 353359 59200
rect 354630 59258 354690 59606
rect 355734 59394 355794 59878
rect 355888 59530 355948 60044
rect 356900 59666 356960 60044
rect 357912 59802 357972 60044
rect 358924 59938 358984 60044
rect 359936 59938 359996 60044
rect 361040 59938 361100 60044
rect 358924 59878 359842 59938
rect 359936 59878 360026 59938
rect 361040 59878 361130 59938
rect 359457 59802 359523 59805
rect 357912 59800 359523 59802
rect 357912 59744 359462 59800
rect 359518 59744 359523 59800
rect 357912 59742 359523 59744
rect 359457 59739 359523 59742
rect 359457 59666 359523 59669
rect 359782 59666 359842 59878
rect 359966 59802 360026 59878
rect 360929 59802 360995 59805
rect 359966 59800 360995 59802
rect 359966 59744 360934 59800
rect 360990 59744 360995 59800
rect 359966 59742 360995 59744
rect 360929 59739 360995 59742
rect 361070 59666 361130 59878
rect 356900 59664 359523 59666
rect 356900 59608 359462 59664
rect 359518 59608 359523 59664
rect 356900 59606 359523 59608
rect 359457 59603 359523 59606
rect 359598 59606 359842 59666
rect 361040 59606 361130 59666
rect 362052 59666 362112 60044
rect 362861 59666 362927 59669
rect 362052 59664 362927 59666
rect 362052 59608 362866 59664
rect 362922 59608 362927 59664
rect 362052 59606 362927 59608
rect 363064 59666 363124 60044
rect 364076 59802 364136 60044
rect 365180 59938 365240 60044
rect 365180 59878 366098 59938
rect 364241 59802 364307 59805
rect 364076 59800 364307 59802
rect 364076 59744 364246 59800
rect 364302 59744 364307 59800
rect 364076 59742 364307 59744
rect 364241 59739 364307 59742
rect 365897 59666 365963 59669
rect 363064 59664 365963 59666
rect 363064 59608 365902 59664
rect 365958 59608 365963 59664
rect 363064 59606 365963 59608
rect 358261 59530 358327 59533
rect 355888 59528 358327 59530
rect 355888 59472 358266 59528
rect 358322 59472 358327 59528
rect 355888 59470 358327 59472
rect 358261 59467 358327 59470
rect 358077 59394 358143 59397
rect 355734 59392 358143 59394
rect 355734 59336 358082 59392
rect 358138 59336 358143 59392
rect 355734 59334 358143 59336
rect 359598 59394 359658 59606
rect 359733 59530 359799 59533
rect 360837 59530 360903 59533
rect 359733 59528 360903 59530
rect 359733 59472 359738 59528
rect 359794 59472 360842 59528
rect 360898 59472 360903 59528
rect 359733 59470 360903 59472
rect 361040 59530 361100 59606
rect 362861 59603 362927 59606
rect 365897 59603 365963 59606
rect 363597 59530 363663 59533
rect 361040 59528 363663 59530
rect 361040 59472 363602 59528
rect 363658 59472 363663 59528
rect 361040 59470 363663 59472
rect 359733 59467 359799 59470
rect 360837 59467 360903 59470
rect 363597 59467 363663 59470
rect 364241 59530 364307 59533
rect 365805 59530 365871 59533
rect 364241 59528 365871 59530
rect 364241 59472 364246 59528
rect 364302 59472 365810 59528
rect 365866 59472 365871 59528
rect 364241 59470 365871 59472
rect 364241 59467 364307 59470
rect 365805 59467 365871 59470
rect 360929 59394 360995 59397
rect 362217 59394 362283 59397
rect 359598 59334 360762 59394
rect 358077 59331 358143 59334
rect 355317 59258 355383 59261
rect 354630 59256 355383 59258
rect 354630 59200 355322 59256
rect 355378 59200 355383 59256
rect 354630 59198 355383 59200
rect 360702 59258 360762 59334
rect 360929 59392 362283 59394
rect 360929 59336 360934 59392
rect 360990 59336 362222 59392
rect 362278 59336 362283 59392
rect 360929 59334 362283 59336
rect 360929 59331 360995 59334
rect 362217 59331 362283 59334
rect 362861 59394 362927 59397
rect 364977 59394 365043 59397
rect 362861 59392 365043 59394
rect 362861 59336 362866 59392
rect 362922 59336 364982 59392
rect 365038 59336 365043 59392
rect 362861 59334 365043 59336
rect 366038 59394 366098 59878
rect 366192 59530 366252 60044
rect 367204 59666 367264 60044
rect 367204 59606 368122 59666
rect 367093 59530 367159 59533
rect 366192 59528 367159 59530
rect 366192 59472 367098 59528
rect 367154 59472 367159 59528
rect 366192 59470 367159 59472
rect 367093 59467 367159 59470
rect 367737 59394 367803 59397
rect 366038 59392 367803 59394
rect 366038 59336 367742 59392
rect 367798 59336 367803 59392
rect 366038 59334 367803 59336
rect 368062 59394 368122 59606
rect 368216 59530 368276 60044
rect 369320 59666 369380 60044
rect 370332 59802 370392 60044
rect 371141 59802 371207 59805
rect 370332 59800 371207 59802
rect 370332 59744 371146 59800
rect 371202 59744 371207 59800
rect 370332 59742 371207 59744
rect 371344 59802 371404 60044
rect 372356 59938 372416 60044
rect 373460 59938 373520 60044
rect 372356 59878 372538 59938
rect 372153 59802 372219 59805
rect 371344 59800 372219 59802
rect 371344 59744 372158 59800
rect 372214 59744 372219 59800
rect 371344 59742 372219 59744
rect 371141 59739 371207 59742
rect 372153 59739 372219 59742
rect 371233 59666 371299 59669
rect 372478 59666 372538 59878
rect 369320 59664 371299 59666
rect 369320 59608 371238 59664
rect 371294 59608 371299 59664
rect 369320 59606 371299 59608
rect 371233 59603 371299 59606
rect 372356 59606 372538 59666
rect 373398 59878 373520 59938
rect 373398 59666 373458 59878
rect 373717 59802 373783 59805
rect 374177 59802 374243 59805
rect 373717 59800 374243 59802
rect 373717 59744 373722 59800
rect 373778 59744 374182 59800
rect 374238 59744 374243 59800
rect 373717 59742 374243 59744
rect 373717 59739 373783 59742
rect 374177 59739 374243 59742
rect 373398 59606 373520 59666
rect 370129 59530 370195 59533
rect 368216 59528 370195 59530
rect 368216 59472 370134 59528
rect 370190 59472 370195 59528
rect 368216 59470 370195 59472
rect 370129 59467 370195 59470
rect 369945 59394 370011 59397
rect 368062 59392 370011 59394
rect 368062 59336 369950 59392
rect 370006 59336 370011 59392
rect 368062 59334 370011 59336
rect 362861 59331 362927 59334
rect 364977 59331 365043 59334
rect 367737 59331 367803 59334
rect 369945 59331 370011 59334
rect 371141 59394 371207 59397
rect 372356 59394 372416 59606
rect 373460 59394 373520 59606
rect 373993 59394 374059 59397
rect 374269 59394 374335 59397
rect 371141 59392 372170 59394
rect 371141 59336 371146 59392
rect 371202 59336 372170 59392
rect 371141 59334 372170 59336
rect 372356 59334 373274 59394
rect 373460 59392 374059 59394
rect 373460 59336 373998 59392
rect 374054 59336 374059 59392
rect 373460 59334 374059 59336
rect 371141 59331 371207 59334
rect 362125 59258 362191 59261
rect 360702 59256 362191 59258
rect 360702 59200 362130 59256
rect 362186 59200 362191 59256
rect 360702 59198 362191 59200
rect 372110 59258 372170 59334
rect 372705 59258 372771 59261
rect 372110 59256 372771 59258
rect 372110 59200 372710 59256
rect 372766 59200 372771 59256
rect 372110 59198 372771 59200
rect 373214 59258 373274 59334
rect 373993 59331 374059 59334
rect 374134 59392 374335 59394
rect 374134 59336 374274 59392
rect 374330 59336 374335 59392
rect 374134 59334 374335 59336
rect 374472 59394 374532 60044
rect 375484 59666 375544 60044
rect 376496 59805 376556 60044
rect 376477 59800 376556 59805
rect 376477 59744 376482 59800
rect 376538 59744 376556 59800
rect 376477 59742 376556 59744
rect 376753 59802 376819 59805
rect 377600 59802 377660 60044
rect 376753 59800 377660 59802
rect 376753 59744 376758 59800
rect 376814 59744 377660 59800
rect 376753 59742 377660 59744
rect 376477 59739 376543 59742
rect 376753 59739 376819 59742
rect 378409 59666 378475 59669
rect 375484 59664 378475 59666
rect 375484 59608 378414 59664
rect 378470 59608 378475 59664
rect 375484 59606 378475 59608
rect 378409 59603 378475 59606
rect 376477 59530 376543 59533
rect 378225 59530 378291 59533
rect 376477 59528 378291 59530
rect 376477 59472 376482 59528
rect 376538 59472 378230 59528
rect 378286 59472 378291 59528
rect 376477 59470 378291 59472
rect 376477 59467 376543 59470
rect 378225 59467 378291 59470
rect 376845 59394 376911 59397
rect 374472 59392 376911 59394
rect 374472 59336 376850 59392
rect 376906 59336 376911 59392
rect 374472 59334 376911 59336
rect 378612 59394 378672 60044
rect 379624 59394 379684 60044
rect 380636 59530 380696 60044
rect 381740 59666 381800 60044
rect 382752 59802 382812 60044
rect 383764 59938 383824 60044
rect 384776 59938 384836 60044
rect 383764 59878 384498 59938
rect 384776 59878 385096 59938
rect 384438 59805 384498 59878
rect 384113 59802 384179 59805
rect 382752 59800 384179 59802
rect 382752 59744 384118 59800
rect 384174 59744 384179 59800
rect 382752 59742 384179 59744
rect 384438 59800 384547 59805
rect 384438 59744 384486 59800
rect 384542 59744 384547 59800
rect 384438 59742 384547 59744
rect 384113 59739 384179 59742
rect 384481 59739 384547 59742
rect 383745 59666 383811 59669
rect 381740 59664 383811 59666
rect 381740 59608 383750 59664
rect 383806 59608 383811 59664
rect 381740 59606 383811 59608
rect 383745 59603 383811 59606
rect 382273 59530 382339 59533
rect 380636 59528 382339 59530
rect 380636 59472 382278 59528
rect 382334 59472 382339 59528
rect 380636 59470 382339 59472
rect 382273 59467 382339 59470
rect 382457 59394 382523 59397
rect 378612 59334 379530 59394
rect 379624 59392 382523 59394
rect 379624 59336 382462 59392
rect 382518 59336 382523 59392
rect 379624 59334 382523 59336
rect 374134 59258 374194 59334
rect 374269 59331 374335 59334
rect 376845 59331 376911 59334
rect 373214 59198 374194 59258
rect 379470 59258 379530 59334
rect 382457 59331 382523 59334
rect 380985 59258 381051 59261
rect 379470 59256 381051 59258
rect 379470 59200 380990 59256
rect 381046 59200 381051 59256
rect 379470 59198 381051 59200
rect 385036 59258 385096 59878
rect 385880 59530 385940 60044
rect 386892 59666 386952 60044
rect 387904 59802 387964 60044
rect 388713 59802 388779 59805
rect 387904 59800 388779 59802
rect 387904 59744 388718 59800
rect 388774 59744 388779 59800
rect 387904 59742 388779 59744
rect 388713 59739 388779 59742
rect 386892 59606 388730 59666
rect 387885 59530 387951 59533
rect 385880 59528 387951 59530
rect 385880 59472 387890 59528
rect 387946 59472 387951 59528
rect 385880 59470 387951 59472
rect 387885 59467 387951 59470
rect 385217 59394 385283 59397
rect 386597 59394 386663 59397
rect 385217 59392 386663 59394
rect 385217 59336 385222 59392
rect 385278 59336 386602 59392
rect 386658 59336 386663 59392
rect 385217 59334 386663 59336
rect 385217 59331 385283 59334
rect 386597 59331 386663 59334
rect 386413 59258 386479 59261
rect 385036 59256 386479 59258
rect 385036 59200 386418 59256
rect 386474 59200 386479 59256
rect 385036 59198 386479 59200
rect 388670 59258 388730 59606
rect 388916 59394 388976 60044
rect 389928 59938 389988 60044
rect 389130 59878 389834 59938
rect 389928 59878 390938 59938
rect 389130 59805 389190 59878
rect 389081 59800 389190 59805
rect 389081 59744 389086 59800
rect 389142 59744 389190 59800
rect 389081 59742 389190 59744
rect 389081 59739 389147 59742
rect 389774 59666 389834 59878
rect 390645 59666 390711 59669
rect 389774 59664 390711 59666
rect 389774 59608 390650 59664
rect 390706 59608 390711 59664
rect 389774 59606 390711 59608
rect 390645 59603 390711 59606
rect 390878 59530 390938 59878
rect 391032 59666 391092 60044
rect 392044 59802 392104 60044
rect 392853 59802 392919 59805
rect 392044 59800 392919 59802
rect 392044 59744 392858 59800
rect 392914 59744 392919 59800
rect 392044 59742 392919 59744
rect 392853 59739 392919 59742
rect 391032 59606 392226 59666
rect 392025 59530 392091 59533
rect 390878 59528 392091 59530
rect 390878 59472 392030 59528
rect 392086 59472 392091 59528
rect 390878 59470 392091 59472
rect 392025 59467 392091 59470
rect 390829 59394 390895 59397
rect 388916 59392 390895 59394
rect 388916 59336 390834 59392
rect 390890 59336 390895 59392
rect 388916 59334 390895 59336
rect 392166 59394 392226 59606
rect 393056 59530 393116 60044
rect 393056 59470 393882 59530
rect 393405 59394 393471 59397
rect 392166 59392 393471 59394
rect 392166 59336 393410 59392
rect 393466 59336 393471 59392
rect 392166 59334 393471 59336
rect 390829 59331 390895 59334
rect 393405 59331 393471 59334
rect 389265 59258 389331 59261
rect 388670 59256 389331 59258
rect 388670 59200 389270 59256
rect 389326 59200 389331 59256
rect 388670 59198 389331 59200
rect 393822 59258 393882 59470
rect 394068 59394 394128 60044
rect 394693 59530 394759 59533
rect 395172 59530 395232 60044
rect 394693 59528 395232 59530
rect 394693 59472 394698 59528
rect 394754 59472 395232 59528
rect 394693 59470 395232 59472
rect 394693 59467 394759 59470
rect 396184 59394 396244 60044
rect 397196 59530 397256 60044
rect 398208 59666 398268 60044
rect 399312 59802 399372 60044
rect 400121 59802 400187 59805
rect 399312 59800 400187 59802
rect 399312 59744 400126 59800
rect 400182 59744 400187 59800
rect 399312 59742 400187 59744
rect 400121 59739 400187 59742
rect 400324 59666 400384 60044
rect 398208 59606 400138 59666
rect 400324 59606 401058 59666
rect 399109 59530 399175 59533
rect 397196 59528 399175 59530
rect 397196 59472 399114 59528
rect 399170 59472 399175 59528
rect 397196 59470 399175 59472
rect 400078 59530 400138 59606
rect 400213 59530 400279 59533
rect 400078 59528 400279 59530
rect 400078 59472 400218 59528
rect 400274 59472 400279 59528
rect 400078 59470 400279 59472
rect 399109 59467 399175 59470
rect 400213 59467 400279 59470
rect 398925 59394 398991 59397
rect 394068 59334 396090 59394
rect 396184 59392 398991 59394
rect 396184 59336 398930 59392
rect 398986 59336 398991 59392
rect 396184 59334 398991 59336
rect 396030 59261 396090 59334
rect 398925 59331 398991 59334
rect 394785 59258 394851 59261
rect 393822 59256 394851 59258
rect 393822 59200 394790 59256
rect 394846 59200 394851 59256
rect 393822 59198 394851 59200
rect 396030 59256 396139 59261
rect 396030 59200 396078 59256
rect 396134 59200 396139 59256
rect 396030 59198 396139 59200
rect 400998 59258 401058 59606
rect 401336 59530 401396 60044
rect 402348 59666 402408 60044
rect 403452 59802 403512 60044
rect 404169 59802 404235 59805
rect 403452 59800 404235 59802
rect 403452 59744 404174 59800
rect 404230 59744 404235 59800
rect 403452 59742 404235 59744
rect 404169 59739 404235 59742
rect 404261 59666 404327 59669
rect 402348 59664 404327 59666
rect 402348 59608 404266 59664
rect 404322 59608 404327 59664
rect 402348 59606 404327 59608
rect 404261 59603 404327 59606
rect 403157 59530 403223 59533
rect 401336 59528 403223 59530
rect 401336 59472 403162 59528
rect 403218 59472 403223 59528
rect 401336 59470 403223 59472
rect 404464 59530 404524 60044
rect 405273 59530 405339 59533
rect 404464 59528 405339 59530
rect 404464 59472 405278 59528
rect 405334 59472 405339 59528
rect 404464 59470 405339 59472
rect 405476 59530 405536 60044
rect 406488 59666 406548 60044
rect 407592 59802 407652 60044
rect 408604 59938 408664 60044
rect 409616 59938 409676 60044
rect 408604 59878 409522 59938
rect 409616 59878 409706 59938
rect 409462 59805 409522 59878
rect 407592 59742 409338 59802
rect 409462 59800 409571 59805
rect 409462 59744 409510 59800
rect 409566 59744 409571 59800
rect 409462 59742 409571 59744
rect 408585 59666 408651 59669
rect 406488 59664 408651 59666
rect 406488 59608 408590 59664
rect 408646 59608 408651 59664
rect 406488 59606 408651 59608
rect 408585 59603 408651 59606
rect 407113 59530 407179 59533
rect 405476 59528 407179 59530
rect 405476 59472 407118 59528
rect 407174 59472 407179 59528
rect 405476 59470 407179 59472
rect 403157 59467 403223 59470
rect 405273 59467 405339 59470
rect 407113 59467 407179 59470
rect 402973 59394 403039 59397
rect 401734 59392 403039 59394
rect 401734 59336 402978 59392
rect 403034 59336 403039 59392
rect 401734 59334 403039 59336
rect 401734 59258 401794 59334
rect 402973 59331 403039 59334
rect 404169 59394 404235 59397
rect 405825 59394 405891 59397
rect 404169 59392 405891 59394
rect 404169 59336 404174 59392
rect 404230 59336 405830 59392
rect 405886 59336 405891 59392
rect 404169 59334 405891 59336
rect 409278 59394 409338 59742
rect 409505 59739 409571 59742
rect 409646 59666 409706 59878
rect 409616 59606 409706 59666
rect 409616 59394 409676 59606
rect 410628 59394 410688 60044
rect 411732 59802 411792 60044
rect 412744 59938 412804 60044
rect 412744 59878 413018 59938
rect 412633 59802 412699 59805
rect 411732 59800 412699 59802
rect 411732 59744 412638 59800
rect 412694 59744 412699 59800
rect 411732 59742 412699 59744
rect 412633 59739 412699 59742
rect 412958 59394 413018 59878
rect 413185 59530 413251 59533
rect 413756 59530 413816 60044
rect 413185 59528 413816 59530
rect 413185 59472 413190 59528
rect 413246 59472 413816 59528
rect 413185 59470 413816 59472
rect 414768 59530 414828 60044
rect 415872 59666 415932 60044
rect 416884 59802 416944 60044
rect 417896 59938 417956 60044
rect 418908 59938 418968 60044
rect 417896 59878 418722 59938
rect 418908 59878 419826 59938
rect 418662 59805 418722 59878
rect 416884 59742 418170 59802
rect 418662 59800 418771 59805
rect 418662 59744 418710 59800
rect 418766 59744 418771 59800
rect 418662 59742 418771 59744
rect 415872 59606 417802 59666
rect 416865 59530 416931 59533
rect 414768 59528 416931 59530
rect 414768 59472 416870 59528
rect 416926 59472 416931 59528
rect 414768 59470 416931 59472
rect 413185 59467 413251 59470
rect 416865 59467 416931 59470
rect 415577 59394 415643 59397
rect 409278 59334 409522 59394
rect 409616 59334 410442 59394
rect 410628 59334 412650 59394
rect 412958 59392 415643 59394
rect 412958 59336 415582 59392
rect 415638 59336 415643 59392
rect 412958 59334 415643 59336
rect 417742 59394 417802 59606
rect 418110 59530 418170 59742
rect 418705 59739 418771 59742
rect 419625 59530 419691 59533
rect 418110 59528 419691 59530
rect 418110 59472 419630 59528
rect 419686 59472 419691 59528
rect 418110 59470 419691 59472
rect 419625 59467 419691 59470
rect 418245 59394 418311 59397
rect 417742 59392 418311 59394
rect 417742 59336 418250 59392
rect 418306 59336 418311 59392
rect 417742 59334 418311 59336
rect 419766 59394 419826 59878
rect 419920 59530 419980 60044
rect 420821 59530 420887 59533
rect 419920 59528 420887 59530
rect 419920 59472 420826 59528
rect 420882 59472 420887 59528
rect 419920 59470 420887 59472
rect 420821 59467 420887 59470
rect 421024 59394 421084 60044
rect 422036 59530 422096 60044
rect 423048 59666 423108 60044
rect 423673 59802 423739 59805
rect 424060 59802 424120 60044
rect 423673 59800 424120 59802
rect 423673 59744 423678 59800
rect 423734 59744 424120 59800
rect 423673 59742 424120 59744
rect 423673 59739 423739 59742
rect 424961 59666 425027 59669
rect 423048 59664 425027 59666
rect 423048 59608 424966 59664
rect 425022 59608 425027 59664
rect 423048 59606 425027 59608
rect 424961 59603 425027 59606
rect 423857 59530 423923 59533
rect 422036 59528 423923 59530
rect 422036 59472 423862 59528
rect 423918 59472 423923 59528
rect 422036 59470 423923 59472
rect 423857 59467 423923 59470
rect 423765 59394 423831 59397
rect 419766 59334 420930 59394
rect 421024 59392 423831 59394
rect 421024 59336 423770 59392
rect 423826 59336 423831 59392
rect 421024 59334 423831 59336
rect 425164 59394 425224 60044
rect 425329 59530 425395 59533
rect 426176 59530 426236 60044
rect 425329 59528 426236 59530
rect 425329 59472 425334 59528
rect 425390 59472 426236 59528
rect 425329 59470 426236 59472
rect 427188 59530 427248 60044
rect 428200 59666 428260 60044
rect 429304 59802 429364 60044
rect 430113 59802 430179 59805
rect 429304 59800 430179 59802
rect 429304 59744 430118 59800
rect 430174 59744 430179 59800
rect 429304 59742 430179 59744
rect 430113 59739 430179 59742
rect 428200 59606 430130 59666
rect 429193 59530 429259 59533
rect 427188 59528 429259 59530
rect 427188 59472 429198 59528
rect 429254 59472 429259 59528
rect 427188 59470 429259 59472
rect 425329 59467 425395 59470
rect 429193 59467 429259 59470
rect 427997 59394 428063 59397
rect 425164 59392 428063 59394
rect 425164 59336 428002 59392
rect 428058 59336 428063 59392
rect 425164 59334 428063 59336
rect 430070 59394 430130 59606
rect 430316 59530 430376 60044
rect 431328 59938 431388 60044
rect 431328 59878 431418 59938
rect 431358 59666 431418 59878
rect 431493 59802 431559 59805
rect 431953 59802 432019 59805
rect 431493 59800 432019 59802
rect 431493 59744 431498 59800
rect 431554 59744 431958 59800
rect 432014 59744 432019 59800
rect 431493 59742 432019 59744
rect 432340 59802 432400 60044
rect 433149 59802 433215 59805
rect 432340 59800 433215 59802
rect 432340 59744 433154 59800
rect 433210 59744 433215 59800
rect 432340 59742 433215 59744
rect 431493 59739 431559 59742
rect 431953 59739 432019 59742
rect 433149 59739 433215 59742
rect 433241 59666 433307 59669
rect 431358 59664 433307 59666
rect 431358 59608 433246 59664
rect 433302 59608 433307 59664
rect 431358 59606 433307 59608
rect 433241 59603 433307 59606
rect 432137 59530 432203 59533
rect 430316 59528 432203 59530
rect 430316 59472 432142 59528
rect 432198 59472 432203 59528
rect 430316 59470 432203 59472
rect 433444 59530 433504 60044
rect 434253 59530 434319 59533
rect 433444 59528 434319 59530
rect 433444 59472 434258 59528
rect 434314 59472 434319 59528
rect 433444 59470 434319 59472
rect 434456 59530 434516 60044
rect 435468 59666 435528 60044
rect 436480 59802 436540 60044
rect 437584 59938 437644 60044
rect 438596 59938 438656 60044
rect 437584 59878 437674 59938
rect 438596 59878 439514 59938
rect 437473 59802 437539 59805
rect 436480 59800 437539 59802
rect 436480 59744 437478 59800
rect 437534 59744 437539 59800
rect 436480 59742 437539 59744
rect 437473 59739 437539 59742
rect 437381 59666 437447 59669
rect 437614 59666 437674 59878
rect 437749 59802 437815 59805
rect 438853 59802 438919 59805
rect 437749 59800 438919 59802
rect 437749 59744 437754 59800
rect 437810 59744 438858 59800
rect 438914 59744 438919 59800
rect 437749 59742 438919 59744
rect 437749 59739 437815 59742
rect 438853 59739 438919 59742
rect 435468 59664 437447 59666
rect 435468 59608 437386 59664
rect 437442 59608 437447 59664
rect 435468 59606 437447 59608
rect 437381 59603 437447 59606
rect 437584 59606 437674 59666
rect 436185 59530 436251 59533
rect 434456 59528 436251 59530
rect 434456 59472 436190 59528
rect 436246 59472 436251 59528
rect 434456 59470 436251 59472
rect 432137 59467 432203 59470
rect 434253 59467 434319 59470
rect 436185 59467 436251 59470
rect 430665 59394 430731 59397
rect 430070 59392 430731 59394
rect 430070 59336 430670 59392
rect 430726 59336 430731 59392
rect 430070 59334 430731 59336
rect 404169 59331 404235 59334
rect 405825 59331 405891 59334
rect 400998 59198 401794 59258
rect 409462 59258 409522 59334
rect 409965 59258 410031 59261
rect 409462 59256 410031 59258
rect 409462 59200 409970 59256
rect 410026 59200 410031 59256
rect 409462 59198 410031 59200
rect 410382 59258 410442 59334
rect 412590 59261 412650 59334
rect 415577 59331 415643 59334
rect 418245 59331 418311 59334
rect 411437 59258 411503 59261
rect 410382 59256 411503 59258
rect 410382 59200 411442 59256
rect 411498 59200 411503 59256
rect 410382 59198 411503 59200
rect 412590 59256 412699 59261
rect 412590 59200 412638 59256
rect 412694 59200 412699 59256
rect 412590 59198 412699 59200
rect 420870 59258 420930 59334
rect 423765 59331 423831 59334
rect 427997 59331 428063 59334
rect 430665 59331 430731 59334
rect 433149 59394 433215 59397
rect 434713 59394 434779 59397
rect 436369 59394 436435 59397
rect 433149 59392 434779 59394
rect 433149 59336 433154 59392
rect 433210 59336 434718 59392
rect 434774 59336 434779 59392
rect 433149 59334 434779 59336
rect 433149 59331 433215 59334
rect 434713 59331 434779 59334
rect 434854 59392 436435 59394
rect 434854 59336 436374 59392
rect 436430 59336 436435 59392
rect 434854 59334 436435 59336
rect 437584 59394 437644 59606
rect 439454 59394 439514 59878
rect 439608 59530 439668 60044
rect 440620 59666 440680 60044
rect 441061 59666 441127 59669
rect 440620 59664 441127 59666
rect 440620 59608 441066 59664
rect 441122 59608 441127 59664
rect 440620 59606 441127 59608
rect 441061 59603 441127 59606
rect 441724 59530 441784 60044
rect 442736 59666 442796 60044
rect 443748 59802 443808 60044
rect 444465 59802 444531 59805
rect 443748 59800 444531 59802
rect 443748 59744 444470 59800
rect 444526 59744 444531 59800
rect 443748 59742 444531 59744
rect 444465 59739 444531 59742
rect 444557 59666 444623 59669
rect 442736 59664 444623 59666
rect 442736 59608 444562 59664
rect 444618 59608 444623 59664
rect 442736 59606 444623 59608
rect 444760 59666 444820 60044
rect 445864 59802 445924 60044
rect 446673 59802 446739 59805
rect 445864 59800 446739 59802
rect 445864 59744 446678 59800
rect 446734 59744 446739 59800
rect 445864 59742 446739 59744
rect 446673 59739 446739 59742
rect 444760 59606 446690 59666
rect 444557 59603 444623 59606
rect 443545 59530 443611 59533
rect 439608 59470 441630 59530
rect 441724 59528 443611 59530
rect 441724 59472 443550 59528
rect 443606 59472 443611 59528
rect 441724 59470 443611 59472
rect 441061 59394 441127 59397
rect 441570 59394 441630 59470
rect 443545 59467 443611 59470
rect 444465 59530 444531 59533
rect 446397 59530 446463 59533
rect 444465 59528 446463 59530
rect 444465 59472 444470 59528
rect 444526 59472 446402 59528
rect 446458 59472 446463 59528
rect 444465 59470 446463 59472
rect 444465 59467 444531 59470
rect 446397 59467 446463 59470
rect 442257 59394 442323 59397
rect 443637 59394 443703 59397
rect 437584 59334 439330 59394
rect 439454 59334 440434 59394
rect 421005 59258 421071 59261
rect 420870 59256 421071 59258
rect 420870 59200 421010 59256
rect 421066 59200 421071 59256
rect 420870 59198 421071 59200
rect 347405 59195 347471 59198
rect 353293 59195 353359 59198
rect 355317 59195 355383 59198
rect 362125 59195 362191 59198
rect 372705 59195 372771 59198
rect 380985 59195 381051 59198
rect 386413 59195 386479 59198
rect 389265 59195 389331 59198
rect 394785 59195 394851 59198
rect 396073 59195 396139 59198
rect 409965 59195 410031 59198
rect 411437 59195 411503 59198
rect 412633 59195 412699 59198
rect 421005 59195 421071 59198
rect 434253 59258 434319 59261
rect 434854 59258 434914 59334
rect 436369 59331 436435 59334
rect 434253 59256 434914 59258
rect 434253 59200 434258 59256
rect 434314 59200 434914 59256
rect 434253 59198 434914 59200
rect 434253 59195 434319 59198
rect 307385 59120 309794 59122
rect 307385 59064 307390 59120
rect 307446 59064 309794 59120
rect 307385 59062 309794 59064
rect 439270 59122 439330 59334
rect 440374 59258 440434 59334
rect 441061 59392 441354 59394
rect 441061 59336 441066 59392
rect 441122 59336 441354 59392
rect 441061 59334 441354 59336
rect 441570 59392 442323 59394
rect 441570 59336 442262 59392
rect 442318 59336 442323 59392
rect 441570 59334 442323 59336
rect 441061 59331 441127 59334
rect 441061 59258 441127 59261
rect 440374 59256 441127 59258
rect 440374 59200 441066 59256
rect 441122 59200 441127 59256
rect 440374 59198 441127 59200
rect 441294 59258 441354 59334
rect 442257 59331 442323 59334
rect 442398 59392 443703 59394
rect 442398 59336 443642 59392
rect 443698 59336 443703 59392
rect 442398 59334 443703 59336
rect 446630 59394 446690 59606
rect 446876 59530 446936 60044
rect 447888 59666 447948 60044
rect 448697 59666 448763 59669
rect 447888 59664 448763 59666
rect 447888 59608 448702 59664
rect 448758 59608 448763 59664
rect 447888 59606 448763 59608
rect 448900 59666 448960 60044
rect 449709 59666 449775 59669
rect 448900 59664 449775 59666
rect 448900 59608 449714 59664
rect 449770 59608 449775 59664
rect 448900 59606 449775 59608
rect 448697 59603 448763 59606
rect 449709 59603 449775 59606
rect 449157 59530 449223 59533
rect 446876 59528 449223 59530
rect 446876 59472 449162 59528
rect 449218 59472 449223 59528
rect 446876 59470 449223 59472
rect 449157 59467 449223 59470
rect 447777 59394 447843 59397
rect 446630 59392 447843 59394
rect 446630 59336 447782 59392
rect 447838 59336 447843 59392
rect 446630 59334 447843 59336
rect 442398 59258 442458 59334
rect 443637 59331 443703 59334
rect 447777 59331 447843 59334
rect 448697 59394 448763 59397
rect 449912 59394 449972 60044
rect 451016 59394 451076 60044
rect 452028 59530 452088 60044
rect 453040 59666 453100 60044
rect 454052 59802 454112 60044
rect 454953 59802 455019 59805
rect 454052 59800 455019 59802
rect 454052 59744 454958 59800
rect 455014 59744 455019 59800
rect 454052 59742 455019 59744
rect 454953 59739 455019 59742
rect 453040 59606 454970 59666
rect 454677 59530 454743 59533
rect 452028 59528 454743 59530
rect 452028 59472 454682 59528
rect 454738 59472 454743 59528
rect 452028 59470 454743 59472
rect 454677 59467 454743 59470
rect 453297 59394 453363 59397
rect 448697 59392 449818 59394
rect 448697 59336 448702 59392
rect 448758 59336 449818 59392
rect 448697 59334 449818 59336
rect 449912 59334 450922 59394
rect 451016 59392 453363 59394
rect 451016 59336 453302 59392
rect 453358 59336 453363 59392
rect 451016 59334 453363 59336
rect 454910 59394 454970 59606
rect 455156 59530 455216 60044
rect 456168 59666 456228 60044
rect 457180 59802 457240 60044
rect 457989 59802 458055 59805
rect 457180 59800 458055 59802
rect 457180 59744 457994 59800
rect 458050 59744 458055 59800
rect 457180 59742 458055 59744
rect 457989 59739 458055 59742
rect 456168 59606 458098 59666
rect 457437 59530 457503 59533
rect 455156 59528 457503 59530
rect 455156 59472 457442 59528
rect 457498 59472 457503 59528
rect 455156 59470 457503 59472
rect 457437 59467 457503 59470
rect 456057 59394 456123 59397
rect 454910 59392 456123 59394
rect 454910 59336 456062 59392
rect 456118 59336 456123 59392
rect 454910 59334 456123 59336
rect 448697 59331 448763 59334
rect 441294 59198 442458 59258
rect 449758 59258 449818 59334
rect 450537 59258 450603 59261
rect 449758 59256 450603 59258
rect 449758 59200 450542 59256
rect 450598 59200 450603 59256
rect 449758 59198 450603 59200
rect 441061 59195 441127 59198
rect 450537 59195 450603 59198
rect 440877 59122 440943 59125
rect 439270 59120 440943 59122
rect 439270 59064 440882 59120
rect 440938 59064 440943 59120
rect 439270 59062 440943 59064
rect 450862 59122 450922 59334
rect 453297 59331 453363 59334
rect 456057 59331 456123 59334
rect 458038 59258 458098 59606
rect 458192 59394 458252 60044
rect 459296 59938 459356 60044
rect 459296 59878 460122 59938
rect 458357 59802 458423 59805
rect 459921 59802 459987 59805
rect 458357 59800 459987 59802
rect 458357 59744 458362 59800
rect 458418 59744 459926 59800
rect 459982 59744 459987 59800
rect 458357 59742 459987 59744
rect 458357 59739 458423 59742
rect 459921 59739 459987 59742
rect 460062 59530 460122 59878
rect 460308 59666 460368 60044
rect 461117 59666 461183 59669
rect 460308 59664 461183 59666
rect 460308 59608 461122 59664
rect 461178 59608 461183 59664
rect 460308 59606 461183 59608
rect 461117 59603 461183 59606
rect 461117 59530 461183 59533
rect 460062 59528 461183 59530
rect 460062 59472 461122 59528
rect 461178 59472 461183 59528
rect 460062 59470 461183 59472
rect 461117 59467 461183 59470
rect 461117 59394 461183 59397
rect 458192 59392 461183 59394
rect 458192 59336 461122 59392
rect 461178 59336 461183 59392
rect 458192 59334 461183 59336
rect 461320 59394 461380 60044
rect 462332 59530 462392 60044
rect 463233 59530 463299 59533
rect 462332 59528 463299 59530
rect 462332 59472 463238 59528
rect 463294 59472 463299 59528
rect 462332 59470 463299 59472
rect 463436 59530 463496 60044
rect 464448 59666 464508 60044
rect 465460 59802 465520 60044
rect 466472 59938 466532 60044
rect 467576 59938 467636 60044
rect 466472 59878 467482 59938
rect 467576 59878 467666 59938
rect 467281 59802 467347 59805
rect 465460 59800 467347 59802
rect 465460 59744 467286 59800
rect 467342 59744 467347 59800
rect 465460 59742 467347 59744
rect 467281 59739 467347 59742
rect 467097 59666 467163 59669
rect 464448 59664 467163 59666
rect 464448 59608 467102 59664
rect 467158 59608 467163 59664
rect 464448 59606 467163 59608
rect 467097 59603 467163 59606
rect 465717 59530 465783 59533
rect 463436 59528 465783 59530
rect 463436 59472 465722 59528
rect 465778 59472 465783 59528
rect 463436 59470 465783 59472
rect 463233 59467 463299 59470
rect 465717 59467 465783 59470
rect 464337 59394 464403 59397
rect 465901 59394 465967 59397
rect 461320 59392 464403 59394
rect 461320 59336 464342 59392
rect 464398 59336 464403 59392
rect 461320 59334 464403 59336
rect 461117 59331 461183 59334
rect 464337 59331 464403 59334
rect 464478 59392 465967 59394
rect 464478 59336 465906 59392
rect 465962 59336 465967 59392
rect 464478 59334 465967 59336
rect 458817 59258 458883 59261
rect 458038 59256 458883 59258
rect 458038 59200 458822 59256
rect 458878 59200 458883 59256
rect 458038 59198 458883 59200
rect 458817 59195 458883 59198
rect 463233 59258 463299 59261
rect 464478 59258 464538 59334
rect 465901 59331 465967 59334
rect 463233 59256 464538 59258
rect 463233 59200 463238 59256
rect 463294 59200 464538 59256
rect 463233 59198 464538 59200
rect 467422 59258 467482 59878
rect 467606 59666 467666 59878
rect 467576 59606 467666 59666
rect 467576 59394 467636 59606
rect 468588 59530 468648 60044
rect 469600 59666 469660 60044
rect 470612 59802 470672 60044
rect 471716 59938 471776 60044
rect 472728 59938 472788 60044
rect 471716 59878 472634 59938
rect 472728 59878 473554 59938
rect 470612 59742 472450 59802
rect 471973 59666 472039 59669
rect 469600 59664 472039 59666
rect 469600 59608 471978 59664
rect 472034 59608 472039 59664
rect 469600 59606 472039 59608
rect 471973 59603 472039 59606
rect 470685 59530 470751 59533
rect 468588 59528 470751 59530
rect 468588 59472 470690 59528
rect 470746 59472 470751 59528
rect 468588 59470 470751 59472
rect 470685 59467 470751 59470
rect 469857 59394 469923 59397
rect 467576 59392 469923 59394
rect 467576 59336 469862 59392
rect 469918 59336 469923 59392
rect 467576 59334 469923 59336
rect 472390 59394 472450 59742
rect 472574 59666 472634 59878
rect 473353 59666 473419 59669
rect 472574 59664 473419 59666
rect 472574 59608 473358 59664
rect 473414 59608 473419 59664
rect 472574 59606 473419 59608
rect 473353 59603 473419 59606
rect 473494 59530 473554 59878
rect 473740 59666 473800 60044
rect 474549 59666 474615 59669
rect 473740 59664 474615 59666
rect 473740 59608 474554 59664
rect 474610 59608 474615 59664
rect 473740 59606 474615 59608
rect 474752 59666 474812 60044
rect 475856 59802 475916 60044
rect 476868 59938 476928 60044
rect 476868 59878 477786 59938
rect 476021 59802 476087 59805
rect 475856 59800 476087 59802
rect 475856 59744 476026 59800
rect 476082 59744 476087 59800
rect 475856 59742 476087 59744
rect 476021 59739 476087 59742
rect 477585 59666 477651 59669
rect 474752 59664 477651 59666
rect 474752 59608 477590 59664
rect 477646 59608 477651 59664
rect 474752 59606 477651 59608
rect 474549 59603 474615 59606
rect 477585 59603 477651 59606
rect 474733 59530 474799 59533
rect 473494 59528 474799 59530
rect 473494 59472 474738 59528
rect 474794 59472 474799 59528
rect 473494 59470 474799 59472
rect 474733 59467 474799 59470
rect 476021 59530 476087 59533
rect 477726 59530 477786 59878
rect 477880 59666 477940 60044
rect 478892 59802 478952 60044
rect 479904 59938 479964 60044
rect 481008 59938 481068 60044
rect 479904 59878 480914 59938
rect 481008 59878 481880 59938
rect 478892 59742 480730 59802
rect 480253 59666 480319 59669
rect 477880 59664 480319 59666
rect 477880 59608 480258 59664
rect 480314 59608 480319 59664
rect 477880 59606 480319 59608
rect 480253 59603 480319 59606
rect 478873 59530 478939 59533
rect 476021 59528 476682 59530
rect 476021 59472 476026 59528
rect 476082 59472 476682 59528
rect 476021 59470 476682 59472
rect 477726 59528 478939 59530
rect 477726 59472 478878 59528
rect 478934 59472 478939 59528
rect 477726 59470 478939 59472
rect 476021 59467 476087 59470
rect 473537 59394 473603 59397
rect 472390 59392 473603 59394
rect 472390 59336 473542 59392
rect 473598 59336 473603 59392
rect 472390 59334 473603 59336
rect 469857 59331 469923 59334
rect 473537 59331 473603 59334
rect 474549 59394 474615 59397
rect 476205 59394 476271 59397
rect 474549 59392 476271 59394
rect 474549 59336 474554 59392
rect 474610 59336 476210 59392
rect 476266 59336 476271 59392
rect 474549 59334 476271 59336
rect 476622 59394 476682 59470
rect 478873 59467 478939 59470
rect 477585 59394 477651 59397
rect 476622 59392 477651 59394
rect 476622 59336 477590 59392
rect 477646 59336 477651 59392
rect 476622 59334 477651 59336
rect 480670 59394 480730 59742
rect 480854 59666 480914 59878
rect 481633 59666 481699 59669
rect 480854 59664 481699 59666
rect 480854 59608 481638 59664
rect 481694 59608 481699 59664
rect 480854 59606 481699 59608
rect 481633 59603 481699 59606
rect 481820 59530 481880 59878
rect 482020 59666 482080 60044
rect 482829 59666 482895 59669
rect 482020 59664 482895 59666
rect 482020 59608 482834 59664
rect 482890 59608 482895 59664
rect 482020 59606 482895 59608
rect 483032 59666 483092 60044
rect 484044 59802 484104 60044
rect 484853 59802 484919 59805
rect 484044 59800 484919 59802
rect 484044 59744 484858 59800
rect 484914 59744 484919 59800
rect 484044 59742 484919 59744
rect 485148 59802 485208 60044
rect 486160 59938 486220 60044
rect 487172 59938 487232 60044
rect 488184 59938 488244 60044
rect 489288 59938 489348 60044
rect 486160 59878 486250 59938
rect 487172 59878 488090 59938
rect 488184 59878 489010 59938
rect 485773 59802 485839 59805
rect 485148 59800 485839 59802
rect 485148 59744 485778 59800
rect 485834 59744 485839 59800
rect 485148 59742 485839 59744
rect 484853 59739 484919 59742
rect 485773 59739 485839 59742
rect 485957 59666 486023 59669
rect 483032 59664 486023 59666
rect 483032 59608 485962 59664
rect 486018 59608 486023 59664
rect 483032 59606 486023 59608
rect 486190 59666 486250 59878
rect 488030 59805 488090 59878
rect 488030 59800 488139 59805
rect 488030 59744 488078 59800
rect 488134 59744 488139 59800
rect 488030 59742 488139 59744
rect 488073 59739 488139 59742
rect 486190 59606 488090 59666
rect 482829 59603 482895 59606
rect 485957 59603 486023 59606
rect 483013 59530 483079 59533
rect 481820 59528 483079 59530
rect 481820 59472 483018 59528
rect 483074 59472 483079 59528
rect 481820 59470 483079 59472
rect 483013 59467 483079 59470
rect 484853 59530 484919 59533
rect 486141 59530 486207 59533
rect 484853 59528 486207 59530
rect 484853 59472 484858 59528
rect 484914 59472 486146 59528
rect 486202 59472 486207 59528
rect 484853 59470 486207 59472
rect 484853 59467 484919 59470
rect 486141 59467 486207 59470
rect 481817 59394 481883 59397
rect 480670 59392 481883 59394
rect 480670 59336 481822 59392
rect 481878 59336 481883 59392
rect 480670 59334 481883 59336
rect 474549 59331 474615 59334
rect 476205 59331 476271 59334
rect 477585 59331 477651 59334
rect 481817 59331 481883 59334
rect 482829 59394 482895 59397
rect 484485 59394 484551 59397
rect 482829 59392 484551 59394
rect 482829 59336 482834 59392
rect 482890 59336 484490 59392
rect 484546 59336 484551 59392
rect 482829 59334 484551 59336
rect 482829 59331 482895 59334
rect 484485 59331 484551 59334
rect 485773 59394 485839 59397
rect 487245 59394 487311 59397
rect 485773 59392 487311 59394
rect 485773 59336 485778 59392
rect 485834 59336 487250 59392
rect 487306 59336 487311 59392
rect 485773 59334 487311 59336
rect 488030 59394 488090 59606
rect 488950 59530 489010 59878
rect 489134 59878 489348 59938
rect 489134 59666 489194 59878
rect 489361 59802 489427 59805
rect 490097 59802 490163 59805
rect 489361 59800 490163 59802
rect 489361 59744 489366 59800
rect 489422 59744 490102 59800
rect 490158 59744 490163 59800
rect 489361 59742 490163 59744
rect 490300 59802 490360 60044
rect 491017 59802 491083 59805
rect 490300 59800 491083 59802
rect 490300 59744 491022 59800
rect 491078 59744 491083 59800
rect 490300 59742 491083 59744
rect 489361 59739 489427 59742
rect 490097 59739 490163 59742
rect 491017 59739 491083 59742
rect 491109 59666 491175 59669
rect 489134 59664 491175 59666
rect 489134 59608 491114 59664
rect 491170 59608 491175 59664
rect 489134 59606 491175 59608
rect 491109 59603 491175 59606
rect 489913 59530 489979 59533
rect 488950 59528 489979 59530
rect 488950 59472 489918 59528
rect 489974 59472 489979 59528
rect 488950 59470 489979 59472
rect 491312 59530 491372 60044
rect 492121 59530 492187 59533
rect 491312 59528 492187 59530
rect 491312 59472 492126 59528
rect 492182 59472 492187 59528
rect 491312 59470 492187 59472
rect 492324 59530 492384 60044
rect 493428 59666 493488 60044
rect 493428 59606 494346 59666
rect 494053 59530 494119 59533
rect 492324 59528 494119 59530
rect 492324 59472 494058 59528
rect 494114 59472 494119 59528
rect 492324 59470 494119 59472
rect 489913 59467 489979 59470
rect 492121 59467 492187 59470
rect 494053 59467 494119 59470
rect 488625 59394 488691 59397
rect 488030 59392 488691 59394
rect 488030 59336 488630 59392
rect 488686 59336 488691 59392
rect 488030 59334 488691 59336
rect 485773 59331 485839 59334
rect 487245 59331 487311 59334
rect 488625 59331 488691 59334
rect 491017 59394 491083 59397
rect 492673 59394 492739 59397
rect 491017 59392 492739 59394
rect 491017 59336 491022 59392
rect 491078 59336 492678 59392
rect 492734 59336 492739 59392
rect 491017 59334 492739 59336
rect 494286 59394 494346 59606
rect 494440 59530 494500 60044
rect 495452 59666 495512 60044
rect 495617 59802 495683 59805
rect 496464 59802 496524 60044
rect 495617 59800 496524 59802
rect 495617 59744 495622 59800
rect 495678 59744 496524 59800
rect 495617 59742 496524 59744
rect 497568 59802 497628 60044
rect 498580 59938 498640 60044
rect 498580 59878 499498 59938
rect 498469 59802 498535 59805
rect 497568 59800 498535 59802
rect 497568 59744 498474 59800
rect 498530 59744 498535 59800
rect 497568 59742 498535 59744
rect 495617 59739 495683 59742
rect 498469 59739 498535 59742
rect 498377 59666 498443 59669
rect 495452 59664 498443 59666
rect 495452 59608 498382 59664
rect 498438 59608 498443 59664
rect 495452 59606 498443 59608
rect 498377 59603 498443 59606
rect 496813 59530 496879 59533
rect 494440 59528 496879 59530
rect 494440 59472 496818 59528
rect 496874 59472 496879 59528
rect 494440 59470 496879 59472
rect 496813 59467 496879 59470
rect 495525 59394 495591 59397
rect 494286 59392 495591 59394
rect 494286 59336 495530 59392
rect 495586 59336 495591 59392
rect 494286 59334 495591 59336
rect 491017 59331 491083 59334
rect 492673 59331 492739 59334
rect 495525 59331 495591 59334
rect 469213 59258 469279 59261
rect 467422 59256 469279 59258
rect 467422 59200 469218 59256
rect 469274 59200 469279 59256
rect 467422 59198 469279 59200
rect 499438 59258 499498 59878
rect 499592 59394 499652 60044
rect 500604 59530 500664 60044
rect 501708 59666 501768 60044
rect 502720 59938 502780 60044
rect 502720 59878 503546 59938
rect 501708 59606 503362 59666
rect 502701 59530 502767 59533
rect 500604 59528 502767 59530
rect 500604 59472 502706 59528
rect 502762 59472 502767 59528
rect 500604 59470 502767 59472
rect 502701 59467 502767 59470
rect 502517 59394 502583 59397
rect 499592 59392 502583 59394
rect 499592 59336 502522 59392
rect 502578 59336 502583 59392
rect 499592 59334 502583 59336
rect 502517 59331 502583 59334
rect 501045 59258 501111 59261
rect 499438 59256 501111 59258
rect 499438 59200 501050 59256
rect 501106 59200 501111 59256
rect 499438 59198 501111 59200
rect 503302 59258 503362 59606
rect 503486 59394 503546 59878
rect 503732 59530 503792 60044
rect 504744 59938 504804 60044
rect 505848 59938 505908 60044
rect 504590 59878 504804 59938
rect 505694 59878 505908 59938
rect 504590 59666 504650 59878
rect 505694 59666 505754 59878
rect 506860 59802 506920 60044
rect 507872 59938 507932 60044
rect 507872 59878 508698 59938
rect 508638 59805 508698 59878
rect 506860 59742 508146 59802
rect 508638 59800 508747 59805
rect 508638 59744 508686 59800
rect 508742 59744 508747 59800
rect 508638 59742 508747 59744
rect 507853 59666 507919 59669
rect 504590 59606 504804 59666
rect 505694 59664 507919 59666
rect 505694 59608 507858 59664
rect 507914 59608 507919 59664
rect 505694 59606 507919 59608
rect 504541 59530 504607 59533
rect 503732 59528 504607 59530
rect 503732 59472 504546 59528
rect 504602 59472 504607 59528
rect 503732 59470 504607 59472
rect 504744 59530 504804 59606
rect 507853 59603 507919 59606
rect 506473 59530 506539 59533
rect 504744 59528 506539 59530
rect 504744 59472 506478 59528
rect 506534 59472 506539 59528
rect 504744 59470 506539 59472
rect 504541 59467 504607 59470
rect 506473 59467 506539 59470
rect 505185 59394 505251 59397
rect 503486 59392 505251 59394
rect 503486 59336 505190 59392
rect 505246 59336 505251 59392
rect 503486 59334 505251 59336
rect 508086 59394 508146 59742
rect 508681 59739 508747 59742
rect 508884 59530 508944 60044
rect 509896 59938 509956 60044
rect 509896 59878 510906 59938
rect 509049 59802 509115 59805
rect 509049 59800 509250 59802
rect 509049 59744 509054 59800
rect 509110 59744 509250 59800
rect 509049 59742 509250 59744
rect 509049 59739 509115 59742
rect 509190 59666 509250 59742
rect 510705 59666 510771 59669
rect 509190 59664 510771 59666
rect 509190 59608 510710 59664
rect 510766 59608 510771 59664
rect 509190 59606 510771 59608
rect 510705 59603 510771 59606
rect 510846 59530 510906 59878
rect 511000 59666 511060 60044
rect 512012 59802 512072 60044
rect 512821 59802 512887 59805
rect 512012 59800 512887 59802
rect 512012 59744 512826 59800
rect 512882 59744 512887 59800
rect 512012 59742 512887 59744
rect 512821 59739 512887 59742
rect 511000 59606 512930 59666
rect 511993 59530 512059 59533
rect 508884 59470 509802 59530
rect 510846 59528 512059 59530
rect 510846 59472 511998 59528
rect 512054 59472 512059 59528
rect 510846 59470 512059 59472
rect 509233 59394 509299 59397
rect 508086 59392 509299 59394
rect 508086 59336 509238 59392
rect 509294 59336 509299 59392
rect 508086 59334 509299 59336
rect 509742 59394 509802 59470
rect 511993 59467 512059 59470
rect 510705 59394 510771 59397
rect 509742 59392 510771 59394
rect 509742 59336 510710 59392
rect 510766 59336 510771 59392
rect 509742 59334 510771 59336
rect 512870 59394 512930 59606
rect 513024 59530 513084 60044
rect 514036 59666 514096 60044
rect 515140 59802 515200 60044
rect 515949 59802 516015 59805
rect 515140 59800 516015 59802
rect 515140 59744 515954 59800
rect 516010 59744 516015 59800
rect 515140 59742 516015 59744
rect 516152 59802 516212 60044
rect 516961 59802 517027 59805
rect 516152 59800 517027 59802
rect 516152 59744 516966 59800
rect 517022 59744 517027 59800
rect 516152 59742 517027 59744
rect 515949 59739 516015 59742
rect 516961 59739 517027 59742
rect 516133 59666 516199 59669
rect 514036 59664 516199 59666
rect 514036 59608 516138 59664
rect 516194 59608 516199 59664
rect 514036 59606 516199 59608
rect 516133 59603 516199 59606
rect 515029 59530 515095 59533
rect 513024 59528 515095 59530
rect 513024 59472 515034 59528
rect 515090 59472 515095 59528
rect 513024 59470 515095 59472
rect 517164 59530 517224 60044
rect 518176 59938 518236 60044
rect 518176 59878 518266 59938
rect 518206 59666 518266 59878
rect 518341 59802 518407 59805
rect 518985 59802 519051 59805
rect 518341 59800 519051 59802
rect 518341 59744 518346 59800
rect 518402 59744 518990 59800
rect 519046 59744 519051 59800
rect 518341 59742 519051 59744
rect 519280 59802 519340 60044
rect 520089 59802 520155 59805
rect 519280 59800 520155 59802
rect 519280 59744 520094 59800
rect 520150 59744 520155 59800
rect 519280 59742 520155 59744
rect 518341 59739 518407 59742
rect 518985 59739 519051 59742
rect 520089 59739 520155 59742
rect 520292 59666 520352 60044
rect 521304 59802 521364 60044
rect 522021 59802 522087 59805
rect 521304 59800 522087 59802
rect 521304 59744 522026 59800
rect 522082 59744 522087 59800
rect 521304 59742 522087 59744
rect 522021 59739 522087 59742
rect 522113 59666 522179 59669
rect 518206 59606 519738 59666
rect 520292 59664 522179 59666
rect 520292 59608 522118 59664
rect 522174 59608 522179 59664
rect 520292 59606 522179 59608
rect 522316 59666 522376 60044
rect 523420 59802 523480 60044
rect 524229 59802 524295 59805
rect 523420 59800 524295 59802
rect 523420 59744 524234 59800
rect 524290 59744 524295 59800
rect 523420 59742 524295 59744
rect 524432 59802 524492 60044
rect 525241 59802 525307 59805
rect 524432 59800 525307 59802
rect 524432 59744 525246 59800
rect 525302 59744 525307 59800
rect 524432 59742 525307 59744
rect 524229 59739 524295 59742
rect 525241 59739 525307 59742
rect 524505 59666 524571 59669
rect 522316 59664 524571 59666
rect 522316 59608 524510 59664
rect 524566 59608 524571 59664
rect 522316 59606 524571 59608
rect 519077 59530 519143 59533
rect 517164 59528 519143 59530
rect 517164 59472 519082 59528
rect 519138 59472 519143 59528
rect 517164 59470 519143 59472
rect 519678 59530 519738 59606
rect 522113 59603 522179 59606
rect 524505 59603 524571 59606
rect 520365 59530 520431 59533
rect 519678 59528 520431 59530
rect 519678 59472 520370 59528
rect 520426 59472 520431 59528
rect 519678 59470 520431 59472
rect 515029 59467 515095 59470
rect 519077 59467 519143 59470
rect 520365 59467 520431 59470
rect 522021 59530 522087 59533
rect 523033 59530 523099 59533
rect 522021 59528 523099 59530
rect 522021 59472 522026 59528
rect 522082 59472 523038 59528
rect 523094 59472 523099 59528
rect 522021 59470 523099 59472
rect 522021 59467 522087 59470
rect 523033 59467 523099 59470
rect 513465 59394 513531 59397
rect 512870 59392 513531 59394
rect 512870 59336 513470 59392
rect 513526 59336 513531 59392
rect 512870 59334 513531 59336
rect 505185 59331 505251 59334
rect 509233 59331 509299 59334
rect 510705 59331 510771 59334
rect 513465 59331 513531 59334
rect 515949 59394 516015 59397
rect 517605 59394 517671 59397
rect 515949 59392 517671 59394
rect 515949 59336 515954 59392
rect 516010 59336 517610 59392
rect 517666 59336 517671 59392
rect 515949 59334 517671 59336
rect 515949 59331 516015 59334
rect 517605 59331 517671 59334
rect 520089 59394 520155 59397
rect 521745 59394 521811 59397
rect 520089 59392 521811 59394
rect 520089 59336 520094 59392
rect 520150 59336 521750 59392
rect 521806 59336 521811 59392
rect 520089 59334 521811 59336
rect 520089 59331 520155 59334
rect 521745 59331 521811 59334
rect 522113 59394 522179 59397
rect 523217 59394 523283 59397
rect 522113 59392 523283 59394
rect 522113 59336 522118 59392
rect 522174 59336 523222 59392
rect 523278 59336 523283 59392
rect 522113 59334 523283 59336
rect 522113 59331 522179 59334
rect 523217 59331 523283 59334
rect 524229 59394 524295 59397
rect 525444 59394 525504 60044
rect 526456 59394 526516 60044
rect 527560 59802 527620 60044
rect 528572 59938 528632 60044
rect 528572 59878 528754 59938
rect 528694 59805 528754 59878
rect 527560 59742 528570 59802
rect 528510 59666 528570 59742
rect 528645 59800 528754 59805
rect 528645 59744 528650 59800
rect 528706 59744 528754 59800
rect 528645 59742 528754 59744
rect 528645 59739 528711 59742
rect 528510 59606 528754 59666
rect 528553 59394 528619 59397
rect 524229 59392 525258 59394
rect 524229 59336 524234 59392
rect 524290 59336 525258 59392
rect 524229 59334 525258 59336
rect 525444 59334 526362 59394
rect 526456 59392 528619 59394
rect 526456 59336 528558 59392
rect 528614 59336 528619 59392
rect 526456 59334 528619 59336
rect 528694 59394 528754 59606
rect 529013 59530 529079 59533
rect 529584 59530 529644 60044
rect 529013 59528 529644 59530
rect 529013 59472 529018 59528
rect 529074 59472 529644 59528
rect 529013 59470 529644 59472
rect 530596 59530 530656 60044
rect 531700 59666 531760 60044
rect 532712 59802 532772 60044
rect 533724 59938 533784 60044
rect 533724 59878 533906 59938
rect 533705 59802 533771 59805
rect 532712 59800 533771 59802
rect 532712 59744 533710 59800
rect 533766 59744 533771 59800
rect 532712 59742 533771 59744
rect 533705 59739 533771 59742
rect 533846 59666 533906 59878
rect 531700 59606 533538 59666
rect 532693 59530 532759 59533
rect 530596 59528 532759 59530
rect 530596 59472 532698 59528
rect 532754 59472 532759 59528
rect 530596 59470 532759 59472
rect 529013 59467 529079 59470
rect 532693 59467 532759 59470
rect 529933 59394 529999 59397
rect 528694 59392 529999 59394
rect 528694 59336 529938 59392
rect 529994 59336 529999 59392
rect 528694 59334 529999 59336
rect 533478 59394 533538 59606
rect 533724 59606 533906 59666
rect 534736 59666 534796 60044
rect 535545 59666 535611 59669
rect 534736 59664 535611 59666
rect 534736 59608 535550 59664
rect 535606 59608 535611 59664
rect 534736 59606 535611 59608
rect 535840 59666 535900 60044
rect 536852 59802 536912 60044
rect 537661 59802 537727 59805
rect 536852 59800 537727 59802
rect 536852 59744 537666 59800
rect 537722 59744 537727 59800
rect 536852 59742 537727 59744
rect 537661 59739 537727 59742
rect 535840 59606 537034 59666
rect 533724 59530 533784 59606
rect 535545 59603 535611 59606
rect 535821 59530 535887 59533
rect 533724 59528 535887 59530
rect 533724 59472 535826 59528
rect 535882 59472 535887 59528
rect 533724 59470 535887 59472
rect 535821 59467 535887 59470
rect 534073 59394 534139 59397
rect 533478 59392 534139 59394
rect 533478 59336 534078 59392
rect 534134 59336 534139 59392
rect 533478 59334 534139 59336
rect 524229 59331 524295 59334
rect 503805 59258 503871 59261
rect 503302 59256 503871 59258
rect 503302 59200 503810 59256
rect 503866 59200 503871 59256
rect 503302 59198 503871 59200
rect 525198 59258 525258 59334
rect 525793 59258 525859 59261
rect 525198 59256 525859 59258
rect 525198 59200 525798 59256
rect 525854 59200 525859 59256
rect 525198 59198 525859 59200
rect 526302 59258 526362 59334
rect 528553 59331 528619 59334
rect 529933 59331 529999 59334
rect 534073 59331 534139 59334
rect 535545 59394 535611 59397
rect 536833 59394 536899 59397
rect 535545 59392 536899 59394
rect 535545 59336 535550 59392
rect 535606 59336 536838 59392
rect 536894 59336 536899 59392
rect 535545 59334 536899 59336
rect 536974 59394 537034 59606
rect 537864 59530 537924 60044
rect 538876 59530 538936 60044
rect 539888 59666 539948 60044
rect 540789 59666 540855 59669
rect 539888 59664 540855 59666
rect 539888 59608 540794 59664
rect 540850 59608 540855 59664
rect 539888 59606 540855 59608
rect 540992 59666 541052 60044
rect 541801 59666 541867 59669
rect 540992 59664 541867 59666
rect 540992 59608 541806 59664
rect 541862 59608 541867 59664
rect 540992 59606 541867 59608
rect 540789 59603 540855 59606
rect 541801 59603 541867 59606
rect 541065 59530 541131 59533
rect 537864 59470 538690 59530
rect 538876 59528 541131 59530
rect 538876 59472 541070 59528
rect 541126 59472 541131 59528
rect 538876 59470 541131 59472
rect 542004 59530 542064 60044
rect 543016 59666 543076 60044
rect 544028 59802 544088 60044
rect 544929 59802 544995 59805
rect 544028 59800 544995 59802
rect 544028 59744 544934 59800
rect 544990 59744 544995 59800
rect 544028 59742 544995 59744
rect 544929 59739 544995 59742
rect 545132 59666 545192 60044
rect 546144 59802 546204 60044
rect 546953 59802 547019 59805
rect 546144 59800 547019 59802
rect 546144 59744 546958 59800
rect 547014 59744 547019 59800
rect 546144 59742 547019 59744
rect 547156 59802 547216 60044
rect 547689 59802 547755 59805
rect 547156 59800 547755 59802
rect 547156 59744 547694 59800
rect 547750 59744 547755 59800
rect 547156 59742 547755 59744
rect 546953 59739 547019 59742
rect 547689 59739 547755 59742
rect 547873 59666 547939 59669
rect 543016 59606 544946 59666
rect 545132 59664 547939 59666
rect 545132 59608 547878 59664
rect 547934 59608 547939 59664
rect 545132 59606 547939 59608
rect 543825 59530 543891 59533
rect 542004 59528 543891 59530
rect 542004 59472 543830 59528
rect 543886 59472 543891 59528
rect 542004 59470 543891 59472
rect 544886 59530 544946 59606
rect 547873 59603 547939 59606
rect 545113 59530 545179 59533
rect 544886 59528 545179 59530
rect 544886 59472 545118 59528
rect 545174 59472 545179 59528
rect 544886 59470 545179 59472
rect 538305 59394 538371 59397
rect 536974 59392 538371 59394
rect 536974 59336 538310 59392
rect 538366 59336 538371 59392
rect 536974 59334 538371 59336
rect 538630 59394 538690 59470
rect 541065 59467 541131 59470
rect 543825 59467 543891 59470
rect 545113 59467 545179 59470
rect 546953 59530 547019 59533
rect 547965 59530 548031 59533
rect 546953 59528 548031 59530
rect 546953 59472 546958 59528
rect 547014 59472 547970 59528
rect 548026 59472 548031 59528
rect 546953 59470 548031 59472
rect 548168 59530 548228 60044
rect 549272 59666 549332 60044
rect 550081 59666 550147 59669
rect 549272 59664 550147 59666
rect 549272 59608 550086 59664
rect 550142 59608 550147 59664
rect 549272 59606 550147 59608
rect 550284 59666 550344 60044
rect 551296 59666 551356 60044
rect 552308 59802 552368 60044
rect 553412 59938 553472 60044
rect 554424 59938 554484 60044
rect 553412 59878 554330 59938
rect 554424 59878 555250 59938
rect 554270 59805 554330 59878
rect 552308 59742 554146 59802
rect 554270 59800 554379 59805
rect 554270 59744 554318 59800
rect 554374 59744 554379 59800
rect 554270 59742 554379 59744
rect 553393 59666 553459 59669
rect 550284 59606 551202 59666
rect 551296 59664 553459 59666
rect 551296 59608 553398 59664
rect 553454 59608 553459 59664
rect 551296 59606 553459 59608
rect 550081 59603 550147 59606
rect 550633 59530 550699 59533
rect 548168 59528 550699 59530
rect 548168 59472 550638 59528
rect 550694 59472 550699 59528
rect 548168 59470 550699 59472
rect 551142 59530 551202 59606
rect 553393 59603 553459 59606
rect 552289 59530 552355 59533
rect 551142 59528 552355 59530
rect 551142 59472 552294 59528
rect 552350 59472 552355 59528
rect 551142 59470 552355 59472
rect 546953 59467 547019 59470
rect 547965 59467 548031 59470
rect 550633 59467 550699 59470
rect 552289 59467 552355 59470
rect 539593 59394 539659 59397
rect 538630 59392 539659 59394
rect 538630 59336 539598 59392
rect 539654 59336 539659 59392
rect 538630 59334 539659 59336
rect 535545 59331 535611 59334
rect 536833 59331 536899 59334
rect 538305 59331 538371 59334
rect 539593 59331 539659 59334
rect 540789 59394 540855 59397
rect 542445 59394 542511 59397
rect 540789 59392 542511 59394
rect 540789 59336 540794 59392
rect 540850 59336 542450 59392
rect 542506 59336 542511 59392
rect 540789 59334 542511 59336
rect 540789 59331 540855 59334
rect 542445 59331 542511 59334
rect 544929 59394 544995 59397
rect 546493 59394 546559 59397
rect 544929 59392 546559 59394
rect 544929 59336 544934 59392
rect 544990 59336 546498 59392
rect 546554 59336 546559 59392
rect 544929 59334 546559 59336
rect 544929 59331 544995 59334
rect 546493 59331 546559 59334
rect 547689 59394 547755 59397
rect 549253 59394 549319 59397
rect 547689 59392 549319 59394
rect 547689 59336 547694 59392
rect 547750 59336 549258 59392
rect 549314 59336 549319 59392
rect 547689 59334 549319 59336
rect 547689 59331 547755 59334
rect 549253 59331 549319 59334
rect 550081 59394 550147 59397
rect 552105 59394 552171 59397
rect 550081 59392 552171 59394
rect 550081 59336 550086 59392
rect 550142 59336 552110 59392
rect 552166 59336 552171 59392
rect 550081 59334 552171 59336
rect 554086 59394 554146 59742
rect 554313 59739 554379 59742
rect 555190 59530 555250 59878
rect 555436 59666 555496 60044
rect 556448 59938 556508 60044
rect 556448 59878 556538 59938
rect 556478 59802 556538 59878
rect 556613 59802 556679 59805
rect 556478 59800 556679 59802
rect 556478 59744 556618 59800
rect 556674 59744 556679 59800
rect 556478 59742 556679 59744
rect 556613 59739 556679 59742
rect 555436 59606 557458 59666
rect 556521 59530 556587 59533
rect 555190 59528 556587 59530
rect 555190 59472 556526 59528
rect 556582 59472 556587 59528
rect 555190 59470 556587 59472
rect 556521 59467 556587 59470
rect 554773 59394 554839 59397
rect 554086 59392 554839 59394
rect 554086 59336 554778 59392
rect 554834 59336 554839 59392
rect 554086 59334 554839 59336
rect 550081 59331 550147 59334
rect 552105 59331 552171 59334
rect 554773 59331 554839 59334
rect 527173 59258 527239 59261
rect 526302 59256 527239 59258
rect 526302 59200 527178 59256
rect 527234 59200 527239 59256
rect 526302 59198 527239 59200
rect 557398 59258 557458 59606
rect 557552 59394 557612 60044
rect 558564 59530 558624 60044
rect 559576 59802 559636 60044
rect 560385 59802 560451 59805
rect 559576 59800 560451 59802
rect 559576 59744 560390 59800
rect 560446 59744 560451 59800
rect 559576 59742 560451 59744
rect 560385 59739 560451 59742
rect 560588 59666 560648 60044
rect 561489 59666 561555 59669
rect 560588 59664 561555 59666
rect 560588 59608 561494 59664
rect 561550 59608 561555 59664
rect 560588 59606 561555 59608
rect 561489 59603 561555 59606
rect 560569 59530 560635 59533
rect 558564 59528 560635 59530
rect 558564 59472 560574 59528
rect 560630 59472 560635 59528
rect 558564 59470 560635 59472
rect 560569 59467 560635 59470
rect 560385 59394 560451 59397
rect 557552 59392 560451 59394
rect 557552 59336 560390 59392
rect 560446 59336 560451 59392
rect 557552 59334 560451 59336
rect 561692 59394 561752 60044
rect 561857 59530 561923 59533
rect 562704 59530 562764 60044
rect 561857 59528 562764 59530
rect 561857 59472 561862 59528
rect 561918 59472 562764 59528
rect 561857 59470 562764 59472
rect 563716 59530 563776 60044
rect 564728 59666 564788 60044
rect 565832 59802 565892 60044
rect 566641 59802 566707 59805
rect 565832 59800 566707 59802
rect 565832 59744 566646 59800
rect 566702 59744 566707 59800
rect 565832 59742 566707 59744
rect 566641 59739 566707 59742
rect 564728 59606 566106 59666
rect 565813 59530 565879 59533
rect 563716 59528 565879 59530
rect 563716 59472 565818 59528
rect 565874 59472 565879 59528
rect 563716 59470 565879 59472
rect 561857 59467 561923 59470
rect 565813 59467 565879 59470
rect 564617 59394 564683 59397
rect 561692 59392 564683 59394
rect 561692 59336 564622 59392
rect 564678 59336 564683 59392
rect 561692 59334 564683 59336
rect 566046 59394 566106 59606
rect 566844 59530 566904 60044
rect 567856 59938 567916 60044
rect 567702 59878 567916 59938
rect 567009 59802 567075 59805
rect 567285 59802 567351 59805
rect 567009 59800 567351 59802
rect 567009 59744 567014 59800
rect 567070 59744 567290 59800
rect 567346 59744 567351 59800
rect 567009 59742 567351 59744
rect 567009 59739 567075 59742
rect 567285 59739 567351 59742
rect 567702 59666 567762 59878
rect 567702 59606 567916 59666
rect 566844 59470 567762 59530
rect 567193 59394 567259 59397
rect 566046 59392 567259 59394
rect 566046 59336 567198 59392
rect 567254 59336 567259 59392
rect 566046 59334 567259 59336
rect 560385 59331 560451 59334
rect 564617 59331 564683 59334
rect 567193 59331 567259 59334
rect 557625 59258 557691 59261
rect 557398 59256 557691 59258
rect 557398 59200 557630 59256
rect 557686 59200 557691 59256
rect 557398 59198 557691 59200
rect 567702 59258 567762 59470
rect 567856 59394 567916 59606
rect 568868 59530 568928 60044
rect 571333 59530 571399 59533
rect 568868 59528 571399 59530
rect 568868 59472 571338 59528
rect 571394 59472 571399 59528
rect 583520 59516 584960 59756
rect 568868 59470 571399 59472
rect 571333 59467 571399 59470
rect 569953 59394 570019 59397
rect 567856 59392 570019 59394
rect 567856 59336 569958 59392
rect 570014 59336 570019 59392
rect 567856 59334 570019 59336
rect 569953 59331 570019 59334
rect 568849 59258 568915 59261
rect 567702 59256 568915 59258
rect 567702 59200 568854 59256
rect 568910 59200 568915 59256
rect 567702 59198 568915 59200
rect 463233 59195 463299 59198
rect 469213 59195 469279 59198
rect 501045 59195 501111 59198
rect 503805 59195 503871 59198
rect 525793 59195 525859 59198
rect 527173 59195 527239 59198
rect 557625 59195 557691 59198
rect 568849 59195 568915 59198
rect 453481 59122 453547 59125
rect 450862 59120 453547 59122
rect 450862 59064 453486 59120
rect 453542 59064 453547 59120
rect 450862 59062 453547 59064
rect 174905 59059 174971 59062
rect 237005 59059 237071 59062
rect 278037 59059 278103 59062
rect 307385 59059 307451 59062
rect 440877 59059 440943 59062
rect 453481 59059 453547 59062
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
rect 19425 3362 19491 3365
rect 93117 3362 93183 3365
rect 19425 3360 93183 3362
rect 19425 3304 19430 3360
rect 19486 3304 93122 3360
rect 93178 3304 93183 3360
rect 19425 3302 93183 3304
rect 19425 3299 19491 3302
rect 93117 3299 93183 3302
rect 166809 3362 166875 3365
rect 583385 3362 583451 3365
rect 166809 3360 583451 3362
rect 166809 3304 166814 3360
rect 166870 3304 583390 3360
rect 583446 3304 583451 3360
rect 166809 3302 583451 3304
rect 166809 3299 166875 3302
rect 583385 3299 583451 3302
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 390032 60134 420618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 390032 63854 424338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 390032 67574 392058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 390032 74414 398898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 390032 78134 402618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 390032 81854 406338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 390032 85574 410058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 390032 92414 416898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 421174 96134 456618
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 390032 96134 420618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 424894 99854 460338
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 390032 99854 424338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 428614 103574 464058
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 392614 103574 428058
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 390032 103574 392058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 390032 110414 398898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 390032 114134 402618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 390032 117854 406338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 390032 121574 410058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 390032 128414 416898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 390032 132134 420618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 390032 135854 424338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 390032 139574 392058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 390032 146414 398898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 390032 150134 402618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 390032 153854 406338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 390032 157574 410058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 390032 164414 416898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 390032 168134 420618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 390032 171854 424338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 390032 175574 392058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 390032 182414 398898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 390032 186134 402618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 390032 189854 406338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 390032 193574 410058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 390032 200414 416898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 390032 204134 420618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 390032 207854 424338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 390032 211574 392058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 390032 218414 398898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 390032 222134 402618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 390032 225854 406338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 390032 229574 410058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 390032 236414 416898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 390032 240134 420618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 390032 243854 424338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 390032 247574 392058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 390032 254414 398898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 390032 258134 402618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 390032 261854 406338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 390032 265574 410058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 390032 272414 416898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 390032 276134 420618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 390032 279854 424338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 390032 283574 392058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 390032 290414 398898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 390032 294134 402618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 390032 297854 406338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 390032 301574 410058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 390032 308414 416898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 390032 312134 420618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 390032 315854 424338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 390032 319574 392058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 390032 326414 398898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 390032 330134 402618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 390032 333854 406338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 390032 337574 410058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 390032 344414 416898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 390032 348134 420618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 390032 351854 424338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 390032 355574 392058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 390032 362414 398898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 390032 366134 402618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 390032 369854 406338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 390032 373574 410058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 390032 380414 416898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 390032 384134 420618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 390032 387854 424338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 390032 391574 392058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 390032 398414 398898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 390032 402134 402618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 390032 405854 406338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 390032 409574 410058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 390032 416414 416898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 390032 420134 420618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 390032 423854 424338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 390032 427574 392058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 390032 434414 398898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 390032 438134 402618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 390032 441854 406338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 390032 445574 410058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 390032 452414 416898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 390032 456134 420618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 390032 459854 424338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 390032 463574 392058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 390032 470414 398898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 390032 474134 402618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 390032 477854 406338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 390032 481574 410058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 390032 488414 416898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 390032 492134 420618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 390032 495854 424338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 390032 499574 392058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 390032 506414 398898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 390032 510134 402618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 390032 513854 406338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 390032 517574 410058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 390032 524414 416898
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 390032 528134 420618
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 390032 531854 424338
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 390032 535574 392058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 390032 542414 398898
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 390032 546134 402618
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 390032 549854 406338
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 390032 553574 410058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 390032 560414 416898
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 390032 564134 420618
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 390032 567854 424338
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 390032 571574 392058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 58000
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 28894 63854 58000
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 32614 67574 58000
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 39454 74414 58000
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 43174 78134 58000
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 46894 81854 58000
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 50614 85574 58000
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 58000
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 58000
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 28894 99854 58000
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 32614 103574 58000
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 39454 110414 58000
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 43174 114134 58000
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 46894 117854 58000
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 50614 121574 58000
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 58000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 58000
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 28894 135854 58000
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 32614 139574 58000
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 39454 146414 58000
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 43174 150134 58000
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 46894 153854 58000
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 50614 157574 58000
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 57454 164414 58000
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 25174 168134 58000
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 28894 171854 58000
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 32614 175574 58000
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 39454 182414 58000
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 43174 186134 58000
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 46894 189854 58000
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 50614 193574 58000
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 57454 200414 58000
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 58000
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 28894 207854 58000
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 32614 211574 58000
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 39454 218414 58000
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 43174 222134 58000
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 46894 225854 58000
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 50614 229574 58000
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 57454 236414 58000
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 58000
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 28894 243854 58000
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 32614 247574 58000
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 39454 254414 58000
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 43174 258134 58000
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 46894 261854 58000
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 50614 265574 58000
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 57454 272414 58000
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 25174 276134 58000
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 28894 279854 58000
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 32614 283574 58000
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 39454 290414 58000
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 43174 294134 58000
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 46894 297854 58000
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 50614 301574 58000
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 57454 308414 58000
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 25174 312134 58000
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 28894 315854 58000
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 32614 319574 58000
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 39454 326414 58000
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 43174 330134 58000
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 46894 333854 58000
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 50614 337574 58000
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 57454 344414 58000
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 25174 348134 58000
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 28894 351854 58000
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 32614 355574 58000
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 39454 362414 58000
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 43174 366134 58000
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 46894 369854 58000
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 50614 373574 58000
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 57454 380414 58000
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 25174 384134 58000
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 28894 387854 58000
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 32614 391574 58000
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 39454 398414 58000
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 43174 402134 58000
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 46894 405854 58000
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 50614 409574 58000
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 57454 416414 58000
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 25174 420134 58000
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 28894 423854 58000
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 32614 427574 58000
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 39454 434414 58000
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 43174 438134 58000
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 46894 441854 58000
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 50614 445574 58000
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 57454 452414 58000
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 25174 456134 58000
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 28894 459854 58000
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 32614 463574 58000
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 39454 470414 58000
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 43174 474134 58000
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 46894 477854 58000
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 50614 481574 58000
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 57454 488414 58000
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 25174 492134 58000
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 28894 495854 58000
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 32614 499574 58000
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 39454 506414 58000
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 43174 510134 58000
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 46894 513854 58000
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 50614 517574 58000
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 57454 524414 58000
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 25174 528134 58000
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 28894 531854 58000
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 32614 535574 58000
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 39454 542414 58000
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 43174 546134 58000
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 46894 549854 58000
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 50614 553574 58000
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 57454 560414 58000
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 25174 564134 58000
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 28894 567854 58000
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 32614 571574 58000
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 58000 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 58000 388894
rect -6806 388574 58000 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 58000 388574
rect -6806 388306 58000 388338
rect 571956 388894 590730 388926
rect 571956 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 571956 388574 590730 388658
rect 571956 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 571956 388306 590730 388338
rect -4886 385174 58000 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 58000 385174
rect -4886 384854 58000 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 58000 384854
rect -4886 384586 58000 384618
rect 571956 385174 588810 385206
rect 571956 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 571956 384854 588810 384938
rect 571956 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 571956 384586 588810 384618
rect -2966 381454 58000 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 58000 381454
rect -2966 381134 58000 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 58000 381134
rect -2966 380866 58000 380898
rect 571956 381454 586890 381486
rect 571956 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 571956 381134 586890 381218
rect 571956 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 571956 380866 586890 380898
rect -8726 374614 58000 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 58000 374614
rect -8726 374294 58000 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 58000 374294
rect -8726 374026 58000 374058
rect 571956 374614 592650 374646
rect 571956 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect 571956 374294 592650 374378
rect 571956 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect 571956 374026 592650 374058
rect -6806 370894 58000 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 58000 370894
rect -6806 370574 58000 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 58000 370574
rect -6806 370306 58000 370338
rect 571956 370894 590730 370926
rect 571956 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect 571956 370574 590730 370658
rect 571956 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect 571956 370306 590730 370338
rect -4886 367174 58000 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 58000 367174
rect -4886 366854 58000 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 58000 366854
rect -4886 366586 58000 366618
rect 571956 367174 588810 367206
rect 571956 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect 571956 366854 588810 366938
rect 571956 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect 571956 366586 588810 366618
rect -2966 363454 58000 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 58000 363454
rect -2966 363134 58000 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 58000 363134
rect -2966 362866 58000 362898
rect 571956 363454 586890 363486
rect 571956 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect 571956 363134 586890 363218
rect 571956 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect 571956 362866 586890 362898
rect -8726 356614 58000 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 58000 356614
rect -8726 356294 58000 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 58000 356294
rect -8726 356026 58000 356058
rect 571956 356614 592650 356646
rect 571956 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 571956 356294 592650 356378
rect 571956 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 571956 356026 592650 356058
rect -6806 352894 58000 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 58000 352894
rect -6806 352574 58000 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 58000 352574
rect -6806 352306 58000 352338
rect 571956 352894 590730 352926
rect 571956 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 571956 352574 590730 352658
rect 571956 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 571956 352306 590730 352338
rect -4886 349174 58000 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 58000 349174
rect -4886 348854 58000 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 58000 348854
rect -4886 348586 58000 348618
rect 571956 349174 588810 349206
rect 571956 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 571956 348854 588810 348938
rect 571956 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 571956 348586 588810 348618
rect -2966 345454 58000 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 58000 345454
rect -2966 345134 58000 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 58000 345134
rect -2966 344866 58000 344898
rect 571956 345454 586890 345486
rect 571956 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 571956 345134 586890 345218
rect 571956 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 571956 344866 586890 344898
rect -8726 338614 58000 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 58000 338614
rect -8726 338294 58000 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 58000 338294
rect -8726 338026 58000 338058
rect 571956 338614 592650 338646
rect 571956 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect 571956 338294 592650 338378
rect 571956 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect 571956 338026 592650 338058
rect -6806 334894 58000 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 58000 334894
rect -6806 334574 58000 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 58000 334574
rect -6806 334306 58000 334338
rect 571956 334894 590730 334926
rect 571956 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect 571956 334574 590730 334658
rect 571956 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect 571956 334306 590730 334338
rect -4886 331174 58000 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 58000 331174
rect -4886 330854 58000 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 58000 330854
rect -4886 330586 58000 330618
rect 571956 331174 588810 331206
rect 571956 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect 571956 330854 588810 330938
rect 571956 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect 571956 330586 588810 330618
rect -2966 327454 58000 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 58000 327454
rect -2966 327134 58000 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 58000 327134
rect -2966 326866 58000 326898
rect 571956 327454 586890 327486
rect 571956 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect 571956 327134 586890 327218
rect 571956 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect 571956 326866 586890 326898
rect -8726 320614 58000 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 58000 320614
rect -8726 320294 58000 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 58000 320294
rect -8726 320026 58000 320058
rect 571956 320614 592650 320646
rect 571956 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 571956 320294 592650 320378
rect 571956 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 571956 320026 592650 320058
rect -6806 316894 58000 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 58000 316894
rect -6806 316574 58000 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 58000 316574
rect -6806 316306 58000 316338
rect 571956 316894 590730 316926
rect 571956 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 571956 316574 590730 316658
rect 571956 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 571956 316306 590730 316338
rect -4886 313174 58000 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 58000 313174
rect -4886 312854 58000 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 58000 312854
rect -4886 312586 58000 312618
rect 571956 313174 588810 313206
rect 571956 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 571956 312854 588810 312938
rect 571956 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 571956 312586 588810 312618
rect -2966 309454 58000 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 58000 309454
rect -2966 309134 58000 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 58000 309134
rect -2966 308866 58000 308898
rect 571956 309454 586890 309486
rect 571956 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 571956 309134 586890 309218
rect 571956 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 571956 308866 586890 308898
rect -8726 302614 58000 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 58000 302614
rect -8726 302294 58000 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 58000 302294
rect -8726 302026 58000 302058
rect 571956 302614 592650 302646
rect 571956 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect 571956 302294 592650 302378
rect 571956 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect 571956 302026 592650 302058
rect -6806 298894 58000 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 58000 298894
rect -6806 298574 58000 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 58000 298574
rect -6806 298306 58000 298338
rect 571956 298894 590730 298926
rect 571956 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect 571956 298574 590730 298658
rect 571956 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect 571956 298306 590730 298338
rect -4886 295174 58000 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 58000 295174
rect -4886 294854 58000 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 58000 294854
rect -4886 294586 58000 294618
rect 571956 295174 588810 295206
rect 571956 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect 571956 294854 588810 294938
rect 571956 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect 571956 294586 588810 294618
rect -2966 291454 58000 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 58000 291454
rect -2966 291134 58000 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 58000 291134
rect -2966 290866 58000 290898
rect 571956 291454 586890 291486
rect 571956 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect 571956 291134 586890 291218
rect 571956 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect 571956 290866 586890 290898
rect -8726 284614 58000 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 58000 284614
rect -8726 284294 58000 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 58000 284294
rect -8726 284026 58000 284058
rect 571956 284614 592650 284646
rect 571956 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 571956 284294 592650 284378
rect 571956 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 571956 284026 592650 284058
rect -6806 280894 58000 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 58000 280894
rect -6806 280574 58000 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 58000 280574
rect -6806 280306 58000 280338
rect 571956 280894 590730 280926
rect 571956 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 571956 280574 590730 280658
rect 571956 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 571956 280306 590730 280338
rect -4886 277174 58000 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 58000 277174
rect -4886 276854 58000 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 58000 276854
rect -4886 276586 58000 276618
rect 571956 277174 588810 277206
rect 571956 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 571956 276854 588810 276938
rect 571956 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 571956 276586 588810 276618
rect -2966 273454 58000 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 58000 273454
rect -2966 273134 58000 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 58000 273134
rect -2966 272866 58000 272898
rect 571956 273454 586890 273486
rect 571956 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 571956 273134 586890 273218
rect 571956 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 571956 272866 586890 272898
rect -8726 266614 58000 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 58000 266614
rect -8726 266294 58000 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 58000 266294
rect -8726 266026 58000 266058
rect 571956 266614 592650 266646
rect 571956 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect 571956 266294 592650 266378
rect 571956 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect 571956 266026 592650 266058
rect -6806 262894 58000 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 58000 262894
rect -6806 262574 58000 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 58000 262574
rect -6806 262306 58000 262338
rect 571956 262894 590730 262926
rect 571956 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect 571956 262574 590730 262658
rect 571956 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect 571956 262306 590730 262338
rect -4886 259174 58000 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 58000 259174
rect -4886 258854 58000 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 58000 258854
rect -4886 258586 58000 258618
rect 571956 259174 588810 259206
rect 571956 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect 571956 258854 588810 258938
rect 571956 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect 571956 258586 588810 258618
rect -2966 255454 58000 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 58000 255454
rect -2966 255134 58000 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 58000 255134
rect -2966 254866 58000 254898
rect 571956 255454 586890 255486
rect 571956 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect 571956 255134 586890 255218
rect 571956 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect 571956 254866 586890 254898
rect -8726 248614 58000 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 58000 248614
rect -8726 248294 58000 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 58000 248294
rect -8726 248026 58000 248058
rect 571956 248614 592650 248646
rect 571956 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 571956 248294 592650 248378
rect 571956 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 571956 248026 592650 248058
rect -6806 244894 58000 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 58000 244894
rect -6806 244574 58000 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 58000 244574
rect -6806 244306 58000 244338
rect 571956 244894 590730 244926
rect 571956 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 571956 244574 590730 244658
rect 571956 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 571956 244306 590730 244338
rect -4886 241174 58000 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 58000 241174
rect -4886 240854 58000 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 58000 240854
rect -4886 240586 58000 240618
rect 571956 241174 588810 241206
rect 571956 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 571956 240854 588810 240938
rect 571956 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 571956 240586 588810 240618
rect -2966 237454 58000 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 58000 237454
rect -2966 237134 58000 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 58000 237134
rect -2966 236866 58000 236898
rect 571956 237454 586890 237486
rect 571956 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 571956 237134 586890 237218
rect 571956 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 571956 236866 586890 236898
rect -8726 230614 58000 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 58000 230614
rect -8726 230294 58000 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 58000 230294
rect -8726 230026 58000 230058
rect 571956 230614 592650 230646
rect 571956 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect 571956 230294 592650 230378
rect 571956 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect 571956 230026 592650 230058
rect -6806 226894 58000 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 58000 226894
rect -6806 226574 58000 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 58000 226574
rect -6806 226306 58000 226338
rect 571956 226894 590730 226926
rect 571956 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect 571956 226574 590730 226658
rect 571956 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect 571956 226306 590730 226338
rect -4886 223174 58000 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 58000 223174
rect -4886 222854 58000 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 58000 222854
rect -4886 222586 58000 222618
rect 571956 223174 588810 223206
rect 571956 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect 571956 222854 588810 222938
rect 571956 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect 571956 222586 588810 222618
rect -2966 219454 58000 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 58000 219454
rect -2966 219134 58000 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 58000 219134
rect -2966 218866 58000 218898
rect 571956 219454 586890 219486
rect 571956 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect 571956 219134 586890 219218
rect 571956 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect 571956 218866 586890 218898
rect -8726 212614 58000 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 58000 212614
rect -8726 212294 58000 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 58000 212294
rect -8726 212026 58000 212058
rect 571956 212614 592650 212646
rect 571956 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 571956 212294 592650 212378
rect 571956 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 571956 212026 592650 212058
rect -6806 208894 58000 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 58000 208894
rect -6806 208574 58000 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 58000 208574
rect -6806 208306 58000 208338
rect 571956 208894 590730 208926
rect 571956 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 571956 208574 590730 208658
rect 571956 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 571956 208306 590730 208338
rect -4886 205174 58000 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 58000 205174
rect -4886 204854 58000 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 58000 204854
rect -4886 204586 58000 204618
rect 571956 205174 588810 205206
rect 571956 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 571956 204854 588810 204938
rect 571956 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 571956 204586 588810 204618
rect -2966 201454 58000 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 58000 201454
rect -2966 201134 58000 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 58000 201134
rect -2966 200866 58000 200898
rect 571956 201454 586890 201486
rect 571956 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 571956 201134 586890 201218
rect 571956 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 571956 200866 586890 200898
rect -8726 194614 58000 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 58000 194614
rect -8726 194294 58000 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 58000 194294
rect -8726 194026 58000 194058
rect 571956 194614 592650 194646
rect 571956 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect 571956 194294 592650 194378
rect 571956 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect 571956 194026 592650 194058
rect -6806 190894 58000 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 58000 190894
rect -6806 190574 58000 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 58000 190574
rect -6806 190306 58000 190338
rect 571956 190894 590730 190926
rect 571956 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect 571956 190574 590730 190658
rect 571956 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect 571956 190306 590730 190338
rect -4886 187174 58000 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 58000 187174
rect -4886 186854 58000 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 58000 186854
rect -4886 186586 58000 186618
rect 571956 187174 588810 187206
rect 571956 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect 571956 186854 588810 186938
rect 571956 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect 571956 186586 588810 186618
rect -2966 183454 58000 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 58000 183454
rect -2966 183134 58000 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 58000 183134
rect -2966 182866 58000 182898
rect 571956 183454 586890 183486
rect 571956 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect 571956 183134 586890 183218
rect 571956 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect 571956 182866 586890 182898
rect -8726 176614 58000 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 58000 176614
rect -8726 176294 58000 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 58000 176294
rect -8726 176026 58000 176058
rect 571956 176614 592650 176646
rect 571956 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 571956 176294 592650 176378
rect 571956 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 571956 176026 592650 176058
rect -6806 172894 58000 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 58000 172894
rect -6806 172574 58000 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 58000 172574
rect -6806 172306 58000 172338
rect 571956 172894 590730 172926
rect 571956 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 571956 172574 590730 172658
rect 571956 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 571956 172306 590730 172338
rect -4886 169174 58000 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 58000 169174
rect -4886 168854 58000 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 58000 168854
rect -4886 168586 58000 168618
rect 571956 169174 588810 169206
rect 571956 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 571956 168854 588810 168938
rect 571956 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 571956 168586 588810 168618
rect -2966 165454 58000 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 58000 165454
rect -2966 165134 58000 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 58000 165134
rect -2966 164866 58000 164898
rect 571956 165454 586890 165486
rect 571956 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 571956 165134 586890 165218
rect 571956 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 571956 164866 586890 164898
rect -8726 158614 58000 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 58000 158614
rect -8726 158294 58000 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 58000 158294
rect -8726 158026 58000 158058
rect 571956 158614 592650 158646
rect 571956 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect 571956 158294 592650 158378
rect 571956 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect 571956 158026 592650 158058
rect -6806 154894 58000 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 58000 154894
rect -6806 154574 58000 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 58000 154574
rect -6806 154306 58000 154338
rect 571956 154894 590730 154926
rect 571956 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect 571956 154574 590730 154658
rect 571956 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect 571956 154306 590730 154338
rect -4886 151174 58000 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 58000 151174
rect -4886 150854 58000 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 58000 150854
rect -4886 150586 58000 150618
rect 571956 151174 588810 151206
rect 571956 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect 571956 150854 588810 150938
rect 571956 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect 571956 150586 588810 150618
rect -2966 147454 58000 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 58000 147454
rect -2966 147134 58000 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 58000 147134
rect -2966 146866 58000 146898
rect 571956 147454 586890 147486
rect 571956 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect 571956 147134 586890 147218
rect 571956 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect 571956 146866 586890 146898
rect -8726 140614 58000 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 58000 140614
rect -8726 140294 58000 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 58000 140294
rect -8726 140026 58000 140058
rect 571956 140614 592650 140646
rect 571956 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 571956 140294 592650 140378
rect 571956 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 571956 140026 592650 140058
rect -6806 136894 58000 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 58000 136894
rect -6806 136574 58000 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 58000 136574
rect -6806 136306 58000 136338
rect 571956 136894 590730 136926
rect 571956 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 571956 136574 590730 136658
rect 571956 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 571956 136306 590730 136338
rect -4886 133174 58000 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 58000 133174
rect -4886 132854 58000 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 58000 132854
rect -4886 132586 58000 132618
rect 571956 133174 588810 133206
rect 571956 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 571956 132854 588810 132938
rect 571956 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 571956 132586 588810 132618
rect -2966 129454 58000 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 58000 129454
rect -2966 129134 58000 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 58000 129134
rect -2966 128866 58000 128898
rect 571956 129454 586890 129486
rect 571956 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 571956 129134 586890 129218
rect 571956 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 571956 128866 586890 128898
rect -8726 122614 58000 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 58000 122614
rect -8726 122294 58000 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 58000 122294
rect -8726 122026 58000 122058
rect 571956 122614 592650 122646
rect 571956 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect 571956 122294 592650 122378
rect 571956 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect 571956 122026 592650 122058
rect -6806 118894 58000 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 58000 118894
rect -6806 118574 58000 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 58000 118574
rect -6806 118306 58000 118338
rect 571956 118894 590730 118926
rect 571956 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect 571956 118574 590730 118658
rect 571956 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect 571956 118306 590730 118338
rect -4886 115174 58000 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 58000 115174
rect -4886 114854 58000 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 58000 114854
rect -4886 114586 58000 114618
rect 571956 115174 588810 115206
rect 571956 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect 571956 114854 588810 114938
rect 571956 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect 571956 114586 588810 114618
rect -2966 111454 58000 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 58000 111454
rect -2966 111134 58000 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 58000 111134
rect -2966 110866 58000 110898
rect 571956 111454 586890 111486
rect 571956 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect 571956 111134 586890 111218
rect 571956 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect 571956 110866 586890 110898
rect -8726 104614 58000 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 58000 104614
rect -8726 104294 58000 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 58000 104294
rect -8726 104026 58000 104058
rect 571956 104614 592650 104646
rect 571956 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 571956 104294 592650 104378
rect 571956 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 571956 104026 592650 104058
rect -6806 100894 58000 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 58000 100894
rect -6806 100574 58000 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 58000 100574
rect -6806 100306 58000 100338
rect 571956 100894 590730 100926
rect 571956 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 571956 100574 590730 100658
rect 571956 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 571956 100306 590730 100338
rect -4886 97174 58000 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 58000 97174
rect -4886 96854 58000 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 58000 96854
rect -4886 96586 58000 96618
rect 571956 97174 588810 97206
rect 571956 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 571956 96854 588810 96938
rect 571956 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 571956 96586 588810 96618
rect -2966 93454 58000 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 58000 93454
rect -2966 93134 58000 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 58000 93134
rect -2966 92866 58000 92898
rect 571956 93454 586890 93486
rect 571956 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 571956 93134 586890 93218
rect 571956 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 571956 92866 586890 92898
rect -8726 86614 58000 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 58000 86614
rect -8726 86294 58000 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 58000 86294
rect -8726 86026 58000 86058
rect 571956 86614 592650 86646
rect 571956 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect 571956 86294 592650 86378
rect 571956 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect 571956 86026 592650 86058
rect -6806 82894 58000 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 58000 82894
rect -6806 82574 58000 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 58000 82574
rect -6806 82306 58000 82338
rect 571956 82894 590730 82926
rect 571956 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect 571956 82574 590730 82658
rect 571956 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect 571956 82306 590730 82338
rect -4886 79174 58000 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 58000 79174
rect -4886 78854 58000 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 58000 78854
rect -4886 78586 58000 78618
rect 571956 79174 588810 79206
rect 571956 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect 571956 78854 588810 78938
rect 571956 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect 571956 78586 588810 78618
rect -2966 75454 58000 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 58000 75454
rect -2966 75134 58000 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 58000 75134
rect -2966 74866 58000 74898
rect 571956 75454 586890 75486
rect 571956 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect 571956 75134 586890 75218
rect 571956 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect 571956 74866 586890 74898
rect -8726 68614 58000 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 58000 68614
rect -8726 68294 58000 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 58000 68294
rect -8726 68026 58000 68058
rect 571956 68614 592650 68646
rect 571956 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 571956 68294 592650 68378
rect 571956 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 571956 68026 592650 68058
rect -6806 64894 58000 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 58000 64894
rect -6806 64574 58000 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 58000 64574
rect -6806 64306 58000 64338
rect 571956 64894 590730 64926
rect 571956 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 571956 64574 590730 64658
rect 571956 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 571956 64306 590730 64338
rect -4886 61174 58000 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 58000 61174
rect -4886 60854 58000 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 58000 60854
rect -4886 60586 58000 60618
rect 571956 61174 588810 61206
rect 571956 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 571956 60854 588810 60938
rect 571956 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 571956 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use azadi_soc_top_caravel  mprj
timestamp 0
transform 1 0 60000 0 1 60000
box 0 0 509956 328032
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 58000 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s 571956 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 58000 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s 571956 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 58000 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s 571956 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 58000 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s 571956 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 58000 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s 571956 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 58000 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s 571956 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 58000 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s 571956 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 58000 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s 571956 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 58000 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s 571956 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 390032 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 390032 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 390032 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 390032 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 390032 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 390032 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 390032 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 390032 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 390032 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 390032 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 390032 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 390032 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 390032 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 390032 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 58000 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s 571956 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 58000 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s 571956 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 58000 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s 571956 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 58000 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s 571956 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 58000 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s 571956 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 58000 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s 571956 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 58000 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s 571956 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 58000 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s 571956 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 58000 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s 571956 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 390032 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 390032 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 390032 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 390032 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 390032 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 390032 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 390032 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 390032 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 390032 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 390032 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 390032 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 390032 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 390032 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 390032 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 58000 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s 571956 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 58000 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s 571956 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 58000 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s 571956 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 58000 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s 571956 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 58000 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s 571956 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 58000 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s 571956 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 58000 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s 571956 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 58000 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s 571956 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 58000 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s 571956 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 390032 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 390032 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 390032 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 390032 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 390032 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 390032 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 390032 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 390032 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 390032 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 390032 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 390032 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 390032 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 390032 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 390032 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 58000 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s 571956 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 58000 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s 571956 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 58000 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s 571956 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 58000 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s 571956 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 58000 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s 571956 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 58000 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s 571956 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 58000 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s 571956 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 58000 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s 571956 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 58000 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s 571956 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 390032 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 390032 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 390032 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 390032 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 390032 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 390032 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 390032 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 390032 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 390032 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 390032 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 390032 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 390032 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 390032 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 390032 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 58000 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 571956 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 58000 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 571956 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 58000 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 571956 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 58000 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 571956 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 58000 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 571956 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 58000 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 571956 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 58000 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 571956 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 58000 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 571956 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 58000 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 571956 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 58000 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 571956 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 390032 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 390032 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 390032 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 390032 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 390032 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 390032 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 390032 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 390032 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 390032 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 390032 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 390032 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 390032 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 390032 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 390032 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 390032 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 58000 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 571956 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 58000 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 571956 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 58000 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 571956 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 58000 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 571956 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 58000 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 571956 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 58000 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 571956 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 58000 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 571956 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 58000 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 571956 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 58000 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 571956 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 390032 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 390032 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 390032 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 390032 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 390032 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 390032 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 390032 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 390032 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 390032 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 390032 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 390032 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 390032 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 390032 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 390032 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 390032 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 58000 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 571956 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 58000 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 571956 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 58000 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 571956 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 58000 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 571956 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 58000 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 571956 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 58000 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 571956 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 58000 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 571956 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 58000 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 571956 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 58000 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 571956 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 390032 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 390032 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 390032 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 390032 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 390032 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 390032 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 390032 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 390032 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 390032 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 390032 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 390032 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 390032 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 390032 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 390032 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 58000 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 571956 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 58000 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 571956 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 58000 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 571956 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 58000 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 571956 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 58000 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 571956 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 58000 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 571956 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 58000 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 571956 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 58000 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 571956 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 58000 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 571956 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 58000 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 571956 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 390032 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 390032 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 390032 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 390032 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 390032 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 390032 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 390032 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 390032 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 390032 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 390032 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 390032 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 390032 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 390032 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 390032 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 390032 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
