##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Mon Jun  6 00:25:34 2022
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO azadi_soc_top_caravel
  CLASS BLOCK ;
  SIZE 2549.780000 BY 1640.160000 ;
  FOREIGN azadi_soc_top_caravel 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1926 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 538.280000 0.000000 538.580000 0.800000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.608 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 10.324 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 49 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1637.970000 0.800000 1638.270000 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 5.600000 0.000000 5.900000 0.800000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 362.100000 0.000000 362.400000 0.800000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.920000 0.000000 2.220000 0.800000 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 10.660000 0.000000 10.960000 0.800000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 15.720000 0.000000 16.020000 0.800000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 20.780000 0.000000 21.080000 0.800000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 26.300000 0.000000 26.600000 0.800000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.960000 0.000000 197.260000 0.800000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 202.020000 0.000000 202.320000 0.800000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 207.080000 0.000000 207.380000 0.800000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 212.140000 0.000000 212.440000 0.800000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 217.660000 0.000000 217.960000 0.800000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 222.720000 0.000000 223.020000 0.800000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 227.780000 0.000000 228.080000 0.800000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 232.840000 0.000000 233.140000 0.800000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 238.360000 0.000000 238.660000 0.800000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 243.420000 0.000000 243.720000 0.800000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 248.480000 0.000000 248.780000 0.800000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 253.540000 0.000000 253.840000 0.800000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 259.060000 0.000000 259.360000 0.800000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 264.120000 0.000000 264.420000 0.800000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 269.180000 0.000000 269.480000 0.800000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 274.240000 0.000000 274.540000 0.800000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 279.760000 0.000000 280.060000 0.800000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 284.820000 0.000000 285.120000 0.800000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 289.880000 0.000000 290.180000 0.800000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 294.940000 0.000000 295.240000 0.800000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 300.460000 0.000000 300.760000 0.800000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 305.520000 0.000000 305.820000 0.800000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 310.580000 0.000000 310.880000 0.800000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 315.640000 0.000000 315.940000 0.800000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 320.700000 0.000000 321.000000 0.800000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 326.220000 0.000000 326.520000 0.800000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 331.280000 0.000000 331.580000 0.800000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 336.340000 0.000000 336.640000 0.800000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 341.400000 0.000000 341.700000 0.800000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.920000 0.000000 347.220000 0.800000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 351.980000 0.000000 352.280000 0.800000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 357.040000 0.000000 357.340000 0.800000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 367.620000 0.000000 367.920000 0.800000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 372.680000 0.000000 372.980000 0.800000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 377.740000 0.000000 378.040000 0.800000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 382.800000 0.000000 383.100000 0.800000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 388.320000 0.000000 388.620000 0.800000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.380000 0.000000 393.680000 0.800000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 398.440000 0.000000 398.740000 0.800000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 403.500000 0.000000 403.800000 0.800000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 409.020000 0.000000 409.320000 0.800000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 414.080000 0.000000 414.380000 0.800000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 419.140000 0.000000 419.440000 0.800000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 424.200000 0.000000 424.500000 0.800000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 429.720000 0.000000 430.020000 0.800000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 434.780000 0.000000 435.080000 0.800000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 439.840000 0.000000 440.140000 0.800000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 444.900000 0.000000 445.200000 0.800000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 450.420000 0.000000 450.720000 0.800000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 455.480000 0.000000 455.780000 0.800000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 460.540000 0.000000 460.840000 0.800000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 465.600000 0.000000 465.900000 0.800000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 470.660000 0.000000 470.960000 0.800000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.180000 0.000000 476.480000 0.800000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 481.240000 0.000000 481.540000 0.800000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 486.300000 0.000000 486.600000 0.800000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 491.360000 0.000000 491.660000 0.800000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.880000 0.000000 497.180000 0.800000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 501.940000 0.000000 502.240000 0.800000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 507.000000 0.000000 507.300000 0.800000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 512.060000 0.000000 512.360000 0.800000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 517.580000 0.000000 517.880000 0.800000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 522.640000 0.000000 522.940000 0.800000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 527.700000 0.000000 528.000000 0.800000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.526 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.51 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 532.760000 0.000000 533.060000 0.800000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.549 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 31.360000 0.000000 31.660000 0.800000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.53 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 36.420000 0.000000 36.720000 0.800000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.7 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 41.480000 0.000000 41.780000 0.800000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.7 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 47.000000 0.000000 47.300000 0.800000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.53 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 52.060000 0.000000 52.360000 0.800000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.53 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 57.120000 0.000000 57.420000 0.800000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.53 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 62.180000 0.000000 62.480000 0.800000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.53 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 67.700000 0.000000 68.000000 0.800000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.53 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 72.760000 0.000000 73.060000 0.800000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.53 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 77.820000 0.000000 78.120000 0.800000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.53 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 82.880000 0.000000 83.180000 0.800000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.53 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 88.400000 0.000000 88.700000 0.800000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.53 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 93.460000 0.000000 93.760000 0.800000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.53 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 98.520000 0.000000 98.820000 0.800000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.53 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 103.580000 0.000000 103.880000 0.800000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.53 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 109.100000 0.000000 109.400000 0.800000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.53 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 114.160000 0.000000 114.460000 0.800000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.53 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 119.220000 0.000000 119.520000 0.800000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.7 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 124.280000 0.000000 124.580000 0.800000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.7 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 129.800000 0.000000 130.100000 0.800000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.53 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 134.860000 0.000000 135.160000 0.800000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.53 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 139.920000 0.000000 140.220000 0.800000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.53 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 144.980000 0.000000 145.280000 0.800000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.53 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 150.040000 0.000000 150.340000 0.800000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.53 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 155.560000 0.000000 155.860000 0.800000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.53 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 160.620000 0.000000 160.920000 0.800000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.53 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 165.680000 0.000000 165.980000 0.800000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.53 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 170.740000 0.000000 171.040000 0.800000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.53 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 176.260000 0.000000 176.560000 0.800000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.53 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 181.320000 0.000000 181.620000 0.800000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.53 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 186.380000 0.000000 186.680000 0.800000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.549 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 191.440000 0.000000 191.740000 0.800000 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1887.920000 0.000000 1888.220000 0.800000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1892.980000 0.000000 1893.280000 0.800000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1898.040000 0.000000 1898.340000 0.800000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1903.100000 0.000000 1903.400000 0.800000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1908.620000 0.000000 1908.920000 0.800000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1913.680000 0.000000 1913.980000 0.800000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1918.740000 0.000000 1919.040000 0.800000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1923.800000 0.000000 1924.100000 0.800000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1929.320000 0.000000 1929.620000 0.800000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1934.380000 0.000000 1934.680000 0.800000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1939.440000 0.000000 1939.740000 0.800000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1944.500000 0.000000 1944.800000 0.800000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1949.560000 0.000000 1949.860000 0.800000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1955.080000 0.000000 1955.380000 0.800000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1960.140000 0.000000 1960.440000 0.800000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1965.200000 0.000000 1965.500000 0.800000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1970.260000 0.000000 1970.560000 0.800000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1975.780000 0.000000 1976.080000 0.800000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1980.840000 0.000000 1981.140000 0.800000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1985.900000 0.000000 1986.200000 0.800000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1990.960000 0.000000 1991.260000 0.800000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.480000 0.000000 1996.780000 0.800000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2001.540000 0.000000 2001.840000 0.800000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2006.600000 0.000000 2006.900000 0.800000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2011.660000 0.000000 2011.960000 0.800000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2017.180000 0.000000 2017.480000 0.800000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2022.240000 0.000000 2022.540000 0.800000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2027.300000 0.000000 2027.600000 0.800000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2032.360000 0.000000 2032.660000 0.800000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2037.880000 0.000000 2038.180000 0.800000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2042.940000 0.000000 2043.240000 0.800000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2048.000000 0.000000 2048.300000 0.800000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2053.060000 0.000000 2053.360000 0.800000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2058.580000 0.000000 2058.880000 0.800000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2063.640000 0.000000 2063.940000 0.800000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2068.700000 0.000000 2069.000000 0.800000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2073.760000 0.000000 2074.060000 0.800000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2079.280000 0.000000 2079.580000 0.800000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2084.340000 0.000000 2084.640000 0.800000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2089.400000 0.000000 2089.700000 0.800000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2094.460000 0.000000 2094.760000 0.800000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2099.520000 0.000000 2099.820000 0.800000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2105.040000 0.000000 2105.340000 0.800000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2110.100000 0.000000 2110.400000 0.800000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2115.160000 0.000000 2115.460000 0.800000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2120.220000 0.000000 2120.520000 0.800000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2125.740000 0.000000 2126.040000 0.800000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2130.800000 0.000000 2131.100000 0.800000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2135.860000 0.000000 2136.160000 0.800000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2140.920000 0.000000 2141.220000 0.800000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.440000 0.000000 2146.740000 0.800000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2151.500000 0.000000 2151.800000 0.800000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2156.560000 0.000000 2156.860000 0.800000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2161.620000 0.000000 2161.920000 0.800000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2167.140000 0.000000 2167.440000 0.800000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2172.200000 0.000000 2172.500000 0.800000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2177.260000 0.000000 2177.560000 0.800000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2182.320000 0.000000 2182.620000 0.800000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2187.840000 0.000000 2188.140000 0.800000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2192.900000 0.000000 2193.200000 0.800000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2197.960000 0.000000 2198.260000 0.800000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2203.020000 0.000000 2203.320000 0.800000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2208.540000 0.000000 2208.840000 0.800000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2213.600000 0.000000 2213.900000 0.800000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2218.660000 0.000000 2218.960000 0.800000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2223.720000 0.000000 2224.020000 0.800000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2229.240000 0.000000 2229.540000 0.800000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2234.300000 0.000000 2234.600000 0.800000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2239.360000 0.000000 2239.660000 0.800000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2244.420000 0.000000 2244.720000 0.800000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2249.480000 0.000000 2249.780000 0.800000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2255.000000 0.000000 2255.300000 0.800000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2260.060000 0.000000 2260.360000 0.800000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2265.120000 0.000000 2265.420000 0.800000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2270.180000 0.000000 2270.480000 0.800000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2275.700000 0.000000 2276.000000 0.800000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2280.760000 0.000000 2281.060000 0.800000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2285.820000 0.000000 2286.120000 0.800000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2290.880000 0.000000 2291.180000 0.800000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.400000 0.000000 2296.700000 0.800000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2301.460000 0.000000 2301.760000 0.800000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2306.520000 0.000000 2306.820000 0.800000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2311.580000 0.000000 2311.880000 0.800000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2317.100000 0.000000 2317.400000 0.800000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2322.160000 0.000000 2322.460000 0.800000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2327.220000 0.000000 2327.520000 0.800000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2332.280000 0.000000 2332.580000 0.800000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2337.800000 0.000000 2338.100000 0.800000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2342.860000 0.000000 2343.160000 0.800000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2347.920000 0.000000 2348.220000 0.800000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2352.980000 0.000000 2353.280000 0.800000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2358.500000 0.000000 2358.800000 0.800000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2363.560000 0.000000 2363.860000 0.800000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.620000 0.000000 2368.920000 0.800000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2373.680000 0.000000 2373.980000 0.800000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2379.200000 0.000000 2379.500000 0.800000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2384.260000 0.000000 2384.560000 0.800000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2389.320000 0.000000 2389.620000 0.800000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2394.380000 0.000000 2394.680000 0.800000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.440000 0.000000 2399.740000 0.800000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2404.960000 0.000000 2405.260000 0.800000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2410.020000 0.000000 2410.320000 0.800000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2415.080000 0.000000 2415.380000 0.800000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2420.140000 0.000000 2420.440000 0.800000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2425.660000 0.000000 2425.960000 0.800000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2430.720000 0.000000 2431.020000 0.800000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2435.780000 0.000000 2436.080000 0.800000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2440.840000 0.000000 2441.140000 0.800000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2446.360000 0.000000 2446.660000 0.800000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2451.420000 0.000000 2451.720000 0.800000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2456.480000 0.000000 2456.780000 0.800000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2461.540000 0.000000 2461.840000 0.800000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 29.5998 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 158.336 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2467.060000 0.000000 2467.360000 0.800000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 33.1878 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 177.472 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2472.120000 0.000000 2472.420000 0.800000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.6288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 131.824 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2477.180000 0.000000 2477.480000 0.800000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.1808 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 134.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2482.240000 0.000000 2482.540000 0.800000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 29.8728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 159.792 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2487.760000 0.000000 2488.060000 0.800000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.4848 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.056 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2492.820000 0.000000 2493.120000 0.800000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.9728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 122.992 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2497.880000 0.000000 2498.180000 0.800000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 26.8368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 143.6 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2502.940000 0.000000 2503.240000 0.800000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 55.9728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 298.992 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2508.460000 0.000000 2508.760000 0.800000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.3668 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 167.76 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2513.520000 0.000000 2513.820000 0.800000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 34.3578 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 183.712 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2518.580000 0.000000 2518.880000 0.800000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.8358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 132.928 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2523.640000 0.000000 2523.940000 0.800000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.1408 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 107.888 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2529.160000 0.000000 2529.460000 0.800000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 99.4998 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 531.136 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2534.220000 0.000000 2534.520000 0.800000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 53.4048 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 285.296 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2539.280000 0.000000 2539.580000 0.800000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.9688 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.304 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2544.340000 0.000000 2544.640000 0.800000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.752 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.936 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 504.05 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2690.65 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1225.980000 0.000000 1226.280000 0.800000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1231.040000 0.000000 1231.340000 0.800000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1236.100000 0.000000 1236.400000 0.800000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1241.160000 0.000000 1241.460000 0.800000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1246.680000 0.000000 1246.980000 0.800000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1251.740000 0.000000 1252.040000 0.800000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1256.800000 0.000000 1257.100000 0.800000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1261.860000 0.000000 1262.160000 0.800000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1267.380000 0.000000 1267.680000 0.800000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1272.440000 0.000000 1272.740000 0.800000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1277.500000 0.000000 1277.800000 0.800000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1282.560000 0.000000 1282.860000 0.800000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1288.080000 0.000000 1288.380000 0.800000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1293.140000 0.000000 1293.440000 0.800000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1298.200000 0.000000 1298.500000 0.800000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.888 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2690.46 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1303.260000 0.000000 1303.560000 0.800000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.888 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2690.46 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1308.780000 0.000000 1309.080000 0.800000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1313.840000 0.000000 1314.140000 0.800000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1318.900000 0.000000 1319.200000 0.800000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1323.960000 0.000000 1324.260000 0.800000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1329.480000 0.000000 1329.780000 0.800000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1334.540000 0.000000 1334.840000 0.800000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1339.600000 0.000000 1339.900000 0.800000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1344.660000 0.000000 1344.960000 0.800000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1350.180000 0.000000 1350.480000 0.800000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1355.240000 0.000000 1355.540000 0.800000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1360.300000 0.000000 1360.600000 0.800000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1365.360000 0.000000 1365.660000 0.800000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.888 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2690.46 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1370.420000 0.000000 1370.720000 0.800000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.888 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2690.46 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1375.940000 0.000000 1376.240000 0.800000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1381.000000 0.000000 1381.300000 0.800000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1386.060000 0.000000 1386.360000 0.800000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1391.120000 0.000000 1391.420000 0.800000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1396.640000 0.000000 1396.940000 0.800000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1401.700000 0.000000 1402.000000 0.800000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1406.760000 0.000000 1407.060000 0.800000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1411.820000 0.000000 1412.120000 0.800000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1417.340000 0.000000 1417.640000 0.800000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1422.400000 0.000000 1422.700000 0.800000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1427.460000 0.000000 1427.760000 0.800000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1432.520000 0.000000 1432.820000 0.800000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1438.040000 0.000000 1438.340000 0.800000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1443.100000 0.000000 1443.400000 0.800000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1448.160000 0.000000 1448.460000 0.800000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.888 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2690.46 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1453.220000 0.000000 1453.520000 0.800000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.888 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2690.46 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1458.740000 0.000000 1459.040000 0.800000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1463.800000 0.000000 1464.100000 0.800000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1468.860000 0.000000 1469.160000 0.800000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1473.920000 0.000000 1474.220000 0.800000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1479.440000 0.000000 1479.740000 0.800000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1484.500000 0.000000 1484.800000 0.800000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1489.560000 0.000000 1489.860000 0.800000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1494.620000 0.000000 1494.920000 0.800000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1499.680000 0.000000 1499.980000 0.800000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1505.200000 0.000000 1505.500000 0.800000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1510.260000 0.000000 1510.560000 0.800000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1515.320000 0.000000 1515.620000 0.800000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1520.380000 0.000000 1520.680000 0.800000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1525.900000 0.000000 1526.200000 0.800000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1530.960000 0.000000 1531.260000 0.800000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.888 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2690.46 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1536.020000 0.000000 1536.320000 0.800000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.888 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2690.46 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1541.080000 0.000000 1541.380000 0.800000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1546.600000 0.000000 1546.900000 0.800000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1551.660000 0.000000 1551.960000 0.800000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1556.720000 0.000000 1557.020000 0.800000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1561.780000 0.000000 1562.080000 0.800000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1567.300000 0.000000 1567.600000 0.800000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1572.360000 0.000000 1572.660000 0.800000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1577.420000 0.000000 1577.720000 0.800000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1582.480000 0.000000 1582.780000 0.800000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1588.000000 0.000000 1588.300000 0.800000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1593.060000 0.000000 1593.360000 0.800000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 503.971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2689.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1598.120000 0.000000 1598.420000 0.800000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 124.752 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 665.936 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 513.534 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2730.82 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1603.180000 0.000000 1603.480000 0.800000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.139 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.416 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 446.854 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2377.69 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 464.91 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2479.51 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1608.700000 0.000000 1609.000000 0.800000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.192 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2334.23 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2436.06 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1613.760000 0.000000 1614.060000 0.800000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.192 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2334.23 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2436.06 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1618.820000 0.000000 1619.120000 0.800000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.192 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2334.23 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2436.06 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1623.880000 0.000000 1624.180000 0.800000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1629.400000 0.000000 1629.700000 0.800000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1634.460000 0.000000 1634.760000 0.800000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1639.520000 0.000000 1639.820000 0.800000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1644.580000 0.000000 1644.880000 0.800000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1649.640000 0.000000 1649.940000 0.800000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1655.160000 0.000000 1655.460000 0.800000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1660.220000 0.000000 1660.520000 0.800000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1665.280000 0.000000 1665.580000 0.800000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1670.340000 0.000000 1670.640000 0.800000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1675.860000 0.000000 1676.160000 0.800000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1680.920000 0.000000 1681.220000 0.800000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1685.980000 0.000000 1686.280000 0.800000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1691.040000 0.000000 1691.340000 0.800000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1696.560000 0.000000 1696.860000 0.800000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.192 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2334.23 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2436.06 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1701.620000 0.000000 1701.920000 0.800000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.192 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2334.23 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2436.06 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1706.680000 0.000000 1706.980000 0.800000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.192 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2334.23 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2436.06 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1711.740000 0.000000 1712.040000 0.800000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.192 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2334.23 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2436.06 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1717.260000 0.000000 1717.560000 0.800000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1722.320000 0.000000 1722.620000 0.800000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1727.380000 0.000000 1727.680000 0.800000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1732.440000 0.000000 1732.740000 0.800000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1737.960000 0.000000 1738.260000 0.800000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1743.020000 0.000000 1743.320000 0.800000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1748.080000 0.000000 1748.380000 0.800000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1753.140000 0.000000 1753.440000 0.800000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1758.660000 0.000000 1758.960000 0.800000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1763.720000 0.000000 1764.020000 0.800000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1768.780000 0.000000 1769.080000 0.800000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1773.840000 0.000000 1774.140000 0.800000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1779.360000 0.000000 1779.660000 0.800000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.192 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2334.23 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2436.06 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1784.420000 0.000000 1784.720000 0.800000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.192 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2334.23 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2436.06 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1789.480000 0.000000 1789.780000 0.800000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1794.540000 0.000000 1794.840000 0.800000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.192 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2334.23 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2436.06 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1799.600000 0.000000 1799.900000 0.800000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.192 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2334.23 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2436.06 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1805.120000 0.000000 1805.420000 0.800000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1810.180000 0.000000 1810.480000 0.800000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1815.240000 0.000000 1815.540000 0.800000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1820.300000 0.000000 1820.600000 0.800000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1825.820000 0.000000 1826.120000 0.800000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1830.880000 0.000000 1831.180000 0.800000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1835.940000 0.000000 1836.240000 0.800000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1841.000000 0.000000 1841.300000 0.800000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1846.520000 0.000000 1846.820000 0.800000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1851.580000 0.000000 1851.880000 0.800000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1856.640000 0.000000 1856.940000 0.800000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1861.700000 0.000000 1862.000000 0.800000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.192 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2334.23 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2436.06 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1867.220000 0.000000 1867.520000 0.800000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.192 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2334.23 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2436.06 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1872.280000 0.000000 1872.580000 0.800000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2333.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.16 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2435.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1877.340000 0.000000 1877.640000 0.800000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.1225 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 497.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 437.195 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2334.46 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 455.251 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2436.28 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.187793 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1882.400000 0.000000 1882.700000 0.800000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 564.040000 0.000000 564.340000 0.800000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 569.100000 0.000000 569.400000 0.800000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.160000 0.000000 574.460000 0.800000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 579.680000 0.000000 579.980000 0.800000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 584.740000 0.000000 585.040000 0.800000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 589.800000 0.000000 590.100000 0.800000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 594.860000 0.000000 595.160000 0.800000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 600.380000 0.000000 600.680000 0.800000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 605.440000 0.000000 605.740000 0.800000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 610.500000 0.000000 610.800000 0.800000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 615.560000 0.000000 615.860000 0.800000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 620.620000 0.000000 620.920000 0.800000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 626.140000 0.000000 626.440000 0.800000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 631.200000 0.000000 631.500000 0.800000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 636.260000 0.000000 636.560000 0.800000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 641.320000 0.000000 641.620000 0.800000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.840000 0.000000 647.140000 0.800000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 651.900000 0.000000 652.200000 0.800000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 656.960000 0.000000 657.260000 0.800000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 662.020000 0.000000 662.320000 0.800000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 667.540000 0.000000 667.840000 0.800000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 672.600000 0.000000 672.900000 0.800000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 677.660000 0.000000 677.960000 0.800000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 682.720000 0.000000 683.020000 0.800000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 688.240000 0.000000 688.540000 0.800000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 693.300000 0.000000 693.600000 0.800000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 698.360000 0.000000 698.660000 0.800000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 703.420000 0.000000 703.720000 0.800000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 708.940000 0.000000 709.240000 0.800000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 714.000000 0.000000 714.300000 0.800000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 719.060000 0.000000 719.360000 0.800000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 724.120000 0.000000 724.420000 0.800000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 729.640000 0.000000 729.940000 0.800000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 734.700000 0.000000 735.000000 0.800000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 739.760000 0.000000 740.060000 0.800000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 744.820000 0.000000 745.120000 0.800000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 750.340000 0.000000 750.640000 0.800000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 755.400000 0.000000 755.700000 0.800000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 760.460000 0.000000 760.760000 0.800000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 765.520000 0.000000 765.820000 0.800000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 770.580000 0.000000 770.880000 0.800000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 776.100000 0.000000 776.400000 0.800000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 781.160000 0.000000 781.460000 0.800000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 786.220000 0.000000 786.520000 0.800000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 791.280000 0.000000 791.580000 0.800000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.800000 0.000000 797.100000 0.800000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 801.860000 0.000000 802.160000 0.800000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 806.920000 0.000000 807.220000 0.800000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 811.980000 0.000000 812.280000 0.800000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.500000 0.000000 817.800000 0.800000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 822.560000 0.000000 822.860000 0.800000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 827.620000 0.000000 827.920000 0.800000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 832.680000 0.000000 832.980000 0.800000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 838.200000 0.000000 838.500000 0.800000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 843.260000 0.000000 843.560000 0.800000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 848.320000 0.000000 848.620000 0.800000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 853.380000 0.000000 853.680000 0.800000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 858.900000 0.000000 859.200000 0.800000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 863.960000 0.000000 864.260000 0.800000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 869.020000 0.000000 869.320000 0.800000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 874.080000 0.000000 874.380000 0.800000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 879.600000 0.000000 879.900000 0.800000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 884.660000 0.000000 884.960000 0.800000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 889.720000 0.000000 890.020000 0.800000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.780000 0.000000 895.080000 0.800000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 900.300000 0.000000 900.600000 0.800000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 905.360000 0.000000 905.660000 0.800000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 910.420000 0.000000 910.720000 0.800000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 915.480000 0.000000 915.780000 0.800000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 920.540000 0.000000 920.840000 0.800000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 926.060000 0.000000 926.360000 0.800000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 931.120000 0.000000 931.420000 0.800000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 936.180000 0.000000 936.480000 0.800000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 941.240000 0.000000 941.540000 0.800000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 946.760000 0.000000 947.060000 0.800000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 951.820000 0.000000 952.120000 0.800000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 956.880000 0.000000 957.180000 0.800000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 961.940000 0.000000 962.240000 0.800000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 967.460000 0.000000 967.760000 0.800000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 972.520000 0.000000 972.820000 0.800000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 977.580000 0.000000 977.880000 0.800000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 982.640000 0.000000 982.940000 0.800000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 988.160000 0.000000 988.460000 0.800000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.220000 0.000000 993.520000 0.800000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 998.280000 0.000000 998.580000 0.800000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1003.340000 0.000000 1003.640000 0.800000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1008.860000 0.000000 1009.160000 0.800000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1013.920000 0.000000 1014.220000 0.800000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1018.980000 0.000000 1019.280000 0.800000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1024.040000 0.000000 1024.340000 0.800000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1029.560000 0.000000 1029.860000 0.800000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1034.620000 0.000000 1034.920000 0.800000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1039.680000 0.000000 1039.980000 0.800000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1044.740000 0.000000 1045.040000 0.800000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1050.260000 0.000000 1050.560000 0.800000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1055.320000 0.000000 1055.620000 0.800000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1060.380000 0.000000 1060.680000 0.800000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1065.440000 0.000000 1065.740000 0.800000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1070.500000 0.000000 1070.800000 0.800000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1076.020000 0.000000 1076.320000 0.800000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1081.080000 0.000000 1081.380000 0.800000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1086.140000 0.000000 1086.440000 0.800000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1091.200000 0.000000 1091.500000 0.800000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.720000 0.000000 1097.020000 0.800000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1101.780000 0.000000 1102.080000 0.800000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1106.840000 0.000000 1107.140000 0.800000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1111.900000 0.000000 1112.200000 0.800000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1117.420000 0.000000 1117.720000 0.800000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1122.480000 0.000000 1122.780000 0.800000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1127.540000 0.000000 1127.840000 0.800000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1132.600000 0.000000 1132.900000 0.800000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1138.120000 0.000000 1138.420000 0.800000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1143.180000 0.000000 1143.480000 0.800000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1148.240000 0.000000 1148.540000 0.800000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1153.300000 0.000000 1153.600000 0.800000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1158.820000 0.000000 1159.120000 0.800000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1163.880000 0.000000 1164.180000 0.800000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1168.940000 0.000000 1169.240000 0.800000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1174.000000 0.000000 1174.300000 0.800000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1179.520000 0.000000 1179.820000 0.800000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1184.580000 0.000000 1184.880000 0.800000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1189.640000 0.000000 1189.940000 0.800000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1194.700000 0.000000 1195.000000 0.800000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1200.220000 0.000000 1200.520000 0.800000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1205.280000 0.000000 1205.580000 0.800000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1210.340000 0.000000 1210.640000 0.800000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1215.400000 0.000000 1215.700000 0.800000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1220.460000 0.000000 1220.760000 0.800000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 742.490000 0.800000 742.790000 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 28.4304 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 153.04 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 711.990000 0.800000 712.290000 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.8946 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 149.712 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 680.880000 0.800000 681.180000 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.4228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 173.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 649.770000 0.800000 650.070000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.1438 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 107.904 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 618.660000 0.800000 618.960000 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 588.160000 0.800000 588.460000 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 557.050000 0.800000 557.350000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 525.940000 0.800000 526.240000 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.6318 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.84 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 495.440000 0.800000 495.740000 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.816 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 464.330000 0.800000 464.630000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.6318 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.84 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 433.220000 0.800000 433.520000 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.1358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.528 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 402.720000 0.800000 403.020000 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.5018 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.48 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 371.610000 0.800000 371.910000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 200.063 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1067.94 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 340.500000 0.800000 340.800000 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 67.6086 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 361.52 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1631.240000 1639.360000 1631.540000 1640.160000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 30.8358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 164.928 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1580.640000 1639.360000 1580.940000 1640.160000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 47.6718 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 254.72 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1529.580000 1639.360000 1529.880000 1640.160000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 37.6251 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 201.608 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1478.520000 1639.360000 1478.820000 1640.160000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.3686 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 168.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1427.460000 1639.360000 1427.760000 1640.160000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.7748 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 281.936 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1376.400000 1639.360000 1376.700000 1640.160000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.7768 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 239.28 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1325.340000 1639.360000 1325.640000 1640.160000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.4446 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 243.312 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1274.740000 1639.360000 1275.040000 1640.160000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1223.680000 1639.360000 1223.980000 1640.160000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 1286.000000 2549.780000 1286.300000 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.6408 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.888 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 1329.920000 2549.780000 1330.220000 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0108 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.528 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 1374.450000 2549.780000 1374.750000 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.4698 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.976 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 1418.370000 2549.780000 1418.670000 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0108 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.528 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 1462.900000 2549.780000 1463.200000 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 1507.430000 2549.780000 1507.730000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1172.620000 1639.360000 1172.920000 1640.160000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.3946 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 189.712 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1121.560000 1639.360000 1121.860000 1640.160000 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1070.500000 1639.360000 1070.800000 1640.160000 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.1938 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 1551.350000 2549.780000 1551.650000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1019.440000 1639.360000 1019.740000 1640.160000 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 968.380000 1639.360000 968.680000 1640.160000 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 28.2708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 151.248 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 917.780000 1639.360000 918.080000 1640.160000 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 1595.880000 2549.780000 1596.180000 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 866.720000 1639.360000 867.020000 1640.160000 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.559 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.69 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1608.690000 0.800000 1608.990000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7698 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.576 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1577.580000 0.800000 1577.880000 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.2738 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.264 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1546.470000 0.800000 1546.770000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.3188 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1515.970000 0.800000 1516.270000 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.9978 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.792 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1484.860000 0.800000 1485.160000 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.1328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 166.512 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1453.750000 0.800000 1454.050000 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.5958 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 147.648 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1423.250000 0.800000 1423.550000 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.6788 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.424 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1392.140000 0.800000 1392.440000 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.1358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.528 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1361.030000 0.800000 1361.330000 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7698 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.576 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1330.530000 0.800000 1330.830000 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.9978 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.792 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1299.420000 0.800000 1299.720000 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.6318 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.84 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1268.310000 0.800000 1268.610000 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.816 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1237.200000 0.800000 1237.500000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.1008 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 129.008 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1206.700000 0.800000 1207.000000 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 60.8121 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 325.272 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2545.260000 1639.360000 2545.560000 1640.160000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 55.1148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 294.416 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2498.340000 1639.360000 2498.640000 1640.160000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.9248 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 122.736 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2447.280000 1639.360000 2447.580000 1640.160000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 57.1878 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 305.472 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2396.220000 1639.360000 2396.520000 1640.160000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.7738 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 239.264 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2345.160000 1639.360000 2345.460000 1640.160000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 41.6706 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 223.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2294.100000 1639.360000 2294.400000 1640.160000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 30.7236 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 164.8 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2243.040000 1639.360000 2243.340000 1640.160000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 47.3928 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 253.232 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2192.440000 1639.360000 2192.740000 1640.160000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 114.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 612.352 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2141.380000 1639.360000 2141.680000 1640.160000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.2018 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.88 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 6.830000 2549.780000 7.130000 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.6172 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 18.0563 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 101.822 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 45.260000 2549.780000 45.560000 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.6172 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 18.0563 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 101.822 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 89.790000 2549.780000 90.090000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.6172 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 18.0563 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 101.822 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 133.710000 2549.780000 134.010000 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.6172 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 18.0563 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 101.822 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 178.240000 2549.780000 178.540000 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.1968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.52 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 222.770000 2549.780000 223.070000 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.6078 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.712 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 266.690000 2549.780000 266.990000 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.6172 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 18.0563 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 101.822 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 311.220000 2549.780000 311.520000 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.5148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.216 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 355.140000 2549.780000 355.440000 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.6172 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 18.0563 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 101.822 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 399.670000 2549.780000 399.970000 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.1938 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 444.200000 2549.780000 444.500000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.3318 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 488.120000 2549.780000 488.420000 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.6922 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 18.0563 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 101.822 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 532.650000 2549.780000 532.950000 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.3798 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.496 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 577.180000 2549.780000 577.480000 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.7908 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 621.100000 2549.780000 621.400000 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.6592 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.128 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 18.0563 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 101.822 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2548.020000 0.000000 2548.320000 0.800000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.8544 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.552 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1175.590000 0.800000 1175.890000 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.7974 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.248 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1144.480000 0.800000 1144.780000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.4284 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.28 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1113.980000 0.800000 1114.280000 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.4764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.536 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1082.870000 0.800000 1083.170000 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.559 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.69 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1051.760000 0.800000 1052.060000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.559 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.69 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1021.260000 0.800000 1021.560000 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.559 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.69 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 990.150000 0.800000 990.450000 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.7164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.816 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 959.040000 0.800000 959.340000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.2004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.064 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 927.930000 0.800000 928.230000 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.3384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.8 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 897.430000 0.800000 897.730000 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.1644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 866.320000 0.800000 866.620000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.6144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.272 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 835.210000 0.800000 835.510000 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.904 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 804.710000 0.800000 805.010000 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.8764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.336 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 773.600000 0.800000 773.900000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 30.9286 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 164.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.7398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2090.320000 1639.360000 2090.620000 1640.160000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 47.2812 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 252.632 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2039.260000 1639.360000 2039.560000 1640.160000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 49.6044 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 264.552 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1988.200000 1639.360000 1988.500000 1640.160000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 47.4774 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 253.208 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1937.140000 1639.360000 1937.440000 1640.160000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 56.3412 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 300.952 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1886.540000 1639.360000 1886.840000 1640.160000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 59.0112 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 315.192 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1835.480000 1639.360000 1835.780000 1640.160000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 63.1254 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 336.664 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1784.420000 1639.360000 1784.720000 1640.160000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.4004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 88.424 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1733.360000 1639.360000 1733.660000 1640.160000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.3554 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.704 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1682.300000 1639.360000 1682.600000 1640.160000 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.01343 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.376 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 665.630000 2549.780000 665.930000 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.93843 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.976 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 709.550000 2549.780000 709.850000 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.01343 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.376 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 754.080000 2549.780000 754.380000 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.01343 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.376 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 798.610000 2549.780000 798.910000 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.1184 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.96 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 842.530000 2549.780000 842.830000 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.1664 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.216 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 887.060000 2549.780000 887.360000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.01343 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.376 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 931.590000 2549.780000 931.890000 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.6922 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 18.0563 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 101.822 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 975.510000 2549.780000 975.810000 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.01343 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.376 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 1020.040000 2549.780000 1020.340000 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.6922 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 18.0563 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 101.822 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 1063.960000 2549.780000 1064.260000 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.6922 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 18.0563 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 101.822 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 1108.490000 2549.780000 1108.790000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.89342 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.256 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 1153.020000 2549.780000 1153.320000 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.2004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.064 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 1196.940000 2549.780000 1197.240000 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.5722 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.184 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.426 LAYER met4  ;
    ANTENNAMAXAREACAR 18.0563 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 101.822 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 1241.470000 2549.780000 1241.770000 ;
    END
  END io_oeb[0]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 309.390000 0.800000 309.690000 ;
    END
  END analog_io[28]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 278.890000 0.800000 279.190000 ;
    END
  END analog_io[27]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 247.780000 0.800000 248.080000 ;
    END
  END analog_io[26]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 216.670000 0.800000 216.970000 ;
    END
  END analog_io[25]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 186.170000 0.800000 186.470000 ;
    END
  END analog_io[24]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 155.060000 0.800000 155.360000 ;
    END
  END analog_io[23]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 123.950000 0.800000 124.250000 ;
    END
  END analog_io[22]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 93.450000 0.800000 93.750000 ;
    END
  END analog_io[21]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 62.340000 0.800000 62.640000 ;
    END
  END analog_io[20]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 31.230000 0.800000 31.530000 ;
    END
  END analog_io[19]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1.950000 0.800000 2.250000 ;
    END
  END analog_io[18]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 815.660000 1639.360000 815.960000 1640.160000 ;
    END
  END analog_io[17]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 764.600000 1639.360000 764.900000 1640.160000 ;
    END
  END analog_io[16]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 713.540000 1639.360000 713.840000 1640.160000 ;
    END
  END analog_io[15]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 662.480000 1639.360000 662.780000 1640.160000 ;
    END
  END analog_io[14]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 611.880000 1639.360000 612.180000 1640.160000 ;
    END
  END analog_io[13]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 560.820000 1639.360000 561.120000 1640.160000 ;
    END
  END analog_io[12]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 509.760000 1639.360000 510.060000 1640.160000 ;
    END
  END analog_io[11]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 458.700000 1639.360000 459.000000 1640.160000 ;
    END
  END analog_io[10]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 407.640000 1639.360000 407.940000 1640.160000 ;
    END
  END analog_io[9]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.580000 1639.360000 356.880000 1640.160000 ;
    END
  END analog_io[8]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 305.980000 1639.360000 306.280000 1640.160000 ;
    END
  END analog_io[7]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.920000 1639.360000 255.220000 1640.160000 ;
    END
  END analog_io[6]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 203.860000 1639.360000 204.160000 1640.160000 ;
    END
  END analog_io[5]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 152.800000 1639.360000 153.100000 1640.160000 ;
    END
  END analog_io[4]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.740000 1639.360000 102.040000 1640.160000 ;
    END
  END analog_io[3]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 50.680000 1639.360000 50.980000 1640.160000 ;
    END
  END analog_io[2]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2548.980000 1637.360000 2549.780000 1637.660000 ;
    END
  END analog_io[1]
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 4.220000 1639.360000 4.520000 1640.160000 ;
    END
  END analog_io[0]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 558.980000 0.000000 559.280000 0.800000 ;
    END
  END user_clock2
  PIN user_irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.549 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 543.340000 0.000000 543.640000 0.800000 ;
    END
  END user_irq[2]
  PIN user_irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.53 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 548.400000 0.000000 548.700000 0.800000 ;
    END
  END user_irq[1]
  PIN user_irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 196.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.53 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 553.460000 0.000000 553.760000 0.800000 ;
    END
  END user_irq[0]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2544.460000 3.460000 2546.060000 1634.660000 ;
    END
    PORT
      LAYER met4 ;
        RECT 3.720000 3.460000 5.320000 1634.660000 ;
    END

# P/G pin shape extracted from block 'azadi_soc_top'
    PORT
      LAYER met4 ;
        RECT 57.555000 1189.800000 59.295000 1584.580000 ;
      LAYER met4 ;
        RECT 532.875000 1189.800000 534.615000 1584.580000 ;
    END
    PORT
      LAYER met4 ;
        RECT 707.335000 1189.800000 709.075000 1584.580000 ;
      LAYER met4 ;
        RECT 1182.655000 1189.800000 1184.395000 1584.580000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1357.115000 1189.800000 1358.855000 1584.580000 ;
      LAYER met4 ;
        RECT 1832.435000 1189.800000 1834.175000 1584.580000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2006.895000 1189.800000 2008.635000 1584.580000 ;
      LAYER met4 ;
        RECT 2482.215000 1189.800000 2483.955000 1584.580000 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.355000 688.015000 58.095000 1082.795000 ;
      LAYER met4 ;
        RECT 531.675000 688.015000 533.415000 1082.795000 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.355000 130.515000 58.095000 525.295000 ;
      LAYER met4 ;
        RECT 531.675000 130.515000 533.415000 525.295000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2006.465000 130.535000 2008.205000 525.315000 ;
      LAYER met4 ;
        RECT 2481.785000 130.535000 2483.525000 525.315000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2006.465000 688.035000 2008.205000 1082.815000 ;
      LAYER met4 ;
        RECT 2481.785000 688.035000 2483.525000 1082.815000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2502.326000 32.075000 2506.325000 1602.635000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2508.325000 26.075000 2512.325000 1608.635000 ;
    END
# end of P/G pin shape extracted from block 'azadi_soc_top'

  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2541.260000 6.660000 2542.860000 1631.460000 ;
    END
    PORT
      LAYER met4 ;
        RECT 6.920000 6.660000 8.520000 1631.460000 ;
    END

# P/G pin shape extracted from block 'azadi_soc_top'
    PORT
      LAYER met4 ;
        RECT 529.475000 1193.200000 531.215000 1581.180000 ;
      LAYER met4 ;
        RECT 60.955000 1193.200000 62.695000 1581.180000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1179.255000 1193.200000 1180.995000 1581.180000 ;
      LAYER met4 ;
        RECT 710.735000 1193.200000 712.475000 1581.180000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1829.035000 1193.200000 1830.775000 1581.180000 ;
      LAYER met4 ;
        RECT 1360.515000 1193.200000 1362.255000 1581.180000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2478.815000 1193.200000 2480.555000 1581.180000 ;
      LAYER met4 ;
        RECT 2010.295000 1193.200000 2012.035000 1581.180000 ;
    END
    PORT
      LAYER met4 ;
        RECT 528.275000 691.415000 530.015000 1079.395000 ;
      LAYER met4 ;
        RECT 59.755000 691.415000 61.495000 1079.395000 ;
    END
    PORT
      LAYER met4 ;
        RECT 528.275000 133.915000 530.015000 521.895000 ;
      LAYER met4 ;
        RECT 59.755000 133.915000 61.495000 521.895000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2478.385000 133.935000 2480.125000 521.915000 ;
      LAYER met4 ;
        RECT 2009.865000 133.935000 2011.605000 521.915000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2478.385000 691.435000 2480.125000 1079.415000 ;
      LAYER met4 ;
        RECT 2009.865000 691.435000 2011.605000 1079.415000 ;
    END
    PORT
      LAYER met4 ;
        RECT 34.885000 32.075000 38.885000 1602.635000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2502.325000 32.075000 2506.325000 1602.635000 ;
    END
# end of P/G pin shape extracted from block 'azadi_soc_top'

  END vccd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 2549.780000 1640.160000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 2549.780000 1640.160000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 2549.780000 1640.160000 ;
    LAYER met3 ;
      RECT 2545.860000 1639.060000 2549.780000 1640.160000 ;
      RECT 2498.940000 1639.060000 2544.960000 1640.160000 ;
      RECT 2447.880000 1639.060000 2498.040000 1640.160000 ;
      RECT 2396.820000 1639.060000 2446.980000 1640.160000 ;
      RECT 2345.760000 1639.060000 2395.920000 1640.160000 ;
      RECT 2294.700000 1639.060000 2344.860000 1640.160000 ;
      RECT 2243.640000 1639.060000 2293.800000 1640.160000 ;
      RECT 2193.040000 1639.060000 2242.740000 1640.160000 ;
      RECT 2141.980000 1639.060000 2192.140000 1640.160000 ;
      RECT 2090.920000 1639.060000 2141.080000 1640.160000 ;
      RECT 2039.860000 1639.060000 2090.020000 1640.160000 ;
      RECT 1988.800000 1639.060000 2038.960000 1640.160000 ;
      RECT 1937.740000 1639.060000 1987.900000 1640.160000 ;
      RECT 1887.140000 1639.060000 1936.840000 1640.160000 ;
      RECT 1836.080000 1639.060000 1886.240000 1640.160000 ;
      RECT 1785.020000 1639.060000 1835.180000 1640.160000 ;
      RECT 1733.960000 1639.060000 1784.120000 1640.160000 ;
      RECT 1682.900000 1639.060000 1733.060000 1640.160000 ;
      RECT 1631.840000 1639.060000 1682.000000 1640.160000 ;
      RECT 1581.240000 1639.060000 1630.940000 1640.160000 ;
      RECT 1530.180000 1639.060000 1580.340000 1640.160000 ;
      RECT 1479.120000 1639.060000 1529.280000 1640.160000 ;
      RECT 1428.060000 1639.060000 1478.220000 1640.160000 ;
      RECT 1377.000000 1639.060000 1427.160000 1640.160000 ;
      RECT 1325.940000 1639.060000 1376.100000 1640.160000 ;
      RECT 1275.340000 1639.060000 1325.040000 1640.160000 ;
      RECT 1224.280000 1639.060000 1274.440000 1640.160000 ;
      RECT 1173.220000 1639.060000 1223.380000 1640.160000 ;
      RECT 1122.160000 1639.060000 1172.320000 1640.160000 ;
      RECT 1071.100000 1639.060000 1121.260000 1640.160000 ;
      RECT 1020.040000 1639.060000 1070.200000 1640.160000 ;
      RECT 968.980000 1639.060000 1019.140000 1640.160000 ;
      RECT 918.380000 1639.060000 968.080000 1640.160000 ;
      RECT 867.320000 1639.060000 917.480000 1640.160000 ;
      RECT 816.260000 1639.060000 866.420000 1640.160000 ;
      RECT 765.200000 1639.060000 815.360000 1640.160000 ;
      RECT 714.140000 1639.060000 764.300000 1640.160000 ;
      RECT 663.080000 1639.060000 713.240000 1640.160000 ;
      RECT 612.480000 1639.060000 662.180000 1640.160000 ;
      RECT 561.420000 1639.060000 611.580000 1640.160000 ;
      RECT 510.360000 1639.060000 560.520000 1640.160000 ;
      RECT 459.300000 1639.060000 509.460000 1640.160000 ;
      RECT 408.240000 1639.060000 458.400000 1640.160000 ;
      RECT 357.180000 1639.060000 407.340000 1640.160000 ;
      RECT 306.580000 1639.060000 356.280000 1640.160000 ;
      RECT 255.520000 1639.060000 305.680000 1640.160000 ;
      RECT 204.460000 1639.060000 254.620000 1640.160000 ;
      RECT 153.400000 1639.060000 203.560000 1640.160000 ;
      RECT 102.340000 1639.060000 152.500000 1640.160000 ;
      RECT 51.280000 1639.060000 101.440000 1640.160000 ;
      RECT 4.820000 1639.060000 50.380000 1640.160000 ;
      RECT 0.000000 1639.060000 3.920000 1640.160000 ;
      RECT 0.000000 1638.570000 2549.780000 1639.060000 ;
      RECT 1.100000 1637.960000 2549.780000 1638.570000 ;
      RECT 1.100000 1637.670000 2548.680000 1637.960000 ;
      RECT 0.000000 1637.060000 2548.680000 1637.670000 ;
      RECT 0.000000 1609.290000 2549.780000 1637.060000 ;
      RECT 1.100000 1608.390000 2549.780000 1609.290000 ;
      RECT 0.000000 1596.480000 2549.780000 1608.390000 ;
      RECT 0.000000 1595.580000 2548.680000 1596.480000 ;
      RECT 0.000000 1578.180000 2549.780000 1595.580000 ;
      RECT 1.100000 1577.280000 2549.780000 1578.180000 ;
      RECT 0.000000 1551.950000 2549.780000 1577.280000 ;
      RECT 0.000000 1551.050000 2548.680000 1551.950000 ;
      RECT 0.000000 1547.070000 2549.780000 1551.050000 ;
      RECT 1.100000 1546.170000 2549.780000 1547.070000 ;
      RECT 0.000000 1516.570000 2549.780000 1546.170000 ;
      RECT 1.100000 1515.670000 2549.780000 1516.570000 ;
      RECT 0.000000 1508.030000 2549.780000 1515.670000 ;
      RECT 0.000000 1507.130000 2548.680000 1508.030000 ;
      RECT 0.000000 1485.460000 2549.780000 1507.130000 ;
      RECT 1.100000 1484.560000 2549.780000 1485.460000 ;
      RECT 0.000000 1463.500000 2549.780000 1484.560000 ;
      RECT 0.000000 1462.600000 2548.680000 1463.500000 ;
      RECT 0.000000 1454.350000 2549.780000 1462.600000 ;
      RECT 1.100000 1453.450000 2549.780000 1454.350000 ;
      RECT 0.000000 1423.850000 2549.780000 1453.450000 ;
      RECT 1.100000 1422.950000 2549.780000 1423.850000 ;
      RECT 0.000000 1418.970000 2549.780000 1422.950000 ;
      RECT 0.000000 1418.070000 2548.680000 1418.970000 ;
      RECT 0.000000 1392.740000 2549.780000 1418.070000 ;
      RECT 1.100000 1391.840000 2549.780000 1392.740000 ;
      RECT 0.000000 1375.050000 2549.780000 1391.840000 ;
      RECT 0.000000 1374.150000 2548.680000 1375.050000 ;
      RECT 0.000000 1361.630000 2549.780000 1374.150000 ;
      RECT 1.100000 1360.730000 2549.780000 1361.630000 ;
      RECT 0.000000 1331.130000 2549.780000 1360.730000 ;
      RECT 1.100000 1330.520000 2549.780000 1331.130000 ;
      RECT 1.100000 1330.230000 2548.680000 1330.520000 ;
      RECT 0.000000 1329.620000 2548.680000 1330.230000 ;
      RECT 0.000000 1300.020000 2549.780000 1329.620000 ;
      RECT 1.100000 1299.120000 2549.780000 1300.020000 ;
      RECT 0.000000 1286.600000 2549.780000 1299.120000 ;
      RECT 0.000000 1285.700000 2548.680000 1286.600000 ;
      RECT 0.000000 1268.910000 2549.780000 1285.700000 ;
      RECT 1.100000 1268.010000 2549.780000 1268.910000 ;
      RECT 0.000000 1242.070000 2549.780000 1268.010000 ;
      RECT 0.000000 1241.170000 2548.680000 1242.070000 ;
      RECT 0.000000 1237.800000 2549.780000 1241.170000 ;
      RECT 1.100000 1236.900000 2549.780000 1237.800000 ;
      RECT 0.000000 1207.300000 2549.780000 1236.900000 ;
      RECT 1.100000 1206.400000 2549.780000 1207.300000 ;
      RECT 0.000000 1197.540000 2549.780000 1206.400000 ;
      RECT 0.000000 1196.640000 2548.680000 1197.540000 ;
      RECT 0.000000 1176.190000 2549.780000 1196.640000 ;
      RECT 1.100000 1175.290000 2549.780000 1176.190000 ;
      RECT 0.000000 1153.620000 2549.780000 1175.290000 ;
      RECT 0.000000 1152.720000 2548.680000 1153.620000 ;
      RECT 0.000000 1145.080000 2549.780000 1152.720000 ;
      RECT 1.100000 1144.180000 2549.780000 1145.080000 ;
      RECT 0.000000 1114.580000 2549.780000 1144.180000 ;
      RECT 1.100000 1113.680000 2549.780000 1114.580000 ;
      RECT 0.000000 1109.090000 2549.780000 1113.680000 ;
      RECT 0.000000 1108.190000 2548.680000 1109.090000 ;
      RECT 0.000000 1083.470000 2549.780000 1108.190000 ;
      RECT 1.100000 1082.570000 2549.780000 1083.470000 ;
      RECT 0.000000 1064.560000 2549.780000 1082.570000 ;
      RECT 0.000000 1063.660000 2548.680000 1064.560000 ;
      RECT 0.000000 1052.360000 2549.780000 1063.660000 ;
      RECT 1.100000 1051.460000 2549.780000 1052.360000 ;
      RECT 0.000000 1021.860000 2549.780000 1051.460000 ;
      RECT 1.100000 1020.960000 2549.780000 1021.860000 ;
      RECT 0.000000 1020.640000 2549.780000 1020.960000 ;
      RECT 0.000000 1019.740000 2548.680000 1020.640000 ;
      RECT 0.000000 990.750000 2549.780000 1019.740000 ;
      RECT 1.100000 989.850000 2549.780000 990.750000 ;
      RECT 0.000000 976.110000 2549.780000 989.850000 ;
      RECT 0.000000 975.210000 2548.680000 976.110000 ;
      RECT 0.000000 959.640000 2549.780000 975.210000 ;
      RECT 1.100000 958.740000 2549.780000 959.640000 ;
      RECT 0.000000 932.190000 2549.780000 958.740000 ;
      RECT 0.000000 931.290000 2548.680000 932.190000 ;
      RECT 0.000000 928.530000 2549.780000 931.290000 ;
      RECT 1.100000 927.630000 2549.780000 928.530000 ;
      RECT 0.000000 898.030000 2549.780000 927.630000 ;
      RECT 1.100000 897.130000 2549.780000 898.030000 ;
      RECT 0.000000 887.660000 2549.780000 897.130000 ;
      RECT 0.000000 886.760000 2548.680000 887.660000 ;
      RECT 0.000000 866.920000 2549.780000 886.760000 ;
      RECT 1.100000 866.020000 2549.780000 866.920000 ;
      RECT 0.000000 843.130000 2549.780000 866.020000 ;
      RECT 0.000000 842.230000 2548.680000 843.130000 ;
      RECT 0.000000 835.810000 2549.780000 842.230000 ;
      RECT 1.100000 834.910000 2549.780000 835.810000 ;
      RECT 0.000000 805.310000 2549.780000 834.910000 ;
      RECT 1.100000 804.410000 2549.780000 805.310000 ;
      RECT 0.000000 799.210000 2549.780000 804.410000 ;
      RECT 0.000000 798.310000 2548.680000 799.210000 ;
      RECT 0.000000 774.200000 2549.780000 798.310000 ;
      RECT 1.100000 773.300000 2549.780000 774.200000 ;
      RECT 0.000000 754.680000 2549.780000 773.300000 ;
      RECT 0.000000 753.780000 2548.680000 754.680000 ;
      RECT 0.000000 743.090000 2549.780000 753.780000 ;
      RECT 1.100000 742.190000 2549.780000 743.090000 ;
      RECT 0.000000 712.590000 2549.780000 742.190000 ;
      RECT 1.100000 711.690000 2549.780000 712.590000 ;
      RECT 0.000000 710.150000 2549.780000 711.690000 ;
      RECT 0.000000 709.250000 2548.680000 710.150000 ;
      RECT 0.000000 681.480000 2549.780000 709.250000 ;
      RECT 1.100000 680.580000 2549.780000 681.480000 ;
      RECT 0.000000 666.230000 2549.780000 680.580000 ;
      RECT 0.000000 665.330000 2548.680000 666.230000 ;
      RECT 0.000000 650.370000 2549.780000 665.330000 ;
      RECT 1.100000 649.470000 2549.780000 650.370000 ;
      RECT 0.000000 621.700000 2549.780000 649.470000 ;
      RECT 0.000000 620.800000 2548.680000 621.700000 ;
      RECT 0.000000 619.260000 2549.780000 620.800000 ;
      RECT 1.100000 618.360000 2549.780000 619.260000 ;
      RECT 0.000000 588.760000 2549.780000 618.360000 ;
      RECT 1.100000 587.860000 2549.780000 588.760000 ;
      RECT 0.000000 577.780000 2549.780000 587.860000 ;
      RECT 0.000000 576.880000 2548.680000 577.780000 ;
      RECT 0.000000 557.650000 2549.780000 576.880000 ;
      RECT 1.100000 556.750000 2549.780000 557.650000 ;
      RECT 0.000000 533.250000 2549.780000 556.750000 ;
      RECT 0.000000 532.350000 2548.680000 533.250000 ;
      RECT 0.000000 526.540000 2549.780000 532.350000 ;
      RECT 1.100000 525.640000 2549.780000 526.540000 ;
      RECT 0.000000 496.040000 2549.780000 525.640000 ;
      RECT 1.100000 495.140000 2549.780000 496.040000 ;
      RECT 0.000000 488.720000 2549.780000 495.140000 ;
      RECT 0.000000 487.820000 2548.680000 488.720000 ;
      RECT 0.000000 464.930000 2549.780000 487.820000 ;
      RECT 1.100000 464.030000 2549.780000 464.930000 ;
      RECT 0.000000 444.800000 2549.780000 464.030000 ;
      RECT 0.000000 443.900000 2548.680000 444.800000 ;
      RECT 0.000000 433.820000 2549.780000 443.900000 ;
      RECT 1.100000 432.920000 2549.780000 433.820000 ;
      RECT 0.000000 403.320000 2549.780000 432.920000 ;
      RECT 1.100000 402.420000 2549.780000 403.320000 ;
      RECT 0.000000 400.270000 2549.780000 402.420000 ;
      RECT 0.000000 399.370000 2548.680000 400.270000 ;
      RECT 0.000000 372.210000 2549.780000 399.370000 ;
      RECT 1.100000 371.310000 2549.780000 372.210000 ;
      RECT 0.000000 355.740000 2549.780000 371.310000 ;
      RECT 0.000000 354.840000 2548.680000 355.740000 ;
      RECT 0.000000 341.100000 2549.780000 354.840000 ;
      RECT 1.100000 340.200000 2549.780000 341.100000 ;
      RECT 0.000000 311.820000 2549.780000 340.200000 ;
      RECT 0.000000 310.920000 2548.680000 311.820000 ;
      RECT 0.000000 309.990000 2549.780000 310.920000 ;
      RECT 1.100000 309.090000 2549.780000 309.990000 ;
      RECT 0.000000 279.490000 2549.780000 309.090000 ;
      RECT 1.100000 278.590000 2549.780000 279.490000 ;
      RECT 0.000000 267.290000 2549.780000 278.590000 ;
      RECT 0.000000 266.390000 2548.680000 267.290000 ;
      RECT 0.000000 248.380000 2549.780000 266.390000 ;
      RECT 1.100000 247.480000 2549.780000 248.380000 ;
      RECT 0.000000 223.370000 2549.780000 247.480000 ;
      RECT 0.000000 222.470000 2548.680000 223.370000 ;
      RECT 0.000000 217.270000 2549.780000 222.470000 ;
      RECT 1.100000 216.370000 2549.780000 217.270000 ;
      RECT 0.000000 186.770000 2549.780000 216.370000 ;
      RECT 1.100000 185.870000 2549.780000 186.770000 ;
      RECT 0.000000 178.840000 2549.780000 185.870000 ;
      RECT 0.000000 177.940000 2548.680000 178.840000 ;
      RECT 0.000000 155.660000 2549.780000 177.940000 ;
      RECT 1.100000 154.760000 2549.780000 155.660000 ;
      RECT 0.000000 134.310000 2549.780000 154.760000 ;
      RECT 0.000000 133.410000 2548.680000 134.310000 ;
      RECT 0.000000 124.550000 2549.780000 133.410000 ;
      RECT 1.100000 123.650000 2549.780000 124.550000 ;
      RECT 0.000000 94.050000 2549.780000 123.650000 ;
      RECT 1.100000 93.150000 2549.780000 94.050000 ;
      RECT 0.000000 90.390000 2549.780000 93.150000 ;
      RECT 0.000000 89.490000 2548.680000 90.390000 ;
      RECT 0.000000 62.940000 2549.780000 89.490000 ;
      RECT 1.100000 62.040000 2549.780000 62.940000 ;
      RECT 0.000000 45.860000 2549.780000 62.040000 ;
      RECT 0.000000 44.960000 2548.680000 45.860000 ;
      RECT 0.000000 31.830000 2549.780000 44.960000 ;
      RECT 1.100000 30.930000 2549.780000 31.830000 ;
      RECT 0.000000 7.430000 2549.780000 30.930000 ;
      RECT 0.000000 6.530000 2548.680000 7.430000 ;
      RECT 0.000000 2.550000 2549.780000 6.530000 ;
      RECT 1.100000 1.650000 2549.780000 2.550000 ;
      RECT 0.000000 1.100000 2549.780000 1.650000 ;
      RECT 2548.620000 0.000000 2549.780000 1.100000 ;
      RECT 2544.940000 0.000000 2547.720000 1.100000 ;
      RECT 2539.880000 0.000000 2544.040000 1.100000 ;
      RECT 2534.820000 0.000000 2538.980000 1.100000 ;
      RECT 2529.760000 0.000000 2533.920000 1.100000 ;
      RECT 2524.240000 0.000000 2528.860000 1.100000 ;
      RECT 2519.180000 0.000000 2523.340000 1.100000 ;
      RECT 2514.120000 0.000000 2518.280000 1.100000 ;
      RECT 2509.060000 0.000000 2513.220000 1.100000 ;
      RECT 2503.540000 0.000000 2508.160000 1.100000 ;
      RECT 2498.480000 0.000000 2502.640000 1.100000 ;
      RECT 2493.420000 0.000000 2497.580000 1.100000 ;
      RECT 2488.360000 0.000000 2492.520000 1.100000 ;
      RECT 2482.840000 0.000000 2487.460000 1.100000 ;
      RECT 2477.780000 0.000000 2481.940000 1.100000 ;
      RECT 2472.720000 0.000000 2476.880000 1.100000 ;
      RECT 2467.660000 0.000000 2471.820000 1.100000 ;
      RECT 2462.140000 0.000000 2466.760000 1.100000 ;
      RECT 2457.080000 0.000000 2461.240000 1.100000 ;
      RECT 2452.020000 0.000000 2456.180000 1.100000 ;
      RECT 2446.960000 0.000000 2451.120000 1.100000 ;
      RECT 2441.440000 0.000000 2446.060000 1.100000 ;
      RECT 2436.380000 0.000000 2440.540000 1.100000 ;
      RECT 2431.320000 0.000000 2435.480000 1.100000 ;
      RECT 2426.260000 0.000000 2430.420000 1.100000 ;
      RECT 2420.740000 0.000000 2425.360000 1.100000 ;
      RECT 2415.680000 0.000000 2419.840000 1.100000 ;
      RECT 2410.620000 0.000000 2414.780000 1.100000 ;
      RECT 2405.560000 0.000000 2409.720000 1.100000 ;
      RECT 2400.040000 0.000000 2404.660000 1.100000 ;
      RECT 2394.980000 0.000000 2399.140000 1.100000 ;
      RECT 2389.920000 0.000000 2394.080000 1.100000 ;
      RECT 2384.860000 0.000000 2389.020000 1.100000 ;
      RECT 2379.800000 0.000000 2383.960000 1.100000 ;
      RECT 2374.280000 0.000000 2378.900000 1.100000 ;
      RECT 2369.220000 0.000000 2373.380000 1.100000 ;
      RECT 2364.160000 0.000000 2368.320000 1.100000 ;
      RECT 2359.100000 0.000000 2363.260000 1.100000 ;
      RECT 2353.580000 0.000000 2358.200000 1.100000 ;
      RECT 2348.520000 0.000000 2352.680000 1.100000 ;
      RECT 2343.460000 0.000000 2347.620000 1.100000 ;
      RECT 2338.400000 0.000000 2342.560000 1.100000 ;
      RECT 2332.880000 0.000000 2337.500000 1.100000 ;
      RECT 2327.820000 0.000000 2331.980000 1.100000 ;
      RECT 2322.760000 0.000000 2326.920000 1.100000 ;
      RECT 2317.700000 0.000000 2321.860000 1.100000 ;
      RECT 2312.180000 0.000000 2316.800000 1.100000 ;
      RECT 2307.120000 0.000000 2311.280000 1.100000 ;
      RECT 2302.060000 0.000000 2306.220000 1.100000 ;
      RECT 2297.000000 0.000000 2301.160000 1.100000 ;
      RECT 2291.480000 0.000000 2296.100000 1.100000 ;
      RECT 2286.420000 0.000000 2290.580000 1.100000 ;
      RECT 2281.360000 0.000000 2285.520000 1.100000 ;
      RECT 2276.300000 0.000000 2280.460000 1.100000 ;
      RECT 2270.780000 0.000000 2275.400000 1.100000 ;
      RECT 2265.720000 0.000000 2269.880000 1.100000 ;
      RECT 2260.660000 0.000000 2264.820000 1.100000 ;
      RECT 2255.600000 0.000000 2259.760000 1.100000 ;
      RECT 2250.080000 0.000000 2254.700000 1.100000 ;
      RECT 2245.020000 0.000000 2249.180000 1.100000 ;
      RECT 2239.960000 0.000000 2244.120000 1.100000 ;
      RECT 2234.900000 0.000000 2239.060000 1.100000 ;
      RECT 2229.840000 0.000000 2234.000000 1.100000 ;
      RECT 2224.320000 0.000000 2228.940000 1.100000 ;
      RECT 2219.260000 0.000000 2223.420000 1.100000 ;
      RECT 2214.200000 0.000000 2218.360000 1.100000 ;
      RECT 2209.140000 0.000000 2213.300000 1.100000 ;
      RECT 2203.620000 0.000000 2208.240000 1.100000 ;
      RECT 2198.560000 0.000000 2202.720000 1.100000 ;
      RECT 2193.500000 0.000000 2197.660000 1.100000 ;
      RECT 2188.440000 0.000000 2192.600000 1.100000 ;
      RECT 2182.920000 0.000000 2187.540000 1.100000 ;
      RECT 2177.860000 0.000000 2182.020000 1.100000 ;
      RECT 2172.800000 0.000000 2176.960000 1.100000 ;
      RECT 2167.740000 0.000000 2171.900000 1.100000 ;
      RECT 2162.220000 0.000000 2166.840000 1.100000 ;
      RECT 2157.160000 0.000000 2161.320000 1.100000 ;
      RECT 2152.100000 0.000000 2156.260000 1.100000 ;
      RECT 2147.040000 0.000000 2151.200000 1.100000 ;
      RECT 2141.520000 0.000000 2146.140000 1.100000 ;
      RECT 2136.460000 0.000000 2140.620000 1.100000 ;
      RECT 2131.400000 0.000000 2135.560000 1.100000 ;
      RECT 2126.340000 0.000000 2130.500000 1.100000 ;
      RECT 2120.820000 0.000000 2125.440000 1.100000 ;
      RECT 2115.760000 0.000000 2119.920000 1.100000 ;
      RECT 2110.700000 0.000000 2114.860000 1.100000 ;
      RECT 2105.640000 0.000000 2109.800000 1.100000 ;
      RECT 2100.120000 0.000000 2104.740000 1.100000 ;
      RECT 2095.060000 0.000000 2099.220000 1.100000 ;
      RECT 2090.000000 0.000000 2094.160000 1.100000 ;
      RECT 2084.940000 0.000000 2089.100000 1.100000 ;
      RECT 2079.880000 0.000000 2084.040000 1.100000 ;
      RECT 2074.360000 0.000000 2078.980000 1.100000 ;
      RECT 2069.300000 0.000000 2073.460000 1.100000 ;
      RECT 2064.240000 0.000000 2068.400000 1.100000 ;
      RECT 2059.180000 0.000000 2063.340000 1.100000 ;
      RECT 2053.660000 0.000000 2058.280000 1.100000 ;
      RECT 2048.600000 0.000000 2052.760000 1.100000 ;
      RECT 2043.540000 0.000000 2047.700000 1.100000 ;
      RECT 2038.480000 0.000000 2042.640000 1.100000 ;
      RECT 2032.960000 0.000000 2037.580000 1.100000 ;
      RECT 2027.900000 0.000000 2032.060000 1.100000 ;
      RECT 2022.840000 0.000000 2027.000000 1.100000 ;
      RECT 2017.780000 0.000000 2021.940000 1.100000 ;
      RECT 2012.260000 0.000000 2016.880000 1.100000 ;
      RECT 2007.200000 0.000000 2011.360000 1.100000 ;
      RECT 2002.140000 0.000000 2006.300000 1.100000 ;
      RECT 1997.080000 0.000000 2001.240000 1.100000 ;
      RECT 1991.560000 0.000000 1996.180000 1.100000 ;
      RECT 1986.500000 0.000000 1990.660000 1.100000 ;
      RECT 1981.440000 0.000000 1985.600000 1.100000 ;
      RECT 1976.380000 0.000000 1980.540000 1.100000 ;
      RECT 1970.860000 0.000000 1975.480000 1.100000 ;
      RECT 1965.800000 0.000000 1969.960000 1.100000 ;
      RECT 1960.740000 0.000000 1964.900000 1.100000 ;
      RECT 1955.680000 0.000000 1959.840000 1.100000 ;
      RECT 1950.160000 0.000000 1954.780000 1.100000 ;
      RECT 1945.100000 0.000000 1949.260000 1.100000 ;
      RECT 1940.040000 0.000000 1944.200000 1.100000 ;
      RECT 1934.980000 0.000000 1939.140000 1.100000 ;
      RECT 1929.920000 0.000000 1934.080000 1.100000 ;
      RECT 1924.400000 0.000000 1929.020000 1.100000 ;
      RECT 1919.340000 0.000000 1923.500000 1.100000 ;
      RECT 1914.280000 0.000000 1918.440000 1.100000 ;
      RECT 1909.220000 0.000000 1913.380000 1.100000 ;
      RECT 1903.700000 0.000000 1908.320000 1.100000 ;
      RECT 1898.640000 0.000000 1902.800000 1.100000 ;
      RECT 1893.580000 0.000000 1897.740000 1.100000 ;
      RECT 1888.520000 0.000000 1892.680000 1.100000 ;
      RECT 1883.000000 0.000000 1887.620000 1.100000 ;
      RECT 1877.940000 0.000000 1882.100000 1.100000 ;
      RECT 1872.880000 0.000000 1877.040000 1.100000 ;
      RECT 1867.820000 0.000000 1871.980000 1.100000 ;
      RECT 1862.300000 0.000000 1866.920000 1.100000 ;
      RECT 1857.240000 0.000000 1861.400000 1.100000 ;
      RECT 1852.180000 0.000000 1856.340000 1.100000 ;
      RECT 1847.120000 0.000000 1851.280000 1.100000 ;
      RECT 1841.600000 0.000000 1846.220000 1.100000 ;
      RECT 1836.540000 0.000000 1840.700000 1.100000 ;
      RECT 1831.480000 0.000000 1835.640000 1.100000 ;
      RECT 1826.420000 0.000000 1830.580000 1.100000 ;
      RECT 1820.900000 0.000000 1825.520000 1.100000 ;
      RECT 1815.840000 0.000000 1820.000000 1.100000 ;
      RECT 1810.780000 0.000000 1814.940000 1.100000 ;
      RECT 1805.720000 0.000000 1809.880000 1.100000 ;
      RECT 1800.200000 0.000000 1804.820000 1.100000 ;
      RECT 1795.140000 0.000000 1799.300000 1.100000 ;
      RECT 1790.080000 0.000000 1794.240000 1.100000 ;
      RECT 1785.020000 0.000000 1789.180000 1.100000 ;
      RECT 1779.960000 0.000000 1784.120000 1.100000 ;
      RECT 1774.440000 0.000000 1779.060000 1.100000 ;
      RECT 1769.380000 0.000000 1773.540000 1.100000 ;
      RECT 1764.320000 0.000000 1768.480000 1.100000 ;
      RECT 1759.260000 0.000000 1763.420000 1.100000 ;
      RECT 1753.740000 0.000000 1758.360000 1.100000 ;
      RECT 1748.680000 0.000000 1752.840000 1.100000 ;
      RECT 1743.620000 0.000000 1747.780000 1.100000 ;
      RECT 1738.560000 0.000000 1742.720000 1.100000 ;
      RECT 1733.040000 0.000000 1737.660000 1.100000 ;
      RECT 1727.980000 0.000000 1732.140000 1.100000 ;
      RECT 1722.920000 0.000000 1727.080000 1.100000 ;
      RECT 1717.860000 0.000000 1722.020000 1.100000 ;
      RECT 1712.340000 0.000000 1716.960000 1.100000 ;
      RECT 1707.280000 0.000000 1711.440000 1.100000 ;
      RECT 1702.220000 0.000000 1706.380000 1.100000 ;
      RECT 1697.160000 0.000000 1701.320000 1.100000 ;
      RECT 1691.640000 0.000000 1696.260000 1.100000 ;
      RECT 1686.580000 0.000000 1690.740000 1.100000 ;
      RECT 1681.520000 0.000000 1685.680000 1.100000 ;
      RECT 1676.460000 0.000000 1680.620000 1.100000 ;
      RECT 1670.940000 0.000000 1675.560000 1.100000 ;
      RECT 1665.880000 0.000000 1670.040000 1.100000 ;
      RECT 1660.820000 0.000000 1664.980000 1.100000 ;
      RECT 1655.760000 0.000000 1659.920000 1.100000 ;
      RECT 1650.240000 0.000000 1654.860000 1.100000 ;
      RECT 1645.180000 0.000000 1649.340000 1.100000 ;
      RECT 1640.120000 0.000000 1644.280000 1.100000 ;
      RECT 1635.060000 0.000000 1639.220000 1.100000 ;
      RECT 1630.000000 0.000000 1634.160000 1.100000 ;
      RECT 1624.480000 0.000000 1629.100000 1.100000 ;
      RECT 1619.420000 0.000000 1623.580000 1.100000 ;
      RECT 1614.360000 0.000000 1618.520000 1.100000 ;
      RECT 1609.300000 0.000000 1613.460000 1.100000 ;
      RECT 1603.780000 0.000000 1608.400000 1.100000 ;
      RECT 1598.720000 0.000000 1602.880000 1.100000 ;
      RECT 1593.660000 0.000000 1597.820000 1.100000 ;
      RECT 1588.600000 0.000000 1592.760000 1.100000 ;
      RECT 1583.080000 0.000000 1587.700000 1.100000 ;
      RECT 1578.020000 0.000000 1582.180000 1.100000 ;
      RECT 1572.960000 0.000000 1577.120000 1.100000 ;
      RECT 1567.900000 0.000000 1572.060000 1.100000 ;
      RECT 1562.380000 0.000000 1567.000000 1.100000 ;
      RECT 1557.320000 0.000000 1561.480000 1.100000 ;
      RECT 1552.260000 0.000000 1556.420000 1.100000 ;
      RECT 1547.200000 0.000000 1551.360000 1.100000 ;
      RECT 1541.680000 0.000000 1546.300000 1.100000 ;
      RECT 1536.620000 0.000000 1540.780000 1.100000 ;
      RECT 1531.560000 0.000000 1535.720000 1.100000 ;
      RECT 1526.500000 0.000000 1530.660000 1.100000 ;
      RECT 1520.980000 0.000000 1525.600000 1.100000 ;
      RECT 1515.920000 0.000000 1520.080000 1.100000 ;
      RECT 1510.860000 0.000000 1515.020000 1.100000 ;
      RECT 1505.800000 0.000000 1509.960000 1.100000 ;
      RECT 1500.280000 0.000000 1504.900000 1.100000 ;
      RECT 1495.220000 0.000000 1499.380000 1.100000 ;
      RECT 1490.160000 0.000000 1494.320000 1.100000 ;
      RECT 1485.100000 0.000000 1489.260000 1.100000 ;
      RECT 1480.040000 0.000000 1484.200000 1.100000 ;
      RECT 1474.520000 0.000000 1479.140000 1.100000 ;
      RECT 1469.460000 0.000000 1473.620000 1.100000 ;
      RECT 1464.400000 0.000000 1468.560000 1.100000 ;
      RECT 1459.340000 0.000000 1463.500000 1.100000 ;
      RECT 1453.820000 0.000000 1458.440000 1.100000 ;
      RECT 1448.760000 0.000000 1452.920000 1.100000 ;
      RECT 1443.700000 0.000000 1447.860000 1.100000 ;
      RECT 1438.640000 0.000000 1442.800000 1.100000 ;
      RECT 1433.120000 0.000000 1437.740000 1.100000 ;
      RECT 1428.060000 0.000000 1432.220000 1.100000 ;
      RECT 1423.000000 0.000000 1427.160000 1.100000 ;
      RECT 1417.940000 0.000000 1422.100000 1.100000 ;
      RECT 1412.420000 0.000000 1417.040000 1.100000 ;
      RECT 1407.360000 0.000000 1411.520000 1.100000 ;
      RECT 1402.300000 0.000000 1406.460000 1.100000 ;
      RECT 1397.240000 0.000000 1401.400000 1.100000 ;
      RECT 1391.720000 0.000000 1396.340000 1.100000 ;
      RECT 1386.660000 0.000000 1390.820000 1.100000 ;
      RECT 1381.600000 0.000000 1385.760000 1.100000 ;
      RECT 1376.540000 0.000000 1380.700000 1.100000 ;
      RECT 1371.020000 0.000000 1375.640000 1.100000 ;
      RECT 1365.960000 0.000000 1370.120000 1.100000 ;
      RECT 1360.900000 0.000000 1365.060000 1.100000 ;
      RECT 1355.840000 0.000000 1360.000000 1.100000 ;
      RECT 1350.780000 0.000000 1354.940000 1.100000 ;
      RECT 1345.260000 0.000000 1349.880000 1.100000 ;
      RECT 1340.200000 0.000000 1344.360000 1.100000 ;
      RECT 1335.140000 0.000000 1339.300000 1.100000 ;
      RECT 1330.080000 0.000000 1334.240000 1.100000 ;
      RECT 1324.560000 0.000000 1329.180000 1.100000 ;
      RECT 1319.500000 0.000000 1323.660000 1.100000 ;
      RECT 1314.440000 0.000000 1318.600000 1.100000 ;
      RECT 1309.380000 0.000000 1313.540000 1.100000 ;
      RECT 1303.860000 0.000000 1308.480000 1.100000 ;
      RECT 1298.800000 0.000000 1302.960000 1.100000 ;
      RECT 1293.740000 0.000000 1297.900000 1.100000 ;
      RECT 1288.680000 0.000000 1292.840000 1.100000 ;
      RECT 1283.160000 0.000000 1287.780000 1.100000 ;
      RECT 1278.100000 0.000000 1282.260000 1.100000 ;
      RECT 1273.040000 0.000000 1277.200000 1.100000 ;
      RECT 1267.980000 0.000000 1272.140000 1.100000 ;
      RECT 1262.460000 0.000000 1267.080000 1.100000 ;
      RECT 1257.400000 0.000000 1261.560000 1.100000 ;
      RECT 1252.340000 0.000000 1256.500000 1.100000 ;
      RECT 1247.280000 0.000000 1251.440000 1.100000 ;
      RECT 1241.760000 0.000000 1246.380000 1.100000 ;
      RECT 1236.700000 0.000000 1240.860000 1.100000 ;
      RECT 1231.640000 0.000000 1235.800000 1.100000 ;
      RECT 1226.580000 0.000000 1230.740000 1.100000 ;
      RECT 1221.060000 0.000000 1225.680000 1.100000 ;
      RECT 1216.000000 0.000000 1220.160000 1.100000 ;
      RECT 1210.940000 0.000000 1215.100000 1.100000 ;
      RECT 1205.880000 0.000000 1210.040000 1.100000 ;
      RECT 1200.820000 0.000000 1204.980000 1.100000 ;
      RECT 1195.300000 0.000000 1199.920000 1.100000 ;
      RECT 1190.240000 0.000000 1194.400000 1.100000 ;
      RECT 1185.180000 0.000000 1189.340000 1.100000 ;
      RECT 1180.120000 0.000000 1184.280000 1.100000 ;
      RECT 1174.600000 0.000000 1179.220000 1.100000 ;
      RECT 1169.540000 0.000000 1173.700000 1.100000 ;
      RECT 1164.480000 0.000000 1168.640000 1.100000 ;
      RECT 1159.420000 0.000000 1163.580000 1.100000 ;
      RECT 1153.900000 0.000000 1158.520000 1.100000 ;
      RECT 1148.840000 0.000000 1153.000000 1.100000 ;
      RECT 1143.780000 0.000000 1147.940000 1.100000 ;
      RECT 1138.720000 0.000000 1142.880000 1.100000 ;
      RECT 1133.200000 0.000000 1137.820000 1.100000 ;
      RECT 1128.140000 0.000000 1132.300000 1.100000 ;
      RECT 1123.080000 0.000000 1127.240000 1.100000 ;
      RECT 1118.020000 0.000000 1122.180000 1.100000 ;
      RECT 1112.500000 0.000000 1117.120000 1.100000 ;
      RECT 1107.440000 0.000000 1111.600000 1.100000 ;
      RECT 1102.380000 0.000000 1106.540000 1.100000 ;
      RECT 1097.320000 0.000000 1101.480000 1.100000 ;
      RECT 1091.800000 0.000000 1096.420000 1.100000 ;
      RECT 1086.740000 0.000000 1090.900000 1.100000 ;
      RECT 1081.680000 0.000000 1085.840000 1.100000 ;
      RECT 1076.620000 0.000000 1080.780000 1.100000 ;
      RECT 1071.100000 0.000000 1075.720000 1.100000 ;
      RECT 1066.040000 0.000000 1070.200000 1.100000 ;
      RECT 1060.980000 0.000000 1065.140000 1.100000 ;
      RECT 1055.920000 0.000000 1060.080000 1.100000 ;
      RECT 1050.860000 0.000000 1055.020000 1.100000 ;
      RECT 1045.340000 0.000000 1049.960000 1.100000 ;
      RECT 1040.280000 0.000000 1044.440000 1.100000 ;
      RECT 1035.220000 0.000000 1039.380000 1.100000 ;
      RECT 1030.160000 0.000000 1034.320000 1.100000 ;
      RECT 1024.640000 0.000000 1029.260000 1.100000 ;
      RECT 1019.580000 0.000000 1023.740000 1.100000 ;
      RECT 1014.520000 0.000000 1018.680000 1.100000 ;
      RECT 1009.460000 0.000000 1013.620000 1.100000 ;
      RECT 1003.940000 0.000000 1008.560000 1.100000 ;
      RECT 998.880000 0.000000 1003.040000 1.100000 ;
      RECT 993.820000 0.000000 997.980000 1.100000 ;
      RECT 988.760000 0.000000 992.920000 1.100000 ;
      RECT 983.240000 0.000000 987.860000 1.100000 ;
      RECT 978.180000 0.000000 982.340000 1.100000 ;
      RECT 973.120000 0.000000 977.280000 1.100000 ;
      RECT 968.060000 0.000000 972.220000 1.100000 ;
      RECT 962.540000 0.000000 967.160000 1.100000 ;
      RECT 957.480000 0.000000 961.640000 1.100000 ;
      RECT 952.420000 0.000000 956.580000 1.100000 ;
      RECT 947.360000 0.000000 951.520000 1.100000 ;
      RECT 941.840000 0.000000 946.460000 1.100000 ;
      RECT 936.780000 0.000000 940.940000 1.100000 ;
      RECT 931.720000 0.000000 935.880000 1.100000 ;
      RECT 926.660000 0.000000 930.820000 1.100000 ;
      RECT 921.140000 0.000000 925.760000 1.100000 ;
      RECT 916.080000 0.000000 920.240000 1.100000 ;
      RECT 911.020000 0.000000 915.180000 1.100000 ;
      RECT 905.960000 0.000000 910.120000 1.100000 ;
      RECT 900.900000 0.000000 905.060000 1.100000 ;
      RECT 895.380000 0.000000 900.000000 1.100000 ;
      RECT 890.320000 0.000000 894.480000 1.100000 ;
      RECT 885.260000 0.000000 889.420000 1.100000 ;
      RECT 880.200000 0.000000 884.360000 1.100000 ;
      RECT 874.680000 0.000000 879.300000 1.100000 ;
      RECT 869.620000 0.000000 873.780000 1.100000 ;
      RECT 864.560000 0.000000 868.720000 1.100000 ;
      RECT 859.500000 0.000000 863.660000 1.100000 ;
      RECT 853.980000 0.000000 858.600000 1.100000 ;
      RECT 848.920000 0.000000 853.080000 1.100000 ;
      RECT 843.860000 0.000000 848.020000 1.100000 ;
      RECT 838.800000 0.000000 842.960000 1.100000 ;
      RECT 833.280000 0.000000 837.900000 1.100000 ;
      RECT 828.220000 0.000000 832.380000 1.100000 ;
      RECT 823.160000 0.000000 827.320000 1.100000 ;
      RECT 818.100000 0.000000 822.260000 1.100000 ;
      RECT 812.580000 0.000000 817.200000 1.100000 ;
      RECT 807.520000 0.000000 811.680000 1.100000 ;
      RECT 802.460000 0.000000 806.620000 1.100000 ;
      RECT 797.400000 0.000000 801.560000 1.100000 ;
      RECT 791.880000 0.000000 796.500000 1.100000 ;
      RECT 786.820000 0.000000 790.980000 1.100000 ;
      RECT 781.760000 0.000000 785.920000 1.100000 ;
      RECT 776.700000 0.000000 780.860000 1.100000 ;
      RECT 771.180000 0.000000 775.800000 1.100000 ;
      RECT 766.120000 0.000000 770.280000 1.100000 ;
      RECT 761.060000 0.000000 765.220000 1.100000 ;
      RECT 756.000000 0.000000 760.160000 1.100000 ;
      RECT 750.940000 0.000000 755.100000 1.100000 ;
      RECT 745.420000 0.000000 750.040000 1.100000 ;
      RECT 740.360000 0.000000 744.520000 1.100000 ;
      RECT 735.300000 0.000000 739.460000 1.100000 ;
      RECT 730.240000 0.000000 734.400000 1.100000 ;
      RECT 724.720000 0.000000 729.340000 1.100000 ;
      RECT 719.660000 0.000000 723.820000 1.100000 ;
      RECT 714.600000 0.000000 718.760000 1.100000 ;
      RECT 709.540000 0.000000 713.700000 1.100000 ;
      RECT 704.020000 0.000000 708.640000 1.100000 ;
      RECT 698.960000 0.000000 703.120000 1.100000 ;
      RECT 693.900000 0.000000 698.060000 1.100000 ;
      RECT 688.840000 0.000000 693.000000 1.100000 ;
      RECT 683.320000 0.000000 687.940000 1.100000 ;
      RECT 678.260000 0.000000 682.420000 1.100000 ;
      RECT 673.200000 0.000000 677.360000 1.100000 ;
      RECT 668.140000 0.000000 672.300000 1.100000 ;
      RECT 662.620000 0.000000 667.240000 1.100000 ;
      RECT 657.560000 0.000000 661.720000 1.100000 ;
      RECT 652.500000 0.000000 656.660000 1.100000 ;
      RECT 647.440000 0.000000 651.600000 1.100000 ;
      RECT 641.920000 0.000000 646.540000 1.100000 ;
      RECT 636.860000 0.000000 641.020000 1.100000 ;
      RECT 631.800000 0.000000 635.960000 1.100000 ;
      RECT 626.740000 0.000000 630.900000 1.100000 ;
      RECT 621.220000 0.000000 625.840000 1.100000 ;
      RECT 616.160000 0.000000 620.320000 1.100000 ;
      RECT 611.100000 0.000000 615.260000 1.100000 ;
      RECT 606.040000 0.000000 610.200000 1.100000 ;
      RECT 600.980000 0.000000 605.140000 1.100000 ;
      RECT 595.460000 0.000000 600.080000 1.100000 ;
      RECT 590.400000 0.000000 594.560000 1.100000 ;
      RECT 585.340000 0.000000 589.500000 1.100000 ;
      RECT 580.280000 0.000000 584.440000 1.100000 ;
      RECT 574.760000 0.000000 579.380000 1.100000 ;
      RECT 569.700000 0.000000 573.860000 1.100000 ;
      RECT 564.640000 0.000000 568.800000 1.100000 ;
      RECT 559.580000 0.000000 563.740000 1.100000 ;
      RECT 554.060000 0.000000 558.680000 1.100000 ;
      RECT 549.000000 0.000000 553.160000 1.100000 ;
      RECT 543.940000 0.000000 548.100000 1.100000 ;
      RECT 538.880000 0.000000 543.040000 1.100000 ;
      RECT 533.360000 0.000000 537.980000 1.100000 ;
      RECT 528.300000 0.000000 532.460000 1.100000 ;
      RECT 523.240000 0.000000 527.400000 1.100000 ;
      RECT 518.180000 0.000000 522.340000 1.100000 ;
      RECT 512.660000 0.000000 517.280000 1.100000 ;
      RECT 507.600000 0.000000 511.760000 1.100000 ;
      RECT 502.540000 0.000000 506.700000 1.100000 ;
      RECT 497.480000 0.000000 501.640000 1.100000 ;
      RECT 491.960000 0.000000 496.580000 1.100000 ;
      RECT 486.900000 0.000000 491.060000 1.100000 ;
      RECT 481.840000 0.000000 486.000000 1.100000 ;
      RECT 476.780000 0.000000 480.940000 1.100000 ;
      RECT 471.260000 0.000000 475.880000 1.100000 ;
      RECT 466.200000 0.000000 470.360000 1.100000 ;
      RECT 461.140000 0.000000 465.300000 1.100000 ;
      RECT 456.080000 0.000000 460.240000 1.100000 ;
      RECT 451.020000 0.000000 455.180000 1.100000 ;
      RECT 445.500000 0.000000 450.120000 1.100000 ;
      RECT 440.440000 0.000000 444.600000 1.100000 ;
      RECT 435.380000 0.000000 439.540000 1.100000 ;
      RECT 430.320000 0.000000 434.480000 1.100000 ;
      RECT 424.800000 0.000000 429.420000 1.100000 ;
      RECT 419.740000 0.000000 423.900000 1.100000 ;
      RECT 414.680000 0.000000 418.840000 1.100000 ;
      RECT 409.620000 0.000000 413.780000 1.100000 ;
      RECT 404.100000 0.000000 408.720000 1.100000 ;
      RECT 399.040000 0.000000 403.200000 1.100000 ;
      RECT 393.980000 0.000000 398.140000 1.100000 ;
      RECT 388.920000 0.000000 393.080000 1.100000 ;
      RECT 383.400000 0.000000 388.020000 1.100000 ;
      RECT 378.340000 0.000000 382.500000 1.100000 ;
      RECT 373.280000 0.000000 377.440000 1.100000 ;
      RECT 368.220000 0.000000 372.380000 1.100000 ;
      RECT 362.700000 0.000000 367.320000 1.100000 ;
      RECT 357.640000 0.000000 361.800000 1.100000 ;
      RECT 352.580000 0.000000 356.740000 1.100000 ;
      RECT 347.520000 0.000000 351.680000 1.100000 ;
      RECT 342.000000 0.000000 346.620000 1.100000 ;
      RECT 336.940000 0.000000 341.100000 1.100000 ;
      RECT 331.880000 0.000000 336.040000 1.100000 ;
      RECT 326.820000 0.000000 330.980000 1.100000 ;
      RECT 321.300000 0.000000 325.920000 1.100000 ;
      RECT 316.240000 0.000000 320.400000 1.100000 ;
      RECT 311.180000 0.000000 315.340000 1.100000 ;
      RECT 306.120000 0.000000 310.280000 1.100000 ;
      RECT 301.060000 0.000000 305.220000 1.100000 ;
      RECT 295.540000 0.000000 300.160000 1.100000 ;
      RECT 290.480000 0.000000 294.640000 1.100000 ;
      RECT 285.420000 0.000000 289.580000 1.100000 ;
      RECT 280.360000 0.000000 284.520000 1.100000 ;
      RECT 274.840000 0.000000 279.460000 1.100000 ;
      RECT 269.780000 0.000000 273.940000 1.100000 ;
      RECT 264.720000 0.000000 268.880000 1.100000 ;
      RECT 259.660000 0.000000 263.820000 1.100000 ;
      RECT 254.140000 0.000000 258.760000 1.100000 ;
      RECT 249.080000 0.000000 253.240000 1.100000 ;
      RECT 244.020000 0.000000 248.180000 1.100000 ;
      RECT 238.960000 0.000000 243.120000 1.100000 ;
      RECT 233.440000 0.000000 238.060000 1.100000 ;
      RECT 228.380000 0.000000 232.540000 1.100000 ;
      RECT 223.320000 0.000000 227.480000 1.100000 ;
      RECT 218.260000 0.000000 222.420000 1.100000 ;
      RECT 212.740000 0.000000 217.360000 1.100000 ;
      RECT 207.680000 0.000000 211.840000 1.100000 ;
      RECT 202.620000 0.000000 206.780000 1.100000 ;
      RECT 197.560000 0.000000 201.720000 1.100000 ;
      RECT 192.040000 0.000000 196.660000 1.100000 ;
      RECT 186.980000 0.000000 191.140000 1.100000 ;
      RECT 181.920000 0.000000 186.080000 1.100000 ;
      RECT 176.860000 0.000000 181.020000 1.100000 ;
      RECT 171.340000 0.000000 175.960000 1.100000 ;
      RECT 166.280000 0.000000 170.440000 1.100000 ;
      RECT 161.220000 0.000000 165.380000 1.100000 ;
      RECT 156.160000 0.000000 160.320000 1.100000 ;
      RECT 150.640000 0.000000 155.260000 1.100000 ;
      RECT 145.580000 0.000000 149.740000 1.100000 ;
      RECT 140.520000 0.000000 144.680000 1.100000 ;
      RECT 135.460000 0.000000 139.620000 1.100000 ;
      RECT 130.400000 0.000000 134.560000 1.100000 ;
      RECT 124.880000 0.000000 129.500000 1.100000 ;
      RECT 119.820000 0.000000 123.980000 1.100000 ;
      RECT 114.760000 0.000000 118.920000 1.100000 ;
      RECT 109.700000 0.000000 113.860000 1.100000 ;
      RECT 104.180000 0.000000 108.800000 1.100000 ;
      RECT 99.120000 0.000000 103.280000 1.100000 ;
      RECT 94.060000 0.000000 98.220000 1.100000 ;
      RECT 89.000000 0.000000 93.160000 1.100000 ;
      RECT 83.480000 0.000000 88.100000 1.100000 ;
      RECT 78.420000 0.000000 82.580000 1.100000 ;
      RECT 73.360000 0.000000 77.520000 1.100000 ;
      RECT 68.300000 0.000000 72.460000 1.100000 ;
      RECT 62.780000 0.000000 67.400000 1.100000 ;
      RECT 57.720000 0.000000 61.880000 1.100000 ;
      RECT 52.660000 0.000000 56.820000 1.100000 ;
      RECT 47.600000 0.000000 51.760000 1.100000 ;
      RECT 42.080000 0.000000 46.700000 1.100000 ;
      RECT 37.020000 0.000000 41.180000 1.100000 ;
      RECT 31.960000 0.000000 36.120000 1.100000 ;
      RECT 26.900000 0.000000 31.060000 1.100000 ;
      RECT 21.380000 0.000000 26.000000 1.100000 ;
      RECT 16.320000 0.000000 20.480000 1.100000 ;
      RECT 11.260000 0.000000 15.420000 1.100000 ;
      RECT 6.200000 0.000000 10.360000 1.100000 ;
      RECT 2.520000 0.000000 5.300000 1.100000 ;
      RECT 0.000000 0.000000 1.620000 1.100000 ;
    LAYER met4 ;
      RECT 0.000000 1634.960000 2549.780000 1640.160000 ;
      RECT 5.620000 1631.760000 2544.160000 1634.960000 ;
      RECT 2543.160000 6.360000 2544.160000 1631.760000 ;
      RECT 8.820000 6.360000 2540.960000 1631.760000 ;
      RECT 5.620000 6.360000 6.620000 1631.760000 ;
      RECT 2546.360000 3.160000 2549.780000 1634.960000 ;
      RECT 5.620000 3.160000 2544.160000 6.360000 ;
      RECT 0.000000 3.160000 3.420000 1634.960000 ;
      RECT 0.000000 0.000000 2549.780000 3.160000 ;
    LAYER met5 ;
      RECT 0.000000 0.000000 2549.780000 1640.160000 ;
  END
END azadi_soc_top_caravel

END LIBRARY
